VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_assaify_mssf_pll
  CLASS BLOCK ;
  FOREIGN tt_um_assaify_mssf_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.391500 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 40.340000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.900500 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.391500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.391500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.500 4.000 225.500 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 5.000 0.500 9.000 225.500 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 86.000 192.770 133.500 193.715 ;
        RECT 86.000 192.730 86.180 192.770 ;
        RECT 86.570 192.730 86.930 192.770 ;
        RECT 87.320 192.730 92.680 192.770 ;
        RECT 93.070 192.730 93.430 192.770 ;
        RECT 93.820 192.730 99.180 192.770 ;
        RECT 99.570 192.730 104.680 192.770 ;
        RECT 105.070 192.730 115.180 192.770 ;
        RECT 115.570 192.730 117.680 192.770 ;
        RECT 118.070 192.730 118.430 192.770 ;
        RECT 118.820 192.730 124.000 192.770 ;
        RECT 124.320 192.730 124.680 192.770 ;
        RECT 125.070 192.730 125.430 192.770 ;
        RECT 125.820 192.730 131.180 192.770 ;
        RECT 131.570 192.730 133.500 192.770 ;
        RECT 86.000 192.645 133.500 192.730 ;
      LAYER nwell ;
        RECT 86.000 190.795 133.500 192.315 ;
      LAYER pwell ;
        RECT 21.250 157.500 25.250 188.500 ;
        RECT 30.750 157.500 34.750 188.500 ;
        RECT 40.250 157.500 44.250 188.500 ;
        RECT 85.500 186.520 133.500 187.465 ;
        RECT 85.500 186.480 92.430 186.520 ;
        RECT 92.820 186.480 108.430 186.520 ;
        RECT 108.820 186.480 124.430 186.520 ;
        RECT 124.820 186.480 133.500 186.520 ;
        RECT 85.500 186.395 133.500 186.480 ;
      LAYER nwell ;
        RECT 85.500 184.545 133.500 186.065 ;
      LAYER pwell ;
        RECT 81.000 176.270 139.250 177.215 ;
        RECT 81.000 176.230 82.930 176.270 ;
        RECT 83.320 176.230 90.180 176.270 ;
        RECT 90.570 176.230 96.180 176.270 ;
        RECT 96.570 176.230 103.180 176.270 ;
        RECT 103.570 176.230 109.180 176.270 ;
        RECT 109.570 176.230 116.180 176.270 ;
        RECT 116.570 176.230 120.680 176.270 ;
        RECT 121.070 176.230 128.430 176.270 ;
        RECT 128.820 176.230 138.680 176.270 ;
        RECT 139.070 176.230 139.250 176.270 ;
        RECT 81.000 176.145 139.250 176.230 ;
      LAYER nwell ;
        RECT 81.000 174.295 139.250 175.815 ;
      LAYER pwell ;
        RECT 81.000 169.270 88.500 170.215 ;
        RECT 81.000 169.230 82.930 169.270 ;
        RECT 83.320 169.230 88.500 169.270 ;
        RECT 81.000 169.145 88.500 169.230 ;
        RECT 90.750 169.270 139.000 170.215 ;
        RECT 90.750 169.230 90.930 169.270 ;
        RECT 91.320 169.230 97.930 169.270 ;
        RECT 98.320 169.230 103.930 169.270 ;
        RECT 104.320 169.230 110.930 169.270 ;
        RECT 111.320 169.230 120.680 169.270 ;
        RECT 121.070 169.230 128.430 169.270 ;
        RECT 128.820 169.230 133.430 169.270 ;
        RECT 133.820 169.230 138.430 169.270 ;
        RECT 138.820 169.230 139.000 169.270 ;
        RECT 90.750 169.145 139.000 169.230 ;
      LAYER nwell ;
        RECT 81.000 167.295 88.500 168.815 ;
        RECT 90.750 167.295 139.000 168.815 ;
      LAYER pwell ;
        RECT 87.500 162.270 144.750 163.215 ;
        RECT 87.500 162.230 87.680 162.270 ;
        RECT 88.070 162.230 96.930 162.270 ;
        RECT 97.320 162.230 107.680 162.270 ;
        RECT 108.070 162.230 117.680 162.270 ;
        RECT 118.070 162.230 130.180 162.270 ;
        RECT 130.570 162.230 144.250 162.270 ;
        RECT 144.570 162.230 144.750 162.270 ;
        RECT 87.500 162.145 144.750 162.230 ;
      LAYER nwell ;
        RECT 87.500 160.295 144.750 161.815 ;
      LAYER pwell ;
        RECT 22.500 155.750 41.500 157.250 ;
        RECT 22.500 155.250 53.000 155.750 ;
        RECT 10.750 149.750 53.000 155.250 ;
      LAYER nwell ;
        RECT 10.750 144.250 41.500 149.750 ;
        RECT 22.500 142.250 41.500 144.250 ;
      LAYER pwell ;
        RECT 41.500 143.750 53.000 149.750 ;
        RECT 114.745 149.015 114.915 149.205 ;
        RECT 116.180 149.065 116.300 149.175 ;
        RECT 119.805 149.015 119.975 149.205 ;
        RECT 125.325 149.015 125.495 149.205 ;
        RECT 126.300 149.065 126.420 149.175 ;
        RECT 131.765 149.015 131.935 149.205 ;
        RECT 137.285 149.015 137.455 149.205 ;
        RECT 138.665 149.015 138.835 149.205 ;
        RECT 114.605 148.205 115.975 149.015 ;
        RECT 116.445 148.205 120.115 149.015 ;
        RECT 120.125 148.205 125.635 149.015 ;
        RECT 125.655 148.145 126.085 148.930 ;
        RECT 126.565 148.205 132.075 149.015 ;
        RECT 132.085 148.205 137.595 149.015 ;
        RECT 137.605 148.205 138.975 149.015 ;
      LAYER nwell ;
        RECT 114.410 144.985 139.170 147.815 ;
      LAYER pwell ;
        RECT 114.605 143.785 115.975 144.595 ;
        RECT 115.985 143.785 117.355 144.595 ;
        RECT 117.535 143.785 120.575 144.695 ;
        RECT 131.395 144.605 132.985 144.695 ;
        RECT 121.045 143.785 124.715 144.595 ;
        RECT 124.725 143.785 130.235 144.595 ;
        RECT 130.415 143.785 132.985 144.605 ;
        RECT 133.005 143.785 136.045 144.695 ;
        RECT 137.605 143.785 138.975 144.595 ;
        RECT 114.745 143.575 114.915 143.785 ;
        RECT 116.180 143.625 116.300 143.735 ;
        RECT 117.045 143.595 117.215 143.785 ;
        RECT 117.535 143.765 117.680 143.785 ;
        RECT 117.510 143.595 117.680 143.765 ;
        RECT 117.965 143.575 118.135 143.765 ;
        RECT 118.430 143.595 118.600 143.765 ;
        RECT 120.780 143.625 120.900 143.735 ;
        RECT 121.700 143.625 121.820 143.735 ;
        RECT 124.405 143.595 124.575 143.785 ;
        RECT 118.455 143.575 118.600 143.595 ;
        RECT 125.325 143.575 125.495 143.765 ;
        RECT 128.545 143.575 128.715 143.765 ;
        RECT 114.605 142.765 115.975 143.575 ;
        RECT 116.445 142.765 118.275 143.575 ;
        RECT 118.455 142.665 121.495 143.575 ;
        RECT 121.965 142.765 125.635 143.575 ;
        RECT 125.655 142.705 126.085 143.490 ;
        RECT 126.105 142.765 128.855 143.575 ;
        RECT 129.005 143.545 129.175 143.765 ;
        RECT 129.925 143.595 130.095 143.785 ;
        RECT 130.415 143.765 130.555 143.785 ;
        RECT 135.900 143.765 136.045 143.785 ;
        RECT 130.385 143.595 130.555 143.765 ;
        RECT 131.820 143.625 131.940 143.735 ;
        RECT 132.230 143.575 132.400 143.765 ;
        RECT 134.580 143.625 134.700 143.735 ;
        RECT 135.900 143.595 136.070 143.765 ;
        RECT 136.365 143.595 136.535 143.765 ;
        RECT 137.285 143.575 137.455 143.765 ;
        RECT 138.665 143.575 138.835 143.785 ;
        RECT 130.220 143.545 131.615 143.575 ;
        RECT 128.880 142.865 131.615 143.545 ;
        RECT 132.085 142.895 134.360 143.575 ;
        RECT 130.205 142.665 131.615 142.865 ;
        RECT 132.990 142.665 134.360 142.895 ;
        RECT 134.845 142.765 137.595 143.575 ;
        RECT 137.605 142.765 138.975 143.575 ;
        RECT 21.250 111.000 25.250 142.000 ;
        RECT 30.750 111.000 34.750 142.000 ;
        RECT 40.250 111.000 44.250 142.000 ;
      LAYER nwell ;
        RECT 114.410 139.545 139.170 142.375 ;
      LAYER pwell ;
        RECT 114.605 138.345 115.975 139.155 ;
        RECT 115.985 138.345 117.815 139.155 ;
        RECT 117.825 139.025 119.170 139.255 ;
        RECT 117.825 138.345 119.655 139.025 ;
        RECT 119.665 138.345 121.035 139.155 ;
        RECT 121.045 138.345 126.555 139.155 ;
        RECT 126.565 138.345 132.075 139.155 ;
        RECT 132.085 138.345 137.595 139.155 ;
        RECT 137.605 138.345 138.975 139.155 ;
        RECT 114.745 138.135 114.915 138.345 ;
        RECT 117.505 138.325 117.675 138.345 ;
        RECT 117.045 138.135 117.215 138.325 ;
        RECT 117.505 138.155 117.680 138.325 ;
        RECT 119.345 138.155 119.515 138.345 ;
        RECT 120.725 138.155 120.895 138.345 ;
        RECT 117.535 138.135 117.680 138.155 ;
        RECT 121.645 138.135 121.815 138.325 ;
        RECT 125.325 138.135 125.495 138.325 ;
        RECT 126.245 138.295 126.415 138.345 ;
        RECT 126.245 138.185 126.420 138.295 ;
        RECT 126.245 138.155 126.415 138.185 ;
        RECT 131.765 138.135 131.935 138.345 ;
        RECT 134.980 138.135 135.150 138.325 ;
        RECT 135.500 138.185 135.620 138.295 ;
        RECT 137.285 138.135 137.455 138.345 ;
        RECT 138.665 138.135 138.835 138.345 ;
        RECT 114.605 137.325 115.975 138.135 ;
        RECT 115.985 137.325 117.355 138.135 ;
        RECT 117.535 137.225 120.575 138.135 ;
        RECT 120.585 137.325 121.955 138.135 ;
        RECT 121.965 137.325 125.635 138.135 ;
        RECT 125.655 137.265 126.085 138.050 ;
        RECT 126.565 137.325 132.075 138.135 ;
        RECT 132.085 137.225 135.295 138.135 ;
        RECT 135.765 137.325 137.595 138.135 ;
        RECT 137.605 137.325 138.975 138.135 ;
      LAYER nwell ;
        RECT 114.410 134.105 139.170 136.935 ;
      LAYER pwell ;
        RECT 114.605 132.905 115.975 133.715 ;
        RECT 116.905 132.905 122.415 133.715 ;
        RECT 122.425 132.905 127.935 133.715 ;
        RECT 127.945 132.905 133.455 133.715 ;
        RECT 133.495 133.615 134.875 133.815 ;
        RECT 133.495 132.935 136.200 133.615 ;
        RECT 133.495 132.905 134.875 132.935 ;
        RECT 114.745 132.695 114.915 132.905 ;
        RECT 116.585 132.750 116.745 132.860 ;
        RECT 117.505 132.695 117.675 132.885 ;
        RECT 117.970 132.695 118.140 132.885 ;
        RECT 121.645 132.740 121.805 132.850 ;
        RECT 122.105 132.715 122.275 132.905 ;
        RECT 125.325 132.695 125.495 132.885 ;
        RECT 126.705 132.740 126.865 132.850 ;
        RECT 127.625 132.715 127.795 132.905 ;
        RECT 130.385 132.695 130.555 132.885 ;
        RECT 132.680 132.695 132.850 132.885 ;
        RECT 133.145 132.715 133.315 132.905 ;
        RECT 135.905 132.885 136.075 132.935 ;
        RECT 136.225 132.905 137.595 133.715 ;
        RECT 137.605 132.905 138.975 133.715 ;
        RECT 135.900 132.715 136.075 132.885 ;
        RECT 135.900 132.695 136.070 132.715 ;
        RECT 137.285 132.695 137.455 132.905 ;
        RECT 138.665 132.695 138.835 132.905 ;
        RECT 114.605 131.885 115.975 132.695 ;
        RECT 115.985 131.885 117.815 132.695 ;
        RECT 117.825 131.785 121.035 132.695 ;
        RECT 121.965 131.885 125.635 132.695 ;
        RECT 125.655 131.825 126.085 132.610 ;
        RECT 127.025 131.885 130.695 132.695 ;
        RECT 130.720 132.015 132.995 132.695 ;
        RECT 130.720 131.785 132.090 132.015 ;
        RECT 133.005 131.785 136.215 132.695 ;
        RECT 136.225 131.885 137.595 132.695 ;
        RECT 137.605 131.885 138.975 132.695 ;
      LAYER nwell ;
        RECT 114.410 128.665 139.170 131.495 ;
      LAYER pwell ;
        RECT 114.605 127.465 115.975 128.275 ;
        RECT 115.985 127.465 117.355 128.275 ;
        RECT 117.365 127.465 120.575 128.375 ;
        RECT 132.775 128.285 134.365 128.375 ;
        RECT 120.585 127.465 126.095 128.275 ;
        RECT 126.105 127.465 131.615 128.275 ;
        RECT 131.795 127.465 134.365 128.285 ;
        RECT 134.845 127.465 137.595 128.275 ;
        RECT 137.605 127.465 138.975 128.275 ;
        RECT 114.745 127.255 114.915 127.465 ;
        RECT 116.180 127.305 116.300 127.415 ;
        RECT 117.045 127.275 117.215 127.465 ;
        RECT 117.510 127.275 117.680 127.465 ;
        RECT 119.805 127.255 119.975 127.445 ;
        RECT 125.325 127.255 125.495 127.445 ;
        RECT 125.785 127.275 125.955 127.465 ;
        RECT 126.300 127.305 126.420 127.415 ;
        RECT 131.305 127.275 131.475 127.465 ;
        RECT 131.795 127.445 131.935 127.465 ;
        RECT 131.765 127.255 131.935 127.445 ;
        RECT 134.580 127.305 134.700 127.415 ;
        RECT 137.285 127.255 137.455 127.465 ;
        RECT 138.665 127.255 138.835 127.465 ;
        RECT 114.605 126.445 115.975 127.255 ;
        RECT 116.445 126.445 120.115 127.255 ;
        RECT 120.125 126.445 125.635 127.255 ;
        RECT 125.655 126.385 126.085 127.170 ;
        RECT 126.565 126.445 132.075 127.255 ;
        RECT 132.085 126.445 137.595 127.255 ;
        RECT 137.605 126.445 138.975 127.255 ;
      LAYER nwell ;
        RECT 114.410 124.450 139.170 126.055 ;
      LAYER pwell ;
        RECT 76.000 114.500 83.000 119.000 ;
        RECT 88.195 118.695 106.305 123.805 ;
      LAYER nwell ;
        RECT 88.195 109.695 106.305 115.555 ;
      LAYER li1 ;
        RECT 81.750 195.250 137.750 195.750 ;
        RECT 21.625 187.875 24.875 188.125 ;
        RECT 21.625 184.375 21.875 187.875 ;
        RECT 23.165 186.750 23.335 187.250 ;
        RECT 22.280 185.480 22.760 186.520 ;
        RECT 23.030 185.480 23.470 186.520 ;
        RECT 23.740 185.480 24.220 186.520 ;
        RECT 23.165 184.750 23.335 185.250 ;
        RECT 24.625 184.375 24.875 187.875 ;
        RECT 21.625 184.125 24.875 184.375 ;
        RECT 21.625 180.625 21.875 184.125 ;
        RECT 23.165 183.000 23.335 183.500 ;
        RECT 22.280 181.730 22.760 182.770 ;
        RECT 23.030 181.730 23.470 182.770 ;
        RECT 23.740 181.730 24.220 182.770 ;
        RECT 23.165 181.000 23.335 181.500 ;
        RECT 24.625 180.625 24.875 184.125 ;
        RECT 21.625 180.375 24.875 180.625 ;
        RECT 21.625 176.875 21.875 180.375 ;
        RECT 23.165 179.250 23.335 179.750 ;
        RECT 22.280 177.980 22.760 179.020 ;
        RECT 23.030 177.980 23.470 179.020 ;
        RECT 23.740 177.980 24.220 179.020 ;
        RECT 23.165 177.250 23.335 177.750 ;
        RECT 24.625 176.875 24.875 180.375 ;
        RECT 21.625 176.625 24.875 176.875 ;
        RECT 21.625 173.125 21.875 176.625 ;
        RECT 23.165 175.500 23.335 176.000 ;
        RECT 22.280 174.230 22.760 175.270 ;
        RECT 23.030 174.230 23.470 175.270 ;
        RECT 23.740 174.230 24.220 175.270 ;
        RECT 23.165 173.500 23.335 174.000 ;
        RECT 24.625 173.125 24.875 176.625 ;
        RECT 21.625 172.875 24.875 173.125 ;
        RECT 21.625 169.375 21.875 172.875 ;
        RECT 23.165 171.750 23.335 172.250 ;
        RECT 22.280 170.480 22.760 171.520 ;
        RECT 23.030 170.480 23.470 171.520 ;
        RECT 23.740 170.480 24.220 171.520 ;
        RECT 23.165 169.750 23.335 170.250 ;
        RECT 24.625 169.375 24.875 172.875 ;
        RECT 21.625 169.125 24.875 169.375 ;
        RECT 21.625 165.625 21.875 169.125 ;
        RECT 23.165 168.000 23.335 168.500 ;
        RECT 22.280 166.730 22.760 167.770 ;
        RECT 23.030 166.730 23.470 167.770 ;
        RECT 23.740 166.730 24.220 167.770 ;
        RECT 23.165 166.000 23.335 166.500 ;
        RECT 24.625 165.625 24.875 169.125 ;
        RECT 21.625 165.375 24.875 165.625 ;
        RECT 21.625 161.875 21.875 165.375 ;
        RECT 23.165 164.250 23.335 164.750 ;
        RECT 22.280 162.980 22.760 164.020 ;
        RECT 23.030 162.980 23.470 164.020 ;
        RECT 23.740 162.980 24.220 164.020 ;
        RECT 23.165 162.250 23.335 162.750 ;
        RECT 24.625 161.875 24.875 165.375 ;
        RECT 21.625 161.625 24.875 161.875 ;
        RECT 21.625 158.125 21.875 161.625 ;
        RECT 23.165 160.500 23.335 161.000 ;
        RECT 22.280 159.230 22.760 160.270 ;
        RECT 23.030 159.230 23.470 160.270 ;
        RECT 23.740 159.230 24.220 160.270 ;
        RECT 23.165 158.500 23.335 159.000 ;
        RECT 24.625 158.125 24.875 161.625 ;
        RECT 21.625 157.875 24.875 158.125 ;
        RECT 31.125 187.875 34.375 188.125 ;
        RECT 31.125 184.375 31.375 187.875 ;
        RECT 32.665 186.750 32.835 187.250 ;
        RECT 31.780 185.480 32.260 186.520 ;
        RECT 32.530 185.480 32.970 186.520 ;
        RECT 33.240 185.480 33.720 186.520 ;
        RECT 32.665 184.750 32.835 185.250 ;
        RECT 34.125 184.375 34.375 187.875 ;
        RECT 31.125 184.125 34.375 184.375 ;
        RECT 31.125 180.625 31.375 184.125 ;
        RECT 32.665 183.000 32.835 183.500 ;
        RECT 31.780 181.730 32.260 182.770 ;
        RECT 32.530 181.730 32.970 182.770 ;
        RECT 33.240 181.730 33.720 182.770 ;
        RECT 32.665 181.000 32.835 181.500 ;
        RECT 34.125 180.625 34.375 184.125 ;
        RECT 31.125 180.375 34.375 180.625 ;
        RECT 31.125 176.875 31.375 180.375 ;
        RECT 32.665 179.250 32.835 179.750 ;
        RECT 31.780 177.980 32.260 179.020 ;
        RECT 32.530 177.980 32.970 179.020 ;
        RECT 33.240 177.980 33.720 179.020 ;
        RECT 32.665 177.250 32.835 177.750 ;
        RECT 34.125 176.875 34.375 180.375 ;
        RECT 31.125 176.625 34.375 176.875 ;
        RECT 31.125 173.125 31.375 176.625 ;
        RECT 32.665 175.500 32.835 176.000 ;
        RECT 31.780 174.230 32.260 175.270 ;
        RECT 32.530 174.230 32.970 175.270 ;
        RECT 33.240 174.230 33.720 175.270 ;
        RECT 32.665 173.500 32.835 174.000 ;
        RECT 34.125 173.125 34.375 176.625 ;
        RECT 31.125 172.875 34.375 173.125 ;
        RECT 31.125 169.375 31.375 172.875 ;
        RECT 32.665 171.750 32.835 172.250 ;
        RECT 31.780 170.480 32.260 171.520 ;
        RECT 32.530 170.480 32.970 171.520 ;
        RECT 33.240 170.480 33.720 171.520 ;
        RECT 32.665 169.750 32.835 170.250 ;
        RECT 34.125 169.375 34.375 172.875 ;
        RECT 31.125 169.125 34.375 169.375 ;
        RECT 31.125 165.625 31.375 169.125 ;
        RECT 32.665 168.000 32.835 168.500 ;
        RECT 31.780 166.730 32.260 167.770 ;
        RECT 32.530 166.730 32.970 167.770 ;
        RECT 33.240 166.730 33.720 167.770 ;
        RECT 32.665 166.000 32.835 166.500 ;
        RECT 34.125 165.625 34.375 169.125 ;
        RECT 31.125 165.375 34.375 165.625 ;
        RECT 31.125 161.875 31.375 165.375 ;
        RECT 32.665 164.250 32.835 164.750 ;
        RECT 31.780 162.980 32.260 164.020 ;
        RECT 32.530 162.980 32.970 164.020 ;
        RECT 33.240 162.980 33.720 164.020 ;
        RECT 32.665 162.250 32.835 162.750 ;
        RECT 34.125 161.875 34.375 165.375 ;
        RECT 31.125 161.625 34.375 161.875 ;
        RECT 31.125 158.125 31.375 161.625 ;
        RECT 32.665 160.500 32.835 161.000 ;
        RECT 31.780 159.230 32.260 160.270 ;
        RECT 32.530 159.230 32.970 160.270 ;
        RECT 33.240 159.230 33.720 160.270 ;
        RECT 32.665 158.500 32.835 159.000 ;
        RECT 34.125 158.125 34.375 161.625 ;
        RECT 31.125 157.875 34.375 158.125 ;
        RECT 40.625 187.875 43.875 188.125 ;
        RECT 40.625 184.375 40.875 187.875 ;
        RECT 42.165 186.750 42.335 187.250 ;
        RECT 41.280 185.480 41.760 186.520 ;
        RECT 42.030 185.480 42.470 186.520 ;
        RECT 42.740 185.480 43.220 186.520 ;
        RECT 42.165 184.750 42.335 185.250 ;
        RECT 43.625 184.375 43.875 187.875 ;
        RECT 40.625 184.125 43.875 184.375 ;
        RECT 40.625 180.625 40.875 184.125 ;
        RECT 42.165 183.000 42.335 183.500 ;
        RECT 41.280 181.730 41.760 182.770 ;
        RECT 42.030 181.730 42.470 182.770 ;
        RECT 42.740 181.730 43.220 182.770 ;
        RECT 42.165 181.000 42.335 181.500 ;
        RECT 43.625 180.625 43.875 184.125 ;
        RECT 81.750 182.250 82.250 195.250 ;
        RECT 86.000 194.135 133.500 194.385 ;
        RECT 86.180 192.770 86.570 194.135 ;
        RECT 86.930 192.770 87.320 194.135 ;
        RECT 87.870 192.935 88.040 194.135 ;
        RECT 88.210 192.935 88.480 193.425 ;
        RECT 88.750 192.935 88.920 194.135 ;
        RECT 89.350 193.615 90.860 193.965 ;
        RECT 89.590 193.105 89.760 193.425 ;
        RECT 89.310 192.935 89.760 193.105 ;
        RECT 90.090 192.935 90.360 193.425 ;
        RECT 91.030 192.935 91.200 194.135 ;
        RECT 91.370 192.935 91.640 193.425 ;
        RECT 88.210 192.025 88.380 192.935 ;
        RECT 89.310 192.645 89.480 192.935 ;
        RECT 88.550 192.315 89.480 192.645 ;
        RECT 89.650 192.640 89.820 192.645 ;
        RECT 90.090 192.640 90.260 192.935 ;
        RECT 89.650 192.315 90.260 192.640 ;
        RECT 91.370 192.565 91.540 192.935 ;
        RECT 90.430 192.395 91.540 192.565 ;
        RECT 86.180 190.375 86.570 191.965 ;
        RECT 86.930 190.375 87.320 191.965 ;
        RECT 87.870 190.375 88.040 192.025 ;
        RECT 88.210 191.085 88.480 192.025 ;
        RECT 88.750 190.375 88.920 192.025 ;
        RECT 89.310 191.085 89.480 192.315 ;
        RECT 90.090 192.025 90.260 192.315 ;
        RECT 91.370 192.025 91.540 192.395 ;
        RECT 91.710 192.315 91.880 192.645 ;
        RECT 89.750 190.375 89.920 192.025 ;
        RECT 90.090 191.085 90.360 192.025 ;
        RECT 90.090 190.700 90.420 190.870 ;
        RECT 90.750 190.375 90.920 192.025 ;
        RECT 91.370 191.085 91.760 192.025 ;
        RECT 92.050 192.000 92.220 193.815 ;
        RECT 92.680 192.770 93.070 194.135 ;
        RECT 93.430 192.770 93.820 194.135 ;
        RECT 94.370 192.935 94.540 194.135 ;
        RECT 94.710 192.935 94.980 193.425 ;
        RECT 95.250 192.935 95.420 194.135 ;
        RECT 95.850 193.615 97.360 193.965 ;
        RECT 96.090 193.105 96.260 193.425 ;
        RECT 95.810 192.935 96.260 193.105 ;
        RECT 96.590 192.935 96.860 193.425 ;
        RECT 97.530 192.935 97.700 194.135 ;
        RECT 97.870 192.935 98.140 193.425 ;
        RECT 94.710 192.025 94.880 192.935 ;
        RECT 95.810 192.645 95.980 192.935 ;
        RECT 95.050 192.315 95.980 192.645 ;
        RECT 96.150 192.640 96.320 192.645 ;
        RECT 96.590 192.640 96.760 192.935 ;
        RECT 96.150 192.315 96.760 192.640 ;
        RECT 97.870 192.565 98.040 192.935 ;
        RECT 96.930 192.395 98.040 192.565 ;
        RECT 91.930 191.500 92.220 192.000 ;
        RECT 91.350 190.700 91.680 190.870 ;
        RECT 92.050 190.670 92.220 191.500 ;
        RECT 92.680 190.375 93.070 191.965 ;
        RECT 93.430 190.375 93.820 191.965 ;
        RECT 94.370 190.375 94.540 192.025 ;
        RECT 94.710 191.085 94.980 192.025 ;
        RECT 95.250 190.375 95.420 192.025 ;
        RECT 95.810 191.085 95.980 192.315 ;
        RECT 96.590 192.025 96.760 192.315 ;
        RECT 97.870 192.025 98.040 192.395 ;
        RECT 98.210 192.315 98.380 192.645 ;
        RECT 96.250 190.375 96.420 192.025 ;
        RECT 96.590 191.085 96.860 192.025 ;
        RECT 96.590 190.700 96.920 190.870 ;
        RECT 97.250 190.375 97.420 192.025 ;
        RECT 97.870 191.085 98.260 192.025 ;
        RECT 98.550 192.000 98.720 193.815 ;
        RECT 99.180 192.770 99.570 194.135 ;
        RECT 100.085 192.935 100.255 194.135 ;
        RECT 100.525 192.935 100.695 193.425 ;
        RECT 100.965 192.935 101.135 194.135 ;
        RECT 101.585 192.935 101.755 194.135 ;
        RECT 102.025 192.935 102.195 193.425 ;
        RECT 102.465 192.935 102.635 194.135 ;
        RECT 103.085 192.935 103.255 194.135 ;
        RECT 103.525 192.935 103.695 193.425 ;
        RECT 103.965 192.935 104.135 194.135 ;
        RECT 104.680 192.770 105.070 194.135 ;
        RECT 105.620 192.935 105.790 194.135 ;
        RECT 105.960 192.935 106.230 193.425 ;
        RECT 106.500 192.935 106.670 194.135 ;
        RECT 107.100 193.615 108.610 193.965 ;
        RECT 107.340 193.105 107.510 193.425 ;
        RECT 107.060 192.935 107.510 193.105 ;
        RECT 107.840 192.935 108.110 193.425 ;
        RECT 108.780 192.935 108.950 194.135 ;
        RECT 109.120 192.935 109.390 193.425 ;
        RECT 100.365 192.645 101.220 192.725 ;
        RECT 101.865 192.645 102.720 192.725 ;
        RECT 103.365 192.645 104.220 192.725 ;
        RECT 100.365 192.315 101.250 192.645 ;
        RECT 101.865 192.315 102.750 192.645 ;
        RECT 103.365 192.315 104.250 192.645 ;
        RECT 100.365 192.235 101.220 192.315 ;
        RECT 101.865 192.235 102.720 192.315 ;
        RECT 103.365 192.235 104.220 192.315 ;
        RECT 105.960 192.025 106.130 192.935 ;
        RECT 107.060 192.645 107.230 192.935 ;
        RECT 106.300 192.315 107.230 192.645 ;
        RECT 107.400 192.640 107.570 192.645 ;
        RECT 107.840 192.640 108.010 192.935 ;
        RECT 107.400 192.315 108.010 192.640 ;
        RECT 109.120 192.565 109.290 192.935 ;
        RECT 108.180 192.395 109.290 192.565 ;
        RECT 98.430 191.500 98.720 192.000 ;
        RECT 97.850 190.700 98.180 190.870 ;
        RECT 98.550 190.670 98.720 191.500 ;
        RECT 99.180 190.375 99.570 191.965 ;
        RECT 100.085 190.375 100.255 192.025 ;
        RECT 100.525 191.085 100.695 192.025 ;
        RECT 100.965 190.375 101.135 192.025 ;
        RECT 101.585 190.375 101.755 192.025 ;
        RECT 102.025 191.085 102.195 192.025 ;
        RECT 102.465 190.375 102.635 192.025 ;
        RECT 103.085 190.375 103.255 192.025 ;
        RECT 103.525 191.085 103.695 192.025 ;
        RECT 103.965 190.375 104.135 192.025 ;
        RECT 104.680 190.375 105.070 191.965 ;
        RECT 105.620 190.375 105.790 192.025 ;
        RECT 105.960 191.085 106.230 192.025 ;
        RECT 106.500 190.375 106.670 192.025 ;
        RECT 107.060 191.085 107.230 192.315 ;
        RECT 107.840 192.025 108.010 192.315 ;
        RECT 109.120 192.025 109.290 192.395 ;
        RECT 109.460 192.315 109.630 192.645 ;
        RECT 107.500 190.375 107.670 192.025 ;
        RECT 107.840 191.085 108.110 192.025 ;
        RECT 107.840 190.700 108.170 190.870 ;
        RECT 108.500 190.375 108.670 192.025 ;
        RECT 109.120 191.085 109.510 192.025 ;
        RECT 109.800 192.000 109.970 193.815 ;
        RECT 110.370 192.935 110.540 194.135 ;
        RECT 110.710 192.935 110.980 193.425 ;
        RECT 111.250 192.935 111.420 194.135 ;
        RECT 111.850 193.615 113.360 193.965 ;
        RECT 112.090 193.105 112.260 193.425 ;
        RECT 111.810 192.935 112.260 193.105 ;
        RECT 112.590 192.935 112.860 193.425 ;
        RECT 113.530 192.935 113.700 194.135 ;
        RECT 113.870 192.935 114.140 193.425 ;
        RECT 110.710 192.025 110.880 192.935 ;
        RECT 111.810 192.645 111.980 192.935 ;
        RECT 111.050 192.315 111.980 192.645 ;
        RECT 112.150 192.640 112.320 192.645 ;
        RECT 112.590 192.640 112.760 192.935 ;
        RECT 112.150 192.315 112.760 192.640 ;
        RECT 113.870 192.565 114.040 192.935 ;
        RECT 112.930 192.395 114.040 192.565 ;
        RECT 109.680 191.500 109.970 192.000 ;
        RECT 109.100 190.700 109.430 190.870 ;
        RECT 109.800 190.670 109.970 191.500 ;
        RECT 110.370 190.375 110.540 192.025 ;
        RECT 110.710 191.085 110.980 192.025 ;
        RECT 111.250 190.375 111.420 192.025 ;
        RECT 111.810 191.085 111.980 192.315 ;
        RECT 112.590 192.025 112.760 192.315 ;
        RECT 113.870 192.025 114.040 192.395 ;
        RECT 114.210 192.315 114.380 192.645 ;
        RECT 112.250 190.375 112.420 192.025 ;
        RECT 112.590 191.085 112.860 192.025 ;
        RECT 112.590 190.700 112.920 190.870 ;
        RECT 113.250 190.375 113.420 192.025 ;
        RECT 113.870 191.085 114.260 192.025 ;
        RECT 114.550 192.000 114.720 193.815 ;
        RECT 115.180 192.770 115.570 194.135 ;
        RECT 116.085 192.935 116.255 194.135 ;
        RECT 116.525 192.935 116.695 193.425 ;
        RECT 116.965 192.935 117.135 194.135 ;
        RECT 117.680 192.770 118.070 194.135 ;
        RECT 118.430 192.770 118.820 194.135 ;
        RECT 119.370 192.935 119.540 194.135 ;
        RECT 119.710 192.935 119.980 193.425 ;
        RECT 120.250 192.935 120.420 194.135 ;
        RECT 120.850 193.615 122.360 193.965 ;
        RECT 121.090 193.105 121.260 193.425 ;
        RECT 120.810 192.935 121.260 193.105 ;
        RECT 121.590 192.935 121.860 193.425 ;
        RECT 122.530 192.935 122.700 194.135 ;
        RECT 122.870 192.935 123.140 193.425 ;
        RECT 116.365 192.645 117.220 192.725 ;
        RECT 116.365 192.315 117.250 192.645 ;
        RECT 116.365 192.235 117.220 192.315 ;
        RECT 119.710 192.025 119.880 192.935 ;
        RECT 120.810 192.645 120.980 192.935 ;
        RECT 120.050 192.315 120.980 192.645 ;
        RECT 121.150 192.640 121.320 192.645 ;
        RECT 121.590 192.640 121.760 192.935 ;
        RECT 121.150 192.315 121.760 192.640 ;
        RECT 122.870 192.565 123.040 192.935 ;
        RECT 121.930 192.395 123.040 192.565 ;
        RECT 114.430 191.500 114.720 192.000 ;
        RECT 113.850 190.700 114.180 190.870 ;
        RECT 114.550 190.670 114.720 191.500 ;
        RECT 115.180 190.375 115.570 191.965 ;
        RECT 116.085 190.375 116.255 192.025 ;
        RECT 116.525 191.085 116.695 192.025 ;
        RECT 116.965 190.375 117.135 192.025 ;
        RECT 117.680 190.375 118.070 191.965 ;
        RECT 118.430 190.375 118.820 191.965 ;
        RECT 119.370 190.375 119.540 192.025 ;
        RECT 119.710 191.085 119.980 192.025 ;
        RECT 120.250 190.375 120.420 192.025 ;
        RECT 120.810 191.085 120.980 192.315 ;
        RECT 121.590 192.025 121.760 192.315 ;
        RECT 122.870 192.025 123.040 192.395 ;
        RECT 123.210 192.315 123.380 192.645 ;
        RECT 121.250 190.375 121.420 192.025 ;
        RECT 121.590 191.085 121.860 192.025 ;
        RECT 121.590 190.700 121.920 190.870 ;
        RECT 122.250 190.375 122.420 192.025 ;
        RECT 122.870 191.085 123.260 192.025 ;
        RECT 123.550 192.000 123.720 193.815 ;
        RECT 123.930 192.770 124.320 194.135 ;
        RECT 124.680 192.770 125.070 194.135 ;
        RECT 125.430 192.770 125.820 194.135 ;
        RECT 126.370 192.935 126.540 194.135 ;
        RECT 126.710 192.935 126.980 193.425 ;
        RECT 127.250 192.935 127.420 194.135 ;
        RECT 127.850 193.615 129.360 193.965 ;
        RECT 128.090 193.105 128.260 193.425 ;
        RECT 127.810 192.935 128.260 193.105 ;
        RECT 128.590 192.935 128.860 193.425 ;
        RECT 129.530 192.935 129.700 194.135 ;
        RECT 129.870 192.935 130.140 193.425 ;
        RECT 126.710 192.025 126.880 192.935 ;
        RECT 127.810 192.645 127.980 192.935 ;
        RECT 127.050 192.315 127.980 192.645 ;
        RECT 128.150 192.640 128.320 192.645 ;
        RECT 128.590 192.640 128.760 192.935 ;
        RECT 128.150 192.315 128.760 192.640 ;
        RECT 129.870 192.565 130.040 192.935 ;
        RECT 128.930 192.395 130.040 192.565 ;
        RECT 123.430 191.500 123.720 192.000 ;
        RECT 122.850 190.700 123.180 190.870 ;
        RECT 123.550 190.670 123.720 191.500 ;
        RECT 123.930 190.375 124.320 191.965 ;
        RECT 124.680 190.375 125.070 191.965 ;
        RECT 125.430 190.375 125.820 191.965 ;
        RECT 126.370 190.375 126.540 192.025 ;
        RECT 126.710 191.085 126.980 192.025 ;
        RECT 127.250 190.375 127.420 192.025 ;
        RECT 127.810 191.085 127.980 192.315 ;
        RECT 128.590 192.025 128.760 192.315 ;
        RECT 129.870 192.025 130.040 192.395 ;
        RECT 130.210 192.315 130.380 192.645 ;
        RECT 128.250 190.375 128.420 192.025 ;
        RECT 128.590 191.085 128.860 192.025 ;
        RECT 128.590 190.700 128.920 190.870 ;
        RECT 129.250 190.375 129.420 192.025 ;
        RECT 129.870 191.085 130.260 192.025 ;
        RECT 130.550 192.000 130.720 193.815 ;
        RECT 131.180 192.770 131.570 194.135 ;
        RECT 132.085 192.935 132.255 194.135 ;
        RECT 132.525 192.935 132.695 193.425 ;
        RECT 132.965 192.935 133.135 194.135 ;
        RECT 132.365 192.645 133.220 192.725 ;
        RECT 132.365 192.315 133.250 192.645 ;
        RECT 132.365 192.235 133.220 192.315 ;
        RECT 130.430 191.500 130.720 192.000 ;
        RECT 129.850 190.700 130.180 190.870 ;
        RECT 130.550 190.670 130.720 191.500 ;
        RECT 131.180 190.375 131.570 191.965 ;
        RECT 132.085 190.375 132.255 192.025 ;
        RECT 132.525 191.085 132.695 192.025 ;
        RECT 132.965 190.375 133.135 192.025 ;
        RECT 86.000 190.125 133.500 190.375 ;
        RECT 85.500 187.885 133.500 188.135 ;
        RECT 85.870 186.685 86.040 187.885 ;
        RECT 86.210 186.685 86.480 187.175 ;
        RECT 86.750 186.685 86.920 187.885 ;
        RECT 87.350 187.365 88.860 187.715 ;
        RECT 87.590 186.855 87.760 187.175 ;
        RECT 87.310 186.685 87.760 186.855 ;
        RECT 88.090 186.685 88.360 187.175 ;
        RECT 89.030 186.685 89.200 187.885 ;
        RECT 89.370 186.685 89.640 187.175 ;
        RECT 86.210 185.775 86.380 186.685 ;
        RECT 87.310 186.395 87.480 186.685 ;
        RECT 86.550 186.065 87.480 186.395 ;
        RECT 87.650 186.390 87.820 186.395 ;
        RECT 88.090 186.390 88.260 186.685 ;
        RECT 87.650 186.065 88.260 186.390 ;
        RECT 89.370 186.315 89.540 186.685 ;
        RECT 88.430 186.145 89.540 186.315 ;
        RECT 85.870 184.125 86.040 185.775 ;
        RECT 86.210 184.835 86.480 185.775 ;
        RECT 86.750 184.125 86.920 185.775 ;
        RECT 87.310 184.835 87.480 186.065 ;
        RECT 88.090 185.775 88.260 186.065 ;
        RECT 89.370 185.775 89.540 186.145 ;
        RECT 89.710 186.065 89.880 186.395 ;
        RECT 87.750 184.125 87.920 185.775 ;
        RECT 88.090 184.835 88.360 185.775 ;
        RECT 88.090 184.450 88.420 184.620 ;
        RECT 88.750 184.125 88.920 185.775 ;
        RECT 89.370 184.835 89.760 185.775 ;
        RECT 90.050 185.750 90.220 187.565 ;
        RECT 90.890 186.685 91.060 187.885 ;
        RECT 90.830 186.345 91.160 186.515 ;
        RECT 91.330 186.115 91.500 187.175 ;
        RECT 91.770 186.685 91.940 187.885 ;
        RECT 92.430 186.520 92.820 187.885 ;
        RECT 93.390 186.685 93.560 187.885 ;
        RECT 93.330 186.345 93.660 186.515 ;
        RECT 90.810 185.945 91.500 186.115 ;
        RECT 91.670 185.945 92.000 186.160 ;
        RECT 93.830 186.115 94.000 187.175 ;
        RECT 94.270 186.685 94.440 187.885 ;
        RECT 95.085 186.685 95.255 187.885 ;
        RECT 95.525 186.685 95.695 187.175 ;
        RECT 95.965 186.685 96.135 187.885 ;
        RECT 96.870 186.685 97.040 187.885 ;
        RECT 97.210 186.685 97.480 187.175 ;
        RECT 97.750 186.685 97.920 187.885 ;
        RECT 98.350 187.365 99.860 187.715 ;
        RECT 98.590 186.855 98.760 187.175 ;
        RECT 98.310 186.685 98.760 186.855 ;
        RECT 99.090 186.685 99.360 187.175 ;
        RECT 100.030 186.685 100.200 187.885 ;
        RECT 100.370 186.685 100.640 187.175 ;
        RECT 95.365 186.395 96.220 186.475 ;
        RECT 93.310 185.945 94.000 186.115 ;
        RECT 94.170 185.945 94.500 186.160 ;
        RECT 95.365 186.065 96.250 186.395 ;
        RECT 95.365 185.985 96.220 186.065 ;
        RECT 97.210 185.775 97.380 186.685 ;
        RECT 98.310 186.395 98.480 186.685 ;
        RECT 97.550 186.065 98.480 186.395 ;
        RECT 98.650 186.390 98.820 186.395 ;
        RECT 99.090 186.390 99.260 186.685 ;
        RECT 98.650 186.065 99.260 186.390 ;
        RECT 100.370 186.315 100.540 186.685 ;
        RECT 99.430 186.145 100.540 186.315 ;
        RECT 89.930 185.250 90.220 185.750 ;
        RECT 89.350 184.450 89.680 184.620 ;
        RECT 90.050 184.420 90.220 185.250 ;
        RECT 90.890 184.835 91.060 185.775 ;
        RECT 91.730 184.125 91.900 185.775 ;
        RECT 92.430 184.125 92.820 185.715 ;
        RECT 93.390 184.835 93.560 185.775 ;
        RECT 94.230 184.125 94.400 185.775 ;
        RECT 95.085 184.125 95.255 185.775 ;
        RECT 95.525 184.835 95.695 185.775 ;
        RECT 95.965 184.125 96.135 185.775 ;
        RECT 96.870 184.125 97.040 185.775 ;
        RECT 97.210 184.835 97.480 185.775 ;
        RECT 97.750 184.125 97.920 185.775 ;
        RECT 98.310 184.835 98.480 186.065 ;
        RECT 99.090 185.775 99.260 186.065 ;
        RECT 100.370 185.775 100.540 186.145 ;
        RECT 100.710 186.065 100.880 186.395 ;
        RECT 98.750 184.125 98.920 185.775 ;
        RECT 99.090 184.835 99.360 185.775 ;
        RECT 99.090 184.450 99.420 184.620 ;
        RECT 99.750 184.125 99.920 185.775 ;
        RECT 100.370 184.835 100.760 185.775 ;
        RECT 101.050 185.750 101.220 187.565 ;
        RECT 101.870 186.685 102.040 187.885 ;
        RECT 102.210 186.685 102.480 187.175 ;
        RECT 102.750 186.685 102.920 187.885 ;
        RECT 103.350 187.365 104.860 187.715 ;
        RECT 103.590 186.855 103.760 187.175 ;
        RECT 103.310 186.685 103.760 186.855 ;
        RECT 104.090 186.685 104.360 187.175 ;
        RECT 105.030 186.685 105.200 187.885 ;
        RECT 105.370 186.685 105.640 187.175 ;
        RECT 102.210 185.775 102.380 186.685 ;
        RECT 103.310 186.395 103.480 186.685 ;
        RECT 102.550 186.065 103.480 186.395 ;
        RECT 103.650 186.390 103.820 186.395 ;
        RECT 104.090 186.390 104.260 186.685 ;
        RECT 103.650 186.065 104.260 186.390 ;
        RECT 105.370 186.315 105.540 186.685 ;
        RECT 104.430 186.145 105.540 186.315 ;
        RECT 100.930 185.250 101.220 185.750 ;
        RECT 100.350 184.450 100.680 184.620 ;
        RECT 101.050 184.420 101.220 185.250 ;
        RECT 101.870 184.125 102.040 185.775 ;
        RECT 102.210 184.835 102.480 185.775 ;
        RECT 102.750 184.125 102.920 185.775 ;
        RECT 103.310 184.835 103.480 186.065 ;
        RECT 104.090 185.775 104.260 186.065 ;
        RECT 105.370 185.775 105.540 186.145 ;
        RECT 105.710 186.065 105.880 186.395 ;
        RECT 103.750 184.125 103.920 185.775 ;
        RECT 104.090 184.835 104.360 185.775 ;
        RECT 104.090 184.450 104.420 184.620 ;
        RECT 104.750 184.125 104.920 185.775 ;
        RECT 105.370 184.835 105.760 185.775 ;
        RECT 106.050 185.750 106.220 187.565 ;
        RECT 106.890 186.685 107.060 187.885 ;
        RECT 106.830 186.345 107.160 186.515 ;
        RECT 107.330 186.115 107.500 187.175 ;
        RECT 107.770 186.685 107.940 187.885 ;
        RECT 108.430 186.520 108.820 187.885 ;
        RECT 109.390 186.685 109.560 187.885 ;
        RECT 109.330 186.345 109.660 186.515 ;
        RECT 106.810 185.945 107.500 186.115 ;
        RECT 107.670 185.945 108.000 186.160 ;
        RECT 109.830 186.115 110.000 187.175 ;
        RECT 110.270 186.685 110.440 187.885 ;
        RECT 111.085 186.685 111.255 187.885 ;
        RECT 111.525 186.685 111.695 187.175 ;
        RECT 111.965 186.685 112.135 187.885 ;
        RECT 112.870 186.685 113.040 187.885 ;
        RECT 113.210 186.685 113.480 187.175 ;
        RECT 113.750 186.685 113.920 187.885 ;
        RECT 114.350 187.365 115.860 187.715 ;
        RECT 114.590 186.855 114.760 187.175 ;
        RECT 114.310 186.685 114.760 186.855 ;
        RECT 115.090 186.685 115.360 187.175 ;
        RECT 116.030 186.685 116.200 187.885 ;
        RECT 116.370 186.685 116.640 187.175 ;
        RECT 111.365 186.395 112.220 186.475 ;
        RECT 109.310 185.945 110.000 186.115 ;
        RECT 110.170 185.945 110.500 186.160 ;
        RECT 111.365 186.065 112.250 186.395 ;
        RECT 111.365 185.985 112.220 186.065 ;
        RECT 113.210 185.775 113.380 186.685 ;
        RECT 114.310 186.395 114.480 186.685 ;
        RECT 113.550 186.065 114.480 186.395 ;
        RECT 114.650 186.390 114.820 186.395 ;
        RECT 115.090 186.390 115.260 186.685 ;
        RECT 114.650 186.065 115.260 186.390 ;
        RECT 116.370 186.315 116.540 186.685 ;
        RECT 115.430 186.145 116.540 186.315 ;
        RECT 105.930 185.250 106.220 185.750 ;
        RECT 105.350 184.450 105.680 184.620 ;
        RECT 106.050 184.420 106.220 185.250 ;
        RECT 106.890 184.835 107.060 185.775 ;
        RECT 107.730 184.125 107.900 185.775 ;
        RECT 108.430 184.125 108.820 185.715 ;
        RECT 109.390 184.835 109.560 185.775 ;
        RECT 110.230 184.125 110.400 185.775 ;
        RECT 111.085 184.125 111.255 185.775 ;
        RECT 111.525 184.835 111.695 185.775 ;
        RECT 111.965 184.125 112.135 185.775 ;
        RECT 112.870 184.125 113.040 185.775 ;
        RECT 113.210 184.835 113.480 185.775 ;
        RECT 113.750 184.125 113.920 185.775 ;
        RECT 114.310 184.835 114.480 186.065 ;
        RECT 115.090 185.775 115.260 186.065 ;
        RECT 116.370 185.775 116.540 186.145 ;
        RECT 116.710 186.065 116.880 186.395 ;
        RECT 114.750 184.125 114.920 185.775 ;
        RECT 115.090 184.835 115.360 185.775 ;
        RECT 115.090 184.450 115.420 184.620 ;
        RECT 115.750 184.125 115.920 185.775 ;
        RECT 116.370 184.835 116.760 185.775 ;
        RECT 117.050 185.750 117.220 187.565 ;
        RECT 117.870 186.685 118.040 187.885 ;
        RECT 118.210 186.685 118.480 187.175 ;
        RECT 118.750 186.685 118.920 187.885 ;
        RECT 119.350 187.365 120.860 187.715 ;
        RECT 119.590 186.855 119.760 187.175 ;
        RECT 119.310 186.685 119.760 186.855 ;
        RECT 120.090 186.685 120.360 187.175 ;
        RECT 121.030 186.685 121.200 187.885 ;
        RECT 121.370 186.685 121.640 187.175 ;
        RECT 118.210 185.775 118.380 186.685 ;
        RECT 119.310 186.395 119.480 186.685 ;
        RECT 118.550 186.065 119.480 186.395 ;
        RECT 119.650 186.390 119.820 186.395 ;
        RECT 120.090 186.390 120.260 186.685 ;
        RECT 119.650 186.065 120.260 186.390 ;
        RECT 121.370 186.315 121.540 186.685 ;
        RECT 120.430 186.145 121.540 186.315 ;
        RECT 116.930 185.250 117.220 185.750 ;
        RECT 116.350 184.450 116.680 184.620 ;
        RECT 117.050 184.420 117.220 185.250 ;
        RECT 117.870 184.125 118.040 185.775 ;
        RECT 118.210 184.835 118.480 185.775 ;
        RECT 118.750 184.125 118.920 185.775 ;
        RECT 119.310 184.835 119.480 186.065 ;
        RECT 120.090 185.775 120.260 186.065 ;
        RECT 121.370 185.775 121.540 186.145 ;
        RECT 121.710 186.065 121.880 186.395 ;
        RECT 119.750 184.125 119.920 185.775 ;
        RECT 120.090 184.835 120.360 185.775 ;
        RECT 120.090 184.450 120.420 184.620 ;
        RECT 120.750 184.125 120.920 185.775 ;
        RECT 121.370 184.835 121.760 185.775 ;
        RECT 122.050 185.750 122.220 187.565 ;
        RECT 122.890 186.685 123.060 187.885 ;
        RECT 122.830 186.345 123.160 186.515 ;
        RECT 123.330 186.115 123.500 187.175 ;
        RECT 123.770 186.685 123.940 187.885 ;
        RECT 124.430 186.520 124.820 187.885 ;
        RECT 125.390 186.685 125.560 187.885 ;
        RECT 125.330 186.345 125.660 186.515 ;
        RECT 122.810 185.945 123.500 186.115 ;
        RECT 123.670 185.945 124.000 186.160 ;
        RECT 125.830 186.115 126.000 187.175 ;
        RECT 126.270 186.685 126.440 187.885 ;
        RECT 127.085 186.685 127.255 187.885 ;
        RECT 127.525 186.685 127.695 187.175 ;
        RECT 127.965 186.685 128.135 187.885 ;
        RECT 128.870 186.685 129.040 187.885 ;
        RECT 129.210 186.685 129.480 187.175 ;
        RECT 129.750 186.685 129.920 187.885 ;
        RECT 130.350 187.365 131.860 187.715 ;
        RECT 130.590 186.855 130.760 187.175 ;
        RECT 130.310 186.685 130.760 186.855 ;
        RECT 131.090 186.685 131.360 187.175 ;
        RECT 132.030 186.685 132.200 187.885 ;
        RECT 132.370 186.685 132.640 187.175 ;
        RECT 127.365 186.395 128.220 186.475 ;
        RECT 125.310 185.945 126.000 186.115 ;
        RECT 126.170 185.945 126.500 186.160 ;
        RECT 127.365 186.065 128.250 186.395 ;
        RECT 127.365 185.985 128.220 186.065 ;
        RECT 129.210 185.775 129.380 186.685 ;
        RECT 130.310 186.395 130.480 186.685 ;
        RECT 129.550 186.065 130.480 186.395 ;
        RECT 130.650 186.390 130.820 186.395 ;
        RECT 131.090 186.390 131.260 186.685 ;
        RECT 130.650 186.065 131.260 186.390 ;
        RECT 132.370 186.315 132.540 186.685 ;
        RECT 131.430 186.145 132.540 186.315 ;
        RECT 121.930 185.250 122.220 185.750 ;
        RECT 121.350 184.450 121.680 184.620 ;
        RECT 122.050 184.420 122.220 185.250 ;
        RECT 122.890 184.835 123.060 185.775 ;
        RECT 123.730 184.125 123.900 185.775 ;
        RECT 124.430 184.125 124.820 185.715 ;
        RECT 125.390 184.835 125.560 185.775 ;
        RECT 126.230 184.125 126.400 185.775 ;
        RECT 127.085 184.125 127.255 185.775 ;
        RECT 127.525 184.835 127.695 185.775 ;
        RECT 127.965 184.125 128.135 185.775 ;
        RECT 128.870 184.125 129.040 185.775 ;
        RECT 129.210 184.835 129.480 185.775 ;
        RECT 129.750 184.125 129.920 185.775 ;
        RECT 130.310 184.835 130.480 186.065 ;
        RECT 131.090 185.775 131.260 186.065 ;
        RECT 132.370 185.775 132.540 186.145 ;
        RECT 132.710 186.065 132.880 186.395 ;
        RECT 130.750 184.125 130.920 185.775 ;
        RECT 131.090 184.835 131.360 185.775 ;
        RECT 131.090 184.450 131.420 184.620 ;
        RECT 131.750 184.125 131.920 185.775 ;
        RECT 132.370 184.835 132.760 185.775 ;
        RECT 133.050 185.750 133.220 187.565 ;
        RECT 132.930 185.250 133.220 185.750 ;
        RECT 132.350 184.450 132.680 184.620 ;
        RECT 133.050 184.420 133.220 185.250 ;
        RECT 85.500 183.875 133.500 184.125 ;
        RECT 137.250 182.250 137.750 195.250 ;
        RECT 81.750 181.750 137.750 182.250 ;
        RECT 40.625 180.375 43.875 180.625 ;
        RECT 40.625 176.875 40.875 180.375 ;
        RECT 42.165 179.250 42.335 179.750 ;
        RECT 41.280 177.980 41.760 179.020 ;
        RECT 42.030 177.980 42.470 179.020 ;
        RECT 42.740 177.980 43.220 179.020 ;
        RECT 42.165 177.250 42.335 177.750 ;
        RECT 43.625 176.875 43.875 180.375 ;
        RECT 40.625 176.625 43.875 176.875 ;
        RECT 40.625 173.125 40.875 176.625 ;
        RECT 42.165 175.500 42.335 176.000 ;
        RECT 41.280 174.230 41.760 175.270 ;
        RECT 42.030 174.230 42.470 175.270 ;
        RECT 42.740 174.230 43.220 175.270 ;
        RECT 42.165 173.500 42.335 174.000 ;
        RECT 43.625 173.125 43.875 176.625 ;
        RECT 40.625 172.875 43.875 173.125 ;
        RECT 40.625 169.375 40.875 172.875 ;
        RECT 42.165 171.750 42.335 172.250 ;
        RECT 41.280 170.480 41.760 171.520 ;
        RECT 42.030 170.480 42.470 171.520 ;
        RECT 42.740 170.480 43.220 171.520 ;
        RECT 42.165 169.750 42.335 170.250 ;
        RECT 43.625 169.375 43.875 172.875 ;
        RECT 40.625 169.125 43.875 169.375 ;
        RECT 40.625 165.625 40.875 169.125 ;
        RECT 42.165 168.000 42.335 168.500 ;
        RECT 41.280 166.730 41.760 167.770 ;
        RECT 42.030 166.730 42.470 167.770 ;
        RECT 42.740 166.730 43.220 167.770 ;
        RECT 42.165 166.000 42.335 166.500 ;
        RECT 43.625 165.625 43.875 169.125 ;
        RECT 40.625 165.375 43.875 165.625 ;
        RECT 40.625 161.875 40.875 165.375 ;
        RECT 42.165 164.250 42.335 164.750 ;
        RECT 41.280 162.980 41.760 164.020 ;
        RECT 42.030 162.980 42.470 164.020 ;
        RECT 42.740 162.980 43.220 164.020 ;
        RECT 42.165 162.250 42.335 162.750 ;
        RECT 43.625 161.875 43.875 165.375 ;
        RECT 40.625 161.625 43.875 161.875 ;
        RECT 40.625 158.125 40.875 161.625 ;
        RECT 42.165 160.500 42.335 161.000 ;
        RECT 41.280 159.230 41.760 160.270 ;
        RECT 42.030 159.230 42.470 160.270 ;
        RECT 42.740 159.230 43.220 160.270 ;
        RECT 42.165 158.500 42.335 159.000 ;
        RECT 43.625 158.125 43.875 161.625 ;
        RECT 40.625 157.875 43.875 158.125 ;
        RECT 77.500 180.750 145.750 181.250 ;
        RECT 22.875 156.625 41.125 156.875 ;
        RECT 11.125 154.625 22.375 154.875 ;
        RECT 11.125 150.375 11.375 154.625 ;
        RECT 11.715 152.155 11.885 154.195 ;
        RECT 12.155 152.155 12.325 154.195 ;
        RECT 12.595 152.155 12.765 154.195 ;
        RECT 13.035 152.155 13.205 154.195 ;
        RECT 13.475 152.155 13.645 154.195 ;
        RECT 13.915 152.155 14.085 154.195 ;
        RECT 14.355 152.155 14.525 154.195 ;
        RECT 14.795 152.155 14.965 154.195 ;
        RECT 15.235 152.155 15.405 154.195 ;
        RECT 15.675 152.155 15.845 154.195 ;
        RECT 16.115 152.155 16.285 154.195 ;
        RECT 13.915 150.750 14.085 151.250 ;
        RECT 16.625 150.375 16.875 154.625 ;
        RECT 17.215 152.155 17.385 154.195 ;
        RECT 17.655 152.155 17.825 154.195 ;
        RECT 18.095 152.155 18.265 154.195 ;
        RECT 18.535 152.155 18.705 154.195 ;
        RECT 18.975 152.155 19.145 154.195 ;
        RECT 19.415 152.155 19.585 154.195 ;
        RECT 19.855 152.155 20.025 154.195 ;
        RECT 20.295 152.155 20.465 154.195 ;
        RECT 20.735 152.155 20.905 154.195 ;
        RECT 21.175 152.155 21.345 154.195 ;
        RECT 21.615 152.155 21.785 154.195 ;
        RECT 19.415 150.750 19.585 151.250 ;
        RECT 22.125 150.375 22.375 154.625 ;
        RECT 11.125 150.125 22.375 150.375 ;
        RECT 22.875 150.375 23.125 156.625 ;
        RECT 23.615 152.230 23.785 156.270 ;
        RECT 24.075 152.230 24.245 156.270 ;
        RECT 24.535 152.230 24.705 156.270 ;
        RECT 24.995 152.230 25.165 156.270 ;
        RECT 25.455 152.230 25.625 156.270 ;
        RECT 25.915 152.230 26.085 156.270 ;
        RECT 26.375 152.230 26.545 156.270 ;
        RECT 26.835 152.230 27.005 156.270 ;
        RECT 27.295 152.230 27.465 156.270 ;
        RECT 27.755 152.230 27.925 156.270 ;
        RECT 28.215 152.230 28.385 156.270 ;
        RECT 25.915 150.750 26.085 151.250 ;
        RECT 28.875 150.375 29.125 156.625 ;
        RECT 29.615 152.230 29.785 156.270 ;
        RECT 30.075 152.230 30.245 156.270 ;
        RECT 30.535 152.230 30.705 156.270 ;
        RECT 30.995 152.230 31.165 156.270 ;
        RECT 31.455 152.230 31.625 156.270 ;
        RECT 31.915 152.230 32.085 156.270 ;
        RECT 32.375 152.230 32.545 156.270 ;
        RECT 32.835 152.230 33.005 156.270 ;
        RECT 33.295 152.230 33.465 156.270 ;
        RECT 33.755 152.230 33.925 156.270 ;
        RECT 34.215 152.230 34.385 156.270 ;
        RECT 31.915 150.750 32.085 151.250 ;
        RECT 34.875 150.375 35.125 156.625 ;
        RECT 35.615 152.230 35.785 156.270 ;
        RECT 36.075 152.230 36.245 156.270 ;
        RECT 36.535 152.230 36.705 156.270 ;
        RECT 36.995 152.230 37.165 156.270 ;
        RECT 37.455 152.230 37.625 156.270 ;
        RECT 37.915 152.230 38.085 156.270 ;
        RECT 38.375 152.230 38.545 156.270 ;
        RECT 38.835 152.230 39.005 156.270 ;
        RECT 39.295 152.230 39.465 156.270 ;
        RECT 39.755 152.230 39.925 156.270 ;
        RECT 40.215 152.230 40.385 156.270 ;
        RECT 37.915 150.750 38.085 151.250 ;
        RECT 40.875 150.375 41.125 156.625 ;
        RECT 77.500 156.750 78.000 180.750 ;
        RECT 81.000 177.635 139.250 177.885 ;
        RECT 81.335 176.435 81.505 177.635 ;
        RECT 81.775 176.435 81.945 176.925 ;
        RECT 82.215 176.435 82.385 177.635 ;
        RECT 82.930 176.270 83.320 177.635 ;
        RECT 83.835 176.435 84.005 177.635 ;
        RECT 84.275 176.435 84.445 176.925 ;
        RECT 84.715 176.435 84.885 177.635 ;
        RECT 85.335 176.435 85.505 177.635 ;
        RECT 85.775 176.435 85.945 176.925 ;
        RECT 86.215 176.435 86.385 177.635 ;
        RECT 87.000 176.435 87.170 176.925 ;
        RECT 87.840 176.435 88.010 177.635 ;
        RECT 88.585 176.435 88.755 177.635 ;
        RECT 89.025 176.435 89.195 176.925 ;
        RECT 89.465 176.435 89.635 177.635 ;
        RECT 90.180 176.270 90.570 177.635 ;
        RECT 81.615 176.145 82.470 176.225 ;
        RECT 84.115 176.145 84.970 176.225 ;
        RECT 85.615 176.145 86.470 176.225 ;
        RECT 81.615 175.815 82.500 176.145 ;
        RECT 84.115 175.815 85.000 176.145 ;
        RECT 85.615 175.815 86.500 176.145 ;
        RECT 87.600 176.095 88.190 176.265 ;
        RECT 88.865 176.145 89.720 176.225 ;
        RECT 81.615 175.735 82.470 175.815 ;
        RECT 84.115 175.735 84.970 175.815 ;
        RECT 85.615 175.735 86.470 175.815 ;
        RECT 87.120 175.695 88.185 175.925 ;
        RECT 88.865 175.815 89.750 176.145 ;
        RECT 88.865 175.735 89.720 175.815 ;
        RECT 81.335 173.875 81.505 175.525 ;
        RECT 81.775 174.585 81.945 175.525 ;
        RECT 82.215 173.875 82.385 175.525 ;
        RECT 82.930 173.875 83.320 175.465 ;
        RECT 83.835 173.875 84.005 175.525 ;
        RECT 84.275 174.585 84.445 175.525 ;
        RECT 84.715 173.875 84.885 175.525 ;
        RECT 85.335 173.875 85.505 175.525 ;
        RECT 85.775 174.585 85.945 175.525 ;
        RECT 86.215 173.875 86.385 175.525 ;
        RECT 86.960 173.875 87.130 175.525 ;
        RECT 87.400 174.585 87.570 175.525 ;
        RECT 87.840 173.875 88.010 175.525 ;
        RECT 88.585 173.875 88.755 175.525 ;
        RECT 89.025 174.585 89.195 175.525 ;
        RECT 89.465 173.875 89.635 175.525 ;
        RECT 90.180 173.875 90.570 175.465 ;
        RECT 91.160 175.270 91.330 177.360 ;
        RECT 91.510 176.435 91.680 176.925 ;
        RECT 91.950 176.435 92.120 177.635 ;
        RECT 92.290 177.160 92.620 177.465 ;
        RECT 93.440 177.095 93.920 177.265 ;
        RECT 94.090 177.160 94.420 177.465 ;
        RECT 91.500 175.935 91.670 176.265 ;
        RECT 92.290 176.250 92.460 176.685 ;
        RECT 92.710 176.515 93.040 176.845 ;
        RECT 93.350 176.435 93.580 176.925 ;
        RECT 91.870 176.080 93.200 176.250 ;
        RECT 91.530 174.370 91.700 175.230 ;
        RECT 91.870 174.585 92.040 176.080 ;
        RECT 93.410 175.910 93.580 176.435 ;
        RECT 93.750 176.080 93.920 177.095 ;
        RECT 94.250 176.265 94.420 176.685 ;
        RECT 94.590 176.435 94.760 177.635 ;
        RECT 95.030 176.435 95.200 176.925 ;
        RECT 95.470 176.435 95.640 177.635 ;
        RECT 96.180 176.270 96.570 177.635 ;
        RECT 97.115 176.435 97.285 177.635 ;
        RECT 97.555 176.435 97.725 176.925 ;
        RECT 97.995 176.435 98.165 177.635 ;
        RECT 99.025 176.435 99.195 177.635 ;
        RECT 99.465 176.435 99.695 176.925 ;
        RECT 99.905 176.435 100.075 177.635 ;
        RECT 100.245 177.295 100.575 177.465 ;
        RECT 100.405 176.790 100.575 177.295 ;
        RECT 100.865 177.095 101.195 177.330 ;
        RECT 94.250 176.095 94.640 176.265 ;
        RECT 97.030 176.145 97.885 176.225 ;
        RECT 92.370 175.740 92.980 175.910 ;
        RECT 93.150 175.740 93.580 175.910 ;
        RECT 92.370 174.540 92.540 175.740 ;
        RECT 91.530 174.200 92.250 174.370 ;
        RECT 92.710 173.875 92.880 175.525 ;
        RECT 93.150 174.585 93.320 175.740 ;
        RECT 94.250 175.525 94.420 176.095 ;
        RECT 94.630 175.740 95.180 175.910 ;
        RECT 97.000 175.815 97.885 176.145 ;
        RECT 99.170 175.865 99.350 176.265 ;
        RECT 97.030 175.735 97.885 175.815 ;
        RECT 98.810 175.695 99.350 175.865 ;
        RECT 99.520 175.525 99.695 176.435 ;
        RECT 99.865 175.695 100.575 176.065 ;
        RECT 93.050 174.045 93.380 174.340 ;
        RECT 93.590 173.875 93.760 175.525 ;
        RECT 94.030 174.585 94.420 175.525 ;
        RECT 93.930 174.200 94.260 174.370 ;
        RECT 94.590 173.875 94.760 175.525 ;
        RECT 95.030 174.585 95.200 175.525 ;
        RECT 95.470 173.875 95.640 175.525 ;
        RECT 96.180 173.875 96.570 175.465 ;
        RECT 97.115 173.875 97.285 175.525 ;
        RECT 97.555 174.585 97.725 175.525 ;
        RECT 97.995 173.875 98.165 175.525 ;
        RECT 98.985 173.875 99.155 175.525 ;
        RECT 99.425 174.585 99.695 175.525 ;
        RECT 99.865 173.875 100.035 175.525 ;
        RECT 100.305 174.540 100.475 175.525 ;
        RECT 100.745 174.585 101.015 176.925 ;
        RECT 101.585 176.435 101.755 177.635 ;
        RECT 101.375 175.740 101.855 176.265 ;
        RECT 101.185 174.540 101.355 175.525 ;
        RECT 100.205 174.045 100.535 174.340 ;
        RECT 101.025 174.215 101.195 174.340 ;
        RECT 100.945 174.045 101.275 174.215 ;
        RECT 101.625 173.875 101.795 175.525 ;
        RECT 102.025 174.585 102.295 176.925 ;
        RECT 102.465 176.435 102.635 177.635 ;
        RECT 103.180 176.270 103.570 177.635 ;
        RECT 102.505 173.875 102.675 175.525 ;
        RECT 103.180 173.875 103.570 175.465 ;
        RECT 104.160 175.270 104.330 177.360 ;
        RECT 104.510 176.435 104.680 176.925 ;
        RECT 104.950 176.435 105.120 177.635 ;
        RECT 105.290 177.160 105.620 177.465 ;
        RECT 106.440 177.095 106.920 177.265 ;
        RECT 107.090 177.160 107.420 177.465 ;
        RECT 104.500 175.935 104.670 176.265 ;
        RECT 105.290 176.250 105.460 176.685 ;
        RECT 105.710 176.515 106.040 176.845 ;
        RECT 106.350 176.435 106.580 176.925 ;
        RECT 104.870 176.080 106.200 176.250 ;
        RECT 104.530 174.370 104.700 175.230 ;
        RECT 104.870 174.585 105.040 176.080 ;
        RECT 106.410 175.910 106.580 176.435 ;
        RECT 106.750 176.080 106.920 177.095 ;
        RECT 107.250 176.265 107.420 176.685 ;
        RECT 107.590 176.435 107.760 177.635 ;
        RECT 108.030 176.435 108.200 176.925 ;
        RECT 108.470 176.435 108.640 177.635 ;
        RECT 109.180 176.270 109.570 177.635 ;
        RECT 110.115 176.435 110.285 177.635 ;
        RECT 110.555 176.435 110.725 176.925 ;
        RECT 110.995 176.435 111.165 177.635 ;
        RECT 112.025 176.435 112.195 177.635 ;
        RECT 112.465 176.435 112.695 176.925 ;
        RECT 112.905 176.435 113.075 177.635 ;
        RECT 113.245 177.295 113.575 177.465 ;
        RECT 113.405 176.790 113.575 177.295 ;
        RECT 113.865 177.095 114.195 177.330 ;
        RECT 107.250 176.095 107.640 176.265 ;
        RECT 110.030 176.145 110.885 176.225 ;
        RECT 105.370 175.740 105.980 175.910 ;
        RECT 106.150 175.740 106.580 175.910 ;
        RECT 105.370 174.540 105.540 175.740 ;
        RECT 104.530 174.200 105.250 174.370 ;
        RECT 105.710 173.875 105.880 175.525 ;
        RECT 106.150 174.585 106.320 175.740 ;
        RECT 107.250 175.525 107.420 176.095 ;
        RECT 107.630 175.740 108.180 175.910 ;
        RECT 110.000 175.815 110.885 176.145 ;
        RECT 112.170 175.865 112.350 176.265 ;
        RECT 110.030 175.735 110.885 175.815 ;
        RECT 111.810 175.695 112.350 175.865 ;
        RECT 112.520 175.525 112.695 176.435 ;
        RECT 112.865 175.695 113.575 176.065 ;
        RECT 106.050 174.045 106.380 174.340 ;
        RECT 106.590 173.875 106.760 175.525 ;
        RECT 107.030 174.585 107.420 175.525 ;
        RECT 106.930 174.200 107.260 174.370 ;
        RECT 107.590 173.875 107.760 175.525 ;
        RECT 108.030 174.585 108.200 175.525 ;
        RECT 108.470 173.875 108.640 175.525 ;
        RECT 109.180 173.875 109.570 175.465 ;
        RECT 110.115 173.875 110.285 175.525 ;
        RECT 110.555 174.585 110.725 175.525 ;
        RECT 110.995 173.875 111.165 175.525 ;
        RECT 111.985 173.875 112.155 175.525 ;
        RECT 112.425 174.585 112.695 175.525 ;
        RECT 112.865 173.875 113.035 175.525 ;
        RECT 113.305 174.540 113.475 175.525 ;
        RECT 113.745 174.585 114.015 176.925 ;
        RECT 114.585 176.435 114.755 177.635 ;
        RECT 114.375 175.740 114.855 176.265 ;
        RECT 114.185 174.540 114.355 175.525 ;
        RECT 113.205 174.045 113.535 174.340 ;
        RECT 114.025 174.215 114.195 174.340 ;
        RECT 113.945 174.045 114.275 174.215 ;
        RECT 114.625 173.875 114.795 175.525 ;
        RECT 115.025 174.585 115.295 176.925 ;
        RECT 115.465 176.435 115.635 177.635 ;
        RECT 116.180 176.270 116.570 177.635 ;
        RECT 117.080 177.295 118.320 177.465 ;
        RECT 118.570 177.295 118.990 177.465 ;
        RECT 115.505 173.875 115.675 175.525 ;
        RECT 116.180 173.875 116.570 175.465 ;
        RECT 117.080 174.520 117.250 177.295 ;
        RECT 117.540 176.955 118.400 177.125 ;
        RECT 117.540 176.435 117.710 176.955 ;
        RECT 118.420 176.265 118.590 176.730 ;
        RECT 118.820 176.435 118.990 177.295 ;
        RECT 119.180 176.435 119.350 177.635 ;
        RECT 119.620 176.435 119.790 176.925 ;
        RECT 120.060 176.435 120.230 177.635 ;
        RECT 120.680 176.270 121.070 177.635 ;
        RECT 121.615 176.435 121.785 177.635 ;
        RECT 122.055 176.435 122.225 176.925 ;
        RECT 122.495 176.435 122.665 177.635 ;
        RECT 123.365 176.435 123.535 177.635 ;
        RECT 123.805 176.435 123.975 176.925 ;
        RECT 124.245 176.435 124.415 177.635 ;
        RECT 125.115 176.435 125.285 177.635 ;
        RECT 125.555 176.435 125.725 176.925 ;
        RECT 125.995 176.435 126.165 177.635 ;
        RECT 126.865 176.435 127.035 177.635 ;
        RECT 127.305 176.435 127.475 176.925 ;
        RECT 127.745 176.435 127.915 177.635 ;
        RECT 128.430 176.270 128.820 177.635 ;
        RECT 129.365 176.435 129.535 177.635 ;
        RECT 129.805 176.435 129.975 176.925 ;
        RECT 130.245 176.435 130.415 177.635 ;
        RECT 131.170 176.435 131.840 176.925 ;
        RECT 132.010 176.435 132.180 177.635 ;
        RECT 132.450 176.435 132.620 176.925 ;
        RECT 132.890 176.435 133.060 177.635 ;
        RECT 117.660 176.035 117.990 176.205 ;
        RECT 118.420 176.095 119.230 176.265 ;
        RECT 121.530 176.145 122.385 176.225 ;
        RECT 123.280 176.145 124.135 176.225 ;
        RECT 125.030 176.145 125.885 176.225 ;
        RECT 126.780 176.145 127.635 176.225 ;
        RECT 129.280 176.145 130.135 176.225 ;
        RECT 118.900 176.035 119.230 176.095 ;
        RECT 119.380 175.865 120.000 175.910 ;
        RECT 117.860 175.695 120.000 175.865 ;
        RECT 121.500 175.815 122.385 176.145 ;
        RECT 123.250 175.815 124.135 176.145 ;
        RECT 125.000 175.815 125.885 176.145 ;
        RECT 126.750 175.815 127.635 176.145 ;
        RECT 129.250 175.815 130.135 176.145 ;
        RECT 131.060 176.095 132.060 176.265 ;
        RECT 131.730 176.075 132.060 176.095 ;
        RECT 121.530 175.735 122.385 175.815 ;
        RECT 123.280 175.735 124.135 175.815 ;
        RECT 125.030 175.735 125.885 175.815 ;
        RECT 126.780 175.735 127.635 175.815 ;
        RECT 129.280 175.735 130.135 175.815 ;
        RECT 131.000 175.695 131.540 175.910 ;
        RECT 132.240 175.905 132.570 175.950 ;
        RECT 131.880 175.735 132.570 175.905 ;
        RECT 117.420 173.875 117.590 175.525 ;
        RECT 117.860 174.585 118.030 175.695 ;
        RECT 117.800 174.045 118.130 174.340 ;
        RECT 118.300 173.875 118.470 175.525 ;
        RECT 118.740 174.585 118.910 175.695 ;
        RECT 118.640 174.045 118.970 174.340 ;
        RECT 119.180 173.875 119.350 175.525 ;
        RECT 119.620 174.585 119.790 175.525 ;
        RECT 120.060 173.875 120.230 175.525 ;
        RECT 120.680 173.875 121.070 175.465 ;
        RECT 121.615 173.875 121.785 175.525 ;
        RECT 122.055 174.585 122.225 175.525 ;
        RECT 122.495 173.875 122.665 175.525 ;
        RECT 123.365 173.875 123.535 175.525 ;
        RECT 123.805 174.585 123.975 175.525 ;
        RECT 124.245 173.875 124.415 175.525 ;
        RECT 125.115 173.875 125.285 175.525 ;
        RECT 125.555 174.585 125.725 175.525 ;
        RECT 125.995 173.875 126.165 175.525 ;
        RECT 126.865 173.875 127.035 175.525 ;
        RECT 127.305 174.585 127.475 175.525 ;
        RECT 127.745 173.875 127.915 175.525 ;
        RECT 128.430 173.875 128.820 175.465 ;
        RECT 129.365 173.875 129.535 175.525 ;
        RECT 129.805 174.585 129.975 175.525 ;
        RECT 130.245 173.875 130.415 175.525 ;
        RECT 131.130 173.875 131.300 175.525 ;
        RECT 131.570 174.585 131.840 175.525 ;
        RECT 132.010 173.875 132.180 175.525 ;
        RECT 132.450 174.585 132.620 175.525 ;
        RECT 132.890 173.875 133.060 175.525 ;
        RECT 133.660 175.270 133.830 177.360 ;
        RECT 134.010 176.435 134.180 176.925 ;
        RECT 134.450 176.435 134.620 177.635 ;
        RECT 134.790 177.160 135.120 177.465 ;
        RECT 135.940 177.095 136.420 177.265 ;
        RECT 136.590 177.160 136.920 177.465 ;
        RECT 134.000 175.935 134.170 176.265 ;
        RECT 134.790 176.250 134.960 176.685 ;
        RECT 135.210 176.515 135.540 176.845 ;
        RECT 135.850 176.435 136.080 176.925 ;
        RECT 134.370 176.080 135.700 176.250 ;
        RECT 134.030 174.370 134.200 175.230 ;
        RECT 134.370 174.585 134.540 176.080 ;
        RECT 135.910 175.910 136.080 176.435 ;
        RECT 136.250 176.080 136.420 177.095 ;
        RECT 136.750 176.265 136.920 176.685 ;
        RECT 137.090 176.435 137.260 177.635 ;
        RECT 137.530 176.435 137.700 176.925 ;
        RECT 137.970 176.435 138.140 177.635 ;
        RECT 138.680 176.270 139.070 177.635 ;
        RECT 136.750 176.095 137.140 176.265 ;
        RECT 134.870 175.740 135.480 175.910 ;
        RECT 135.650 175.740 136.080 175.910 ;
        RECT 134.870 174.540 135.040 175.740 ;
        RECT 134.030 174.200 134.750 174.370 ;
        RECT 135.210 173.875 135.380 175.525 ;
        RECT 135.650 174.585 135.820 175.740 ;
        RECT 136.750 175.525 136.920 176.095 ;
        RECT 137.130 175.740 137.680 175.910 ;
        RECT 135.550 174.045 135.880 174.340 ;
        RECT 136.090 173.875 136.260 175.525 ;
        RECT 136.530 174.585 136.920 175.525 ;
        RECT 136.430 174.200 136.760 174.370 ;
        RECT 137.090 173.875 137.260 175.525 ;
        RECT 137.530 174.585 137.700 175.525 ;
        RECT 137.970 173.875 138.140 175.525 ;
        RECT 138.680 173.875 139.070 175.465 ;
        RECT 81.000 173.625 139.250 173.875 ;
        RECT 81.000 170.635 88.500 170.885 ;
        RECT 90.750 170.635 139.000 170.885 ;
        RECT 81.335 169.435 81.505 170.635 ;
        RECT 81.775 169.435 81.945 169.925 ;
        RECT 82.215 169.435 82.385 170.635 ;
        RECT 82.930 169.270 83.320 170.635 ;
        RECT 83.835 169.435 84.005 170.635 ;
        RECT 84.275 169.435 84.445 169.925 ;
        RECT 84.715 169.435 84.885 170.635 ;
        RECT 85.335 169.435 85.505 170.635 ;
        RECT 85.775 169.435 85.945 169.925 ;
        RECT 86.215 169.435 86.385 170.635 ;
        RECT 87.000 169.435 87.170 169.925 ;
        RECT 87.840 169.435 88.010 170.635 ;
        RECT 90.930 169.270 91.320 170.635 ;
        RECT 91.865 169.435 92.035 170.635 ;
        RECT 81.615 169.145 82.470 169.225 ;
        RECT 84.115 169.145 84.970 169.225 ;
        RECT 85.615 169.145 86.470 169.225 ;
        RECT 81.615 168.815 82.500 169.145 ;
        RECT 84.115 168.815 85.000 169.145 ;
        RECT 85.615 168.815 86.500 169.145 ;
        RECT 87.600 169.095 88.190 169.265 ;
        RECT 81.615 168.735 82.470 168.815 ;
        RECT 84.115 168.735 84.970 168.815 ;
        RECT 85.615 168.735 86.470 168.815 ;
        RECT 87.120 168.695 88.185 168.925 ;
        RECT 81.335 166.875 81.505 168.525 ;
        RECT 81.775 167.585 81.945 168.525 ;
        RECT 82.215 166.875 82.385 168.525 ;
        RECT 82.930 166.875 83.320 168.465 ;
        RECT 83.835 166.875 84.005 168.525 ;
        RECT 84.275 167.585 84.445 168.525 ;
        RECT 84.715 166.875 84.885 168.525 ;
        RECT 85.335 166.875 85.505 168.525 ;
        RECT 85.775 167.585 85.945 168.525 ;
        RECT 86.215 166.875 86.385 168.525 ;
        RECT 86.960 166.875 87.130 168.525 ;
        RECT 87.400 167.585 87.570 168.525 ;
        RECT 87.840 166.875 88.010 168.525 ;
        RECT 90.930 166.875 91.320 168.465 ;
        RECT 91.825 166.875 91.995 168.525 ;
        RECT 92.205 167.585 92.475 169.925 ;
        RECT 92.745 169.435 92.915 170.635 ;
        RECT 93.305 170.095 93.635 170.330 ;
        RECT 93.925 170.295 94.255 170.465 ;
        RECT 92.645 168.740 93.125 169.265 ;
        RECT 92.705 166.875 92.875 168.525 ;
        RECT 93.145 167.540 93.315 168.525 ;
        RECT 93.485 167.585 93.755 169.925 ;
        RECT 93.925 169.790 94.095 170.295 ;
        RECT 94.425 169.435 94.595 170.635 ;
        RECT 94.805 169.435 95.035 169.925 ;
        RECT 95.305 169.435 95.475 170.635 ;
        RECT 96.335 169.435 96.505 170.635 ;
        RECT 96.775 169.435 96.945 169.925 ;
        RECT 97.215 169.435 97.385 170.635 ;
        RECT 93.925 168.695 94.635 169.065 ;
        RECT 94.805 168.525 94.980 169.435 ;
        RECT 97.930 169.270 98.320 170.635 ;
        RECT 98.860 169.435 99.030 170.635 ;
        RECT 99.300 169.435 99.470 169.925 ;
        RECT 99.740 169.435 99.910 170.635 ;
        RECT 100.080 170.160 100.410 170.465 ;
        RECT 100.580 170.095 101.060 170.265 ;
        RECT 101.880 170.160 102.210 170.465 ;
        RECT 100.080 169.265 100.250 169.685 ;
        RECT 95.150 168.865 95.330 169.265 ;
        RECT 96.615 169.145 97.470 169.225 ;
        RECT 95.150 168.695 95.690 168.865 ;
        RECT 96.615 168.815 97.500 169.145 ;
        RECT 99.860 169.095 100.250 169.265 ;
        RECT 96.615 168.735 97.470 168.815 ;
        RECT 99.320 168.740 99.870 168.910 ;
        RECT 100.080 168.525 100.250 169.095 ;
        RECT 100.580 169.080 100.750 170.095 ;
        RECT 100.920 169.435 101.150 169.925 ;
        RECT 101.460 169.515 101.790 169.845 ;
        RECT 100.920 168.910 101.090 169.435 ;
        RECT 102.040 169.250 102.210 169.685 ;
        RECT 102.380 169.435 102.550 170.635 ;
        RECT 102.820 169.435 102.990 169.925 ;
        RECT 101.300 169.080 102.630 169.250 ;
        RECT 100.920 168.740 101.350 168.910 ;
        RECT 101.520 168.740 102.130 168.910 ;
        RECT 94.025 167.540 94.195 168.525 ;
        RECT 93.305 167.215 93.475 167.340 ;
        RECT 93.225 167.045 93.555 167.215 ;
        RECT 93.965 167.045 94.295 167.340 ;
        RECT 94.465 166.875 94.635 168.525 ;
        RECT 94.805 167.585 95.075 168.525 ;
        RECT 95.345 166.875 95.515 168.525 ;
        RECT 96.335 166.875 96.505 168.525 ;
        RECT 96.775 167.585 96.945 168.525 ;
        RECT 97.215 166.875 97.385 168.525 ;
        RECT 97.930 166.875 98.320 168.465 ;
        RECT 98.860 166.875 99.030 168.525 ;
        RECT 99.300 167.585 99.470 168.525 ;
        RECT 99.740 166.875 99.910 168.525 ;
        RECT 100.080 167.585 100.470 168.525 ;
        RECT 100.240 167.200 100.570 167.370 ;
        RECT 100.740 166.875 100.910 168.525 ;
        RECT 101.180 167.585 101.350 168.740 ;
        RECT 101.120 167.045 101.450 167.340 ;
        RECT 101.620 166.875 101.790 168.525 ;
        RECT 101.960 167.540 102.130 168.740 ;
        RECT 102.460 167.585 102.630 169.080 ;
        RECT 102.830 168.935 103.000 169.265 ;
        RECT 103.170 168.270 103.340 170.360 ;
        RECT 103.930 169.270 104.320 170.635 ;
        RECT 104.865 169.435 105.035 170.635 ;
        RECT 102.800 167.370 102.970 168.230 ;
        RECT 102.250 167.200 102.970 167.370 ;
        RECT 103.930 166.875 104.320 168.465 ;
        RECT 104.825 166.875 104.995 168.525 ;
        RECT 105.205 167.585 105.475 169.925 ;
        RECT 105.745 169.435 105.915 170.635 ;
        RECT 106.305 170.095 106.635 170.330 ;
        RECT 106.925 170.295 107.255 170.465 ;
        RECT 105.645 168.740 106.125 169.265 ;
        RECT 105.705 166.875 105.875 168.525 ;
        RECT 106.145 167.540 106.315 168.525 ;
        RECT 106.485 167.585 106.755 169.925 ;
        RECT 106.925 169.790 107.095 170.295 ;
        RECT 107.425 169.435 107.595 170.635 ;
        RECT 107.805 169.435 108.035 169.925 ;
        RECT 108.305 169.435 108.475 170.635 ;
        RECT 109.335 169.435 109.505 170.635 ;
        RECT 109.775 169.435 109.945 169.925 ;
        RECT 110.215 169.435 110.385 170.635 ;
        RECT 106.925 168.695 107.635 169.065 ;
        RECT 107.805 168.525 107.980 169.435 ;
        RECT 110.930 169.270 111.320 170.635 ;
        RECT 111.860 169.435 112.030 170.635 ;
        RECT 112.300 169.435 112.470 169.925 ;
        RECT 112.740 169.435 112.910 170.635 ;
        RECT 113.080 170.160 113.410 170.465 ;
        RECT 113.580 170.095 114.060 170.265 ;
        RECT 114.880 170.160 115.210 170.465 ;
        RECT 113.080 169.265 113.250 169.685 ;
        RECT 108.150 168.865 108.330 169.265 ;
        RECT 109.615 169.145 110.470 169.225 ;
        RECT 108.150 168.695 108.690 168.865 ;
        RECT 109.615 168.815 110.500 169.145 ;
        RECT 112.860 169.095 113.250 169.265 ;
        RECT 109.615 168.735 110.470 168.815 ;
        RECT 112.320 168.740 112.870 168.910 ;
        RECT 113.080 168.525 113.250 169.095 ;
        RECT 113.580 169.080 113.750 170.095 ;
        RECT 113.920 169.435 114.150 169.925 ;
        RECT 114.460 169.515 114.790 169.845 ;
        RECT 113.920 168.910 114.090 169.435 ;
        RECT 115.040 169.250 115.210 169.685 ;
        RECT 115.380 169.435 115.550 170.635 ;
        RECT 115.820 169.435 115.990 169.925 ;
        RECT 114.300 169.080 115.630 169.250 ;
        RECT 113.920 168.740 114.350 168.910 ;
        RECT 114.520 168.740 115.130 168.910 ;
        RECT 107.025 167.540 107.195 168.525 ;
        RECT 106.305 167.215 106.475 167.340 ;
        RECT 106.225 167.045 106.555 167.215 ;
        RECT 106.965 167.045 107.295 167.340 ;
        RECT 107.465 166.875 107.635 168.525 ;
        RECT 107.805 167.585 108.075 168.525 ;
        RECT 108.345 166.875 108.515 168.525 ;
        RECT 109.335 166.875 109.505 168.525 ;
        RECT 109.775 167.585 109.945 168.525 ;
        RECT 110.215 166.875 110.385 168.525 ;
        RECT 110.930 166.875 111.320 168.465 ;
        RECT 111.860 166.875 112.030 168.525 ;
        RECT 112.300 167.585 112.470 168.525 ;
        RECT 112.740 166.875 112.910 168.525 ;
        RECT 113.080 167.585 113.470 168.525 ;
        RECT 113.240 167.200 113.570 167.370 ;
        RECT 113.740 166.875 113.910 168.525 ;
        RECT 114.180 167.585 114.350 168.740 ;
        RECT 114.120 167.045 114.450 167.340 ;
        RECT 114.620 166.875 114.790 168.525 ;
        RECT 114.960 167.540 115.130 168.740 ;
        RECT 115.460 167.585 115.630 169.080 ;
        RECT 115.830 168.935 116.000 169.265 ;
        RECT 116.170 168.270 116.340 170.360 ;
        RECT 120.680 169.270 121.070 170.635 ;
        RECT 121.615 169.435 121.785 170.635 ;
        RECT 122.055 169.435 122.225 169.925 ;
        RECT 122.495 169.435 122.665 170.635 ;
        RECT 123.365 169.435 123.535 170.635 ;
        RECT 123.805 169.435 123.975 169.925 ;
        RECT 124.245 169.435 124.415 170.635 ;
        RECT 125.115 169.435 125.285 170.635 ;
        RECT 125.555 169.435 125.725 169.925 ;
        RECT 125.995 169.435 126.165 170.635 ;
        RECT 126.865 169.435 127.035 170.635 ;
        RECT 127.305 169.435 127.475 169.925 ;
        RECT 127.745 169.435 127.915 170.635 ;
        RECT 128.430 169.270 128.820 170.635 ;
        RECT 129.365 169.435 129.535 170.635 ;
        RECT 129.805 169.435 129.975 169.925 ;
        RECT 130.245 169.435 130.415 170.635 ;
        RECT 131.170 169.435 131.840 169.925 ;
        RECT 132.010 169.435 132.180 170.635 ;
        RECT 132.450 169.435 132.620 169.925 ;
        RECT 132.890 169.435 133.060 170.635 ;
        RECT 133.430 169.270 133.820 170.635 ;
        RECT 134.310 169.435 134.480 170.635 ;
        RECT 134.750 169.435 134.920 170.090 ;
        RECT 135.190 169.435 135.360 170.635 ;
        RECT 135.630 169.435 135.800 169.925 ;
        RECT 136.070 169.435 136.240 170.635 ;
        RECT 136.865 169.435 137.035 170.635 ;
        RECT 137.305 169.435 137.475 169.925 ;
        RECT 137.745 169.435 137.915 170.635 ;
        RECT 138.430 169.270 138.820 170.635 ;
        RECT 121.530 169.145 122.385 169.225 ;
        RECT 123.280 169.145 124.135 169.225 ;
        RECT 125.030 169.145 125.885 169.225 ;
        RECT 126.780 169.145 127.635 169.225 ;
        RECT 129.280 169.145 130.135 169.225 ;
        RECT 121.500 168.815 122.385 169.145 ;
        RECT 123.250 168.815 124.135 169.145 ;
        RECT 125.000 168.815 125.885 169.145 ;
        RECT 126.750 168.815 127.635 169.145 ;
        RECT 129.250 168.815 130.135 169.145 ;
        RECT 131.060 169.095 132.060 169.265 ;
        RECT 134.310 169.095 135.240 169.265 ;
        RECT 136.780 169.145 137.635 169.225 ;
        RECT 131.730 169.075 132.060 169.095 ;
        RECT 121.530 168.735 122.385 168.815 ;
        RECT 123.280 168.735 124.135 168.815 ;
        RECT 125.030 168.735 125.885 168.815 ;
        RECT 126.780 168.735 127.635 168.815 ;
        RECT 129.280 168.735 130.135 168.815 ;
        RECT 131.000 168.695 131.540 168.910 ;
        RECT 132.240 168.905 132.570 168.950 ;
        RECT 131.880 168.735 132.570 168.905 ;
        RECT 134.250 168.695 134.580 168.910 ;
        RECT 135.380 168.740 135.720 168.995 ;
        RECT 136.750 168.815 137.635 169.145 ;
        RECT 136.780 168.735 137.635 168.815 ;
        RECT 115.800 167.370 115.970 168.230 ;
        RECT 115.250 167.200 115.970 167.370 ;
        RECT 120.680 166.875 121.070 168.465 ;
        RECT 121.615 166.875 121.785 168.525 ;
        RECT 122.055 167.585 122.225 168.525 ;
        RECT 122.495 166.875 122.665 168.525 ;
        RECT 123.365 166.875 123.535 168.525 ;
        RECT 123.805 167.585 123.975 168.525 ;
        RECT 124.245 166.875 124.415 168.525 ;
        RECT 125.115 166.875 125.285 168.525 ;
        RECT 125.555 167.585 125.725 168.525 ;
        RECT 125.995 166.875 126.165 168.525 ;
        RECT 126.865 166.875 127.035 168.525 ;
        RECT 127.305 167.585 127.475 168.525 ;
        RECT 127.745 166.875 127.915 168.525 ;
        RECT 128.430 166.875 128.820 168.465 ;
        RECT 129.365 166.875 129.535 168.525 ;
        RECT 129.805 167.585 129.975 168.525 ;
        RECT 130.245 166.875 130.415 168.525 ;
        RECT 131.130 166.875 131.300 168.525 ;
        RECT 131.570 167.585 131.840 168.525 ;
        RECT 132.010 166.875 132.180 168.525 ;
        RECT 132.450 167.585 132.620 168.525 ;
        RECT 132.890 166.875 133.060 168.525 ;
        RECT 133.430 166.875 133.820 168.465 ;
        RECT 134.350 167.585 134.520 168.525 ;
        RECT 135.190 166.875 135.360 168.525 ;
        RECT 135.630 167.585 135.800 168.525 ;
        RECT 136.070 166.875 136.240 168.525 ;
        RECT 136.865 166.875 137.035 168.525 ;
        RECT 137.305 167.585 137.475 168.525 ;
        RECT 137.745 166.875 137.915 168.525 ;
        RECT 138.430 166.875 138.820 168.465 ;
        RECT 81.000 166.625 88.500 166.875 ;
        RECT 90.750 166.625 139.000 166.875 ;
        RECT 87.500 163.635 144.750 163.885 ;
        RECT 87.680 162.270 88.070 163.635 ;
        RECT 88.585 162.435 88.755 163.635 ;
        RECT 89.025 162.435 89.195 162.925 ;
        RECT 89.465 162.435 89.635 163.635 ;
        RECT 90.335 162.435 90.505 163.635 ;
        RECT 90.775 162.435 90.945 162.925 ;
        RECT 91.215 162.435 91.385 163.635 ;
        RECT 92.120 162.435 92.290 163.635 ;
        RECT 92.460 162.435 92.730 162.925 ;
        RECT 93.000 162.435 93.170 163.635 ;
        RECT 93.600 163.115 95.110 163.465 ;
        RECT 93.840 162.605 94.010 162.925 ;
        RECT 93.560 162.435 94.010 162.605 ;
        RECT 94.340 162.435 94.610 162.925 ;
        RECT 95.280 162.435 95.450 163.635 ;
        RECT 95.620 162.435 95.890 162.925 ;
        RECT 88.865 162.145 89.720 162.225 ;
        RECT 90.615 162.145 91.470 162.225 ;
        RECT 88.865 161.815 89.750 162.145 ;
        RECT 90.615 161.815 91.500 162.145 ;
        RECT 88.865 161.735 89.720 161.815 ;
        RECT 90.615 161.735 91.470 161.815 ;
        RECT 92.460 161.525 92.630 162.435 ;
        RECT 93.560 162.145 93.730 162.435 ;
        RECT 92.800 161.815 93.730 162.145 ;
        RECT 93.900 162.140 94.070 162.145 ;
        RECT 94.340 162.140 94.510 162.435 ;
        RECT 93.900 161.815 94.510 162.140 ;
        RECT 95.620 162.065 95.790 162.435 ;
        RECT 94.680 161.895 95.790 162.065 ;
        RECT 87.680 159.875 88.070 161.465 ;
        RECT 88.585 159.875 88.755 161.525 ;
        RECT 89.025 160.585 89.195 161.525 ;
        RECT 89.465 159.875 89.635 161.525 ;
        RECT 90.335 159.875 90.505 161.525 ;
        RECT 90.775 160.585 90.945 161.525 ;
        RECT 91.215 159.875 91.385 161.525 ;
        RECT 92.120 159.875 92.290 161.525 ;
        RECT 92.460 160.585 92.730 161.525 ;
        RECT 93.000 159.875 93.170 161.525 ;
        RECT 93.560 160.585 93.730 161.815 ;
        RECT 94.340 161.525 94.510 161.815 ;
        RECT 95.620 161.525 95.790 161.895 ;
        RECT 95.960 161.815 96.130 162.145 ;
        RECT 94.000 159.875 94.170 161.525 ;
        RECT 94.340 160.585 94.610 161.525 ;
        RECT 94.340 160.200 94.670 160.370 ;
        RECT 95.000 159.875 95.170 161.525 ;
        RECT 95.620 160.585 96.010 161.525 ;
        RECT 96.300 161.500 96.470 163.315 ;
        RECT 96.930 162.270 97.320 163.635 ;
        RECT 97.870 162.435 98.040 163.635 ;
        RECT 98.210 162.435 98.480 162.925 ;
        RECT 98.750 162.435 98.920 163.635 ;
        RECT 99.350 163.115 100.860 163.465 ;
        RECT 99.590 162.605 99.760 162.925 ;
        RECT 99.310 162.435 99.760 162.605 ;
        RECT 100.090 162.435 100.360 162.925 ;
        RECT 101.030 162.435 101.200 163.635 ;
        RECT 101.370 162.435 101.640 162.925 ;
        RECT 98.210 161.525 98.380 162.435 ;
        RECT 99.310 162.145 99.480 162.435 ;
        RECT 98.550 161.815 99.480 162.145 ;
        RECT 99.650 162.140 99.820 162.145 ;
        RECT 100.090 162.140 100.260 162.435 ;
        RECT 99.650 161.815 100.260 162.140 ;
        RECT 101.370 162.065 101.540 162.435 ;
        RECT 100.430 161.895 101.540 162.065 ;
        RECT 96.180 161.000 96.470 161.500 ;
        RECT 95.600 160.200 95.930 160.370 ;
        RECT 96.300 160.170 96.470 161.000 ;
        RECT 96.930 159.875 97.320 161.465 ;
        RECT 97.870 159.875 98.040 161.525 ;
        RECT 98.210 160.585 98.480 161.525 ;
        RECT 98.750 159.875 98.920 161.525 ;
        RECT 99.310 160.585 99.480 161.815 ;
        RECT 100.090 161.525 100.260 161.815 ;
        RECT 101.370 161.525 101.540 161.895 ;
        RECT 101.710 161.815 101.880 162.145 ;
        RECT 99.750 159.875 99.920 161.525 ;
        RECT 100.090 160.585 100.360 161.525 ;
        RECT 100.090 160.200 100.420 160.370 ;
        RECT 100.750 159.875 100.920 161.525 ;
        RECT 101.370 160.585 101.760 161.525 ;
        RECT 102.050 161.500 102.220 163.315 ;
        RECT 102.870 162.435 103.040 163.635 ;
        RECT 103.210 162.435 103.480 162.925 ;
        RECT 103.750 162.435 103.920 163.635 ;
        RECT 104.350 163.115 105.860 163.465 ;
        RECT 104.590 162.605 104.760 162.925 ;
        RECT 104.310 162.435 104.760 162.605 ;
        RECT 105.090 162.435 105.360 162.925 ;
        RECT 106.030 162.435 106.200 163.635 ;
        RECT 106.370 162.435 106.640 162.925 ;
        RECT 103.210 161.525 103.380 162.435 ;
        RECT 104.310 162.145 104.480 162.435 ;
        RECT 103.550 161.815 104.480 162.145 ;
        RECT 104.650 162.140 104.820 162.145 ;
        RECT 105.090 162.140 105.260 162.435 ;
        RECT 104.650 161.815 105.260 162.140 ;
        RECT 106.370 162.065 106.540 162.435 ;
        RECT 105.430 161.895 106.540 162.065 ;
        RECT 101.930 161.000 102.220 161.500 ;
        RECT 101.350 160.200 101.680 160.370 ;
        RECT 102.050 160.170 102.220 161.000 ;
        RECT 102.870 159.875 103.040 161.525 ;
        RECT 103.210 160.585 103.480 161.525 ;
        RECT 103.750 159.875 103.920 161.525 ;
        RECT 104.310 160.585 104.480 161.815 ;
        RECT 105.090 161.525 105.260 161.815 ;
        RECT 106.370 161.525 106.540 161.895 ;
        RECT 106.710 161.815 106.880 162.145 ;
        RECT 104.750 159.875 104.920 161.525 ;
        RECT 105.090 160.585 105.360 161.525 ;
        RECT 105.090 160.200 105.420 160.370 ;
        RECT 105.750 159.875 105.920 161.525 ;
        RECT 106.370 160.585 106.760 161.525 ;
        RECT 107.050 161.500 107.220 163.315 ;
        RECT 107.680 162.270 108.070 163.635 ;
        RECT 108.585 162.435 108.755 163.635 ;
        RECT 109.025 162.435 109.195 162.925 ;
        RECT 109.465 162.435 109.635 163.635 ;
        RECT 110.370 162.435 110.540 163.635 ;
        RECT 110.710 162.435 110.980 162.925 ;
        RECT 111.250 162.435 111.420 163.635 ;
        RECT 111.850 163.115 113.360 163.465 ;
        RECT 112.090 162.605 112.260 162.925 ;
        RECT 111.810 162.435 112.260 162.605 ;
        RECT 112.590 162.435 112.860 162.925 ;
        RECT 113.530 162.435 113.700 163.635 ;
        RECT 113.870 162.435 114.140 162.925 ;
        RECT 108.865 162.145 109.720 162.225 ;
        RECT 108.865 161.815 109.750 162.145 ;
        RECT 108.865 161.735 109.720 161.815 ;
        RECT 110.710 161.525 110.880 162.435 ;
        RECT 111.810 162.145 111.980 162.435 ;
        RECT 111.050 161.815 111.980 162.145 ;
        RECT 112.150 162.140 112.320 162.145 ;
        RECT 112.590 162.140 112.760 162.435 ;
        RECT 112.150 161.815 112.760 162.140 ;
        RECT 113.870 162.065 114.040 162.435 ;
        RECT 112.930 161.895 114.040 162.065 ;
        RECT 106.930 161.000 107.220 161.500 ;
        RECT 106.350 160.200 106.680 160.370 ;
        RECT 107.050 160.170 107.220 161.000 ;
        RECT 107.680 159.875 108.070 161.465 ;
        RECT 108.585 159.875 108.755 161.525 ;
        RECT 109.025 160.585 109.195 161.525 ;
        RECT 109.465 159.875 109.635 161.525 ;
        RECT 110.370 159.875 110.540 161.525 ;
        RECT 110.710 160.585 110.980 161.525 ;
        RECT 111.250 159.875 111.420 161.525 ;
        RECT 111.810 160.585 111.980 161.815 ;
        RECT 112.590 161.525 112.760 161.815 ;
        RECT 113.870 161.525 114.040 161.895 ;
        RECT 114.210 161.815 114.380 162.145 ;
        RECT 112.250 159.875 112.420 161.525 ;
        RECT 112.590 160.585 112.860 161.525 ;
        RECT 112.590 160.200 112.920 160.370 ;
        RECT 113.250 159.875 113.420 161.525 ;
        RECT 113.870 160.585 114.260 161.525 ;
        RECT 114.550 161.500 114.720 163.315 ;
        RECT 115.190 162.435 115.360 163.635 ;
        RECT 115.630 162.435 115.800 162.925 ;
        RECT 116.070 162.435 116.240 163.635 ;
        RECT 116.410 162.435 117.080 162.925 ;
        RECT 117.680 162.270 118.070 163.635 ;
        RECT 118.620 162.435 118.790 163.635 ;
        RECT 118.960 162.435 119.230 162.925 ;
        RECT 119.500 162.435 119.670 163.635 ;
        RECT 120.100 163.115 121.610 163.465 ;
        RECT 120.340 162.605 120.510 162.925 ;
        RECT 120.060 162.435 120.510 162.605 ;
        RECT 120.840 162.435 121.110 162.925 ;
        RECT 121.780 162.435 121.950 163.635 ;
        RECT 122.120 162.435 122.390 162.925 ;
        RECT 116.190 162.095 117.190 162.265 ;
        RECT 116.190 162.075 116.520 162.095 ;
        RECT 115.680 161.905 116.010 161.950 ;
        RECT 115.680 161.735 116.370 161.905 ;
        RECT 116.710 161.695 117.250 161.910 ;
        RECT 118.960 161.525 119.130 162.435 ;
        RECT 120.060 162.145 120.230 162.435 ;
        RECT 119.300 161.815 120.230 162.145 ;
        RECT 120.400 162.140 120.570 162.145 ;
        RECT 120.840 162.140 121.010 162.435 ;
        RECT 120.400 161.815 121.010 162.140 ;
        RECT 122.120 162.065 122.290 162.435 ;
        RECT 121.180 161.895 122.290 162.065 ;
        RECT 114.430 161.000 114.720 161.500 ;
        RECT 113.850 160.200 114.180 160.370 ;
        RECT 114.550 160.170 114.720 161.000 ;
        RECT 115.190 159.875 115.360 161.525 ;
        RECT 115.630 160.585 115.800 161.525 ;
        RECT 116.070 159.875 116.240 161.525 ;
        RECT 116.410 160.585 116.680 161.525 ;
        RECT 116.950 159.875 117.120 161.525 ;
        RECT 117.680 159.875 118.070 161.465 ;
        RECT 118.620 159.875 118.790 161.525 ;
        RECT 118.960 160.585 119.230 161.525 ;
        RECT 119.500 159.875 119.670 161.525 ;
        RECT 120.060 160.585 120.230 161.815 ;
        RECT 120.840 161.525 121.010 161.815 ;
        RECT 122.120 161.525 122.290 161.895 ;
        RECT 122.460 161.815 122.630 162.145 ;
        RECT 120.500 159.875 120.670 161.525 ;
        RECT 120.840 160.585 121.110 161.525 ;
        RECT 120.840 160.200 121.170 160.370 ;
        RECT 121.500 159.875 121.670 161.525 ;
        RECT 122.120 160.585 122.510 161.525 ;
        RECT 122.800 161.500 122.970 163.315 ;
        RECT 123.620 162.435 123.790 163.635 ;
        RECT 123.960 162.435 124.230 162.925 ;
        RECT 124.500 162.435 124.670 163.635 ;
        RECT 125.100 163.115 126.610 163.465 ;
        RECT 125.340 162.605 125.510 162.925 ;
        RECT 125.060 162.435 125.510 162.605 ;
        RECT 125.840 162.435 126.110 162.925 ;
        RECT 126.780 162.435 126.950 163.635 ;
        RECT 127.120 162.435 127.390 162.925 ;
        RECT 123.960 161.525 124.130 162.435 ;
        RECT 125.060 162.145 125.230 162.435 ;
        RECT 124.300 161.815 125.230 162.145 ;
        RECT 125.400 162.140 125.570 162.145 ;
        RECT 125.840 162.140 126.010 162.435 ;
        RECT 125.400 161.815 126.010 162.140 ;
        RECT 127.120 162.065 127.290 162.435 ;
        RECT 126.180 161.895 127.290 162.065 ;
        RECT 122.680 161.000 122.970 161.500 ;
        RECT 122.100 160.200 122.430 160.370 ;
        RECT 122.800 160.170 122.970 161.000 ;
        RECT 123.620 159.875 123.790 161.525 ;
        RECT 123.960 160.585 124.230 161.525 ;
        RECT 124.500 159.875 124.670 161.525 ;
        RECT 125.060 160.585 125.230 161.815 ;
        RECT 125.840 161.525 126.010 161.815 ;
        RECT 127.120 161.525 127.290 161.895 ;
        RECT 127.460 161.815 127.630 162.145 ;
        RECT 125.500 159.875 125.670 161.525 ;
        RECT 125.840 160.585 126.110 161.525 ;
        RECT 125.840 160.200 126.170 160.370 ;
        RECT 126.500 159.875 126.670 161.525 ;
        RECT 127.120 160.585 127.510 161.525 ;
        RECT 127.800 161.500 127.970 163.315 ;
        RECT 128.640 162.435 128.810 163.635 ;
        RECT 128.580 162.095 128.910 162.265 ;
        RECT 129.080 161.865 129.250 162.925 ;
        RECT 129.520 162.435 129.690 163.635 ;
        RECT 130.180 162.270 130.570 163.635 ;
        RECT 131.140 162.435 131.310 163.635 ;
        RECT 131.080 162.095 131.410 162.265 ;
        RECT 128.560 161.695 129.250 161.865 ;
        RECT 129.420 161.695 129.750 161.910 ;
        RECT 131.580 161.865 131.750 162.925 ;
        RECT 132.020 162.435 132.190 163.635 ;
        RECT 132.835 162.435 133.005 163.635 ;
        RECT 133.275 162.435 133.445 162.925 ;
        RECT 133.715 162.435 133.885 163.635 ;
        RECT 134.620 162.435 134.790 163.635 ;
        RECT 134.960 162.435 135.230 162.925 ;
        RECT 135.500 162.435 135.670 163.635 ;
        RECT 136.100 163.115 137.610 163.465 ;
        RECT 136.340 162.605 136.510 162.925 ;
        RECT 136.060 162.435 136.510 162.605 ;
        RECT 136.840 162.435 137.110 162.925 ;
        RECT 137.780 162.435 137.950 163.635 ;
        RECT 138.120 162.435 138.390 162.925 ;
        RECT 133.115 162.145 133.970 162.225 ;
        RECT 131.060 161.695 131.750 161.865 ;
        RECT 131.920 161.695 132.250 161.910 ;
        RECT 133.115 161.815 134.000 162.145 ;
        RECT 133.115 161.735 133.970 161.815 ;
        RECT 134.960 161.525 135.130 162.435 ;
        RECT 136.060 162.145 136.230 162.435 ;
        RECT 135.300 161.815 136.230 162.145 ;
        RECT 136.400 162.140 136.570 162.145 ;
        RECT 136.840 162.140 137.010 162.435 ;
        RECT 136.400 161.815 137.010 162.140 ;
        RECT 138.120 162.065 138.290 162.435 ;
        RECT 137.180 161.895 138.290 162.065 ;
        RECT 127.680 161.000 127.970 161.500 ;
        RECT 127.100 160.200 127.430 160.370 ;
        RECT 127.800 160.170 127.970 161.000 ;
        RECT 128.640 160.585 128.810 161.525 ;
        RECT 129.480 159.875 129.650 161.525 ;
        RECT 130.180 159.875 130.570 161.465 ;
        RECT 131.140 160.585 131.310 161.525 ;
        RECT 131.980 159.875 132.150 161.525 ;
        RECT 132.835 159.875 133.005 161.525 ;
        RECT 133.275 160.585 133.445 161.525 ;
        RECT 133.715 159.875 133.885 161.525 ;
        RECT 134.620 159.875 134.790 161.525 ;
        RECT 134.960 160.585 135.230 161.525 ;
        RECT 135.500 159.875 135.670 161.525 ;
        RECT 136.060 160.585 136.230 161.815 ;
        RECT 136.840 161.525 137.010 161.815 ;
        RECT 138.120 161.525 138.290 161.895 ;
        RECT 138.460 161.815 138.630 162.145 ;
        RECT 136.500 159.875 136.670 161.525 ;
        RECT 136.840 160.585 137.110 161.525 ;
        RECT 136.840 160.200 137.170 160.370 ;
        RECT 137.500 159.875 137.670 161.525 ;
        RECT 138.120 160.585 138.510 161.525 ;
        RECT 138.800 161.500 138.970 163.315 ;
        RECT 139.620 162.435 139.790 163.635 ;
        RECT 139.960 162.435 140.230 162.925 ;
        RECT 140.500 162.435 140.670 163.635 ;
        RECT 141.100 163.115 142.610 163.465 ;
        RECT 141.340 162.605 141.510 162.925 ;
        RECT 141.060 162.435 141.510 162.605 ;
        RECT 141.840 162.435 142.110 162.925 ;
        RECT 142.780 162.435 142.950 163.635 ;
        RECT 143.120 162.435 143.390 162.925 ;
        RECT 139.960 161.525 140.130 162.435 ;
        RECT 141.060 162.145 141.230 162.435 ;
        RECT 140.300 161.815 141.230 162.145 ;
        RECT 141.400 162.140 141.570 162.145 ;
        RECT 141.840 162.140 142.010 162.435 ;
        RECT 141.400 161.815 142.010 162.140 ;
        RECT 143.120 162.065 143.290 162.435 ;
        RECT 142.180 161.895 143.290 162.065 ;
        RECT 138.680 161.000 138.970 161.500 ;
        RECT 138.100 160.200 138.430 160.370 ;
        RECT 138.800 160.170 138.970 161.000 ;
        RECT 139.620 159.875 139.790 161.525 ;
        RECT 139.960 160.585 140.230 161.525 ;
        RECT 140.500 159.875 140.670 161.525 ;
        RECT 141.060 160.585 141.230 161.815 ;
        RECT 141.840 161.525 142.010 161.815 ;
        RECT 143.120 161.525 143.290 161.895 ;
        RECT 143.460 161.815 143.630 162.145 ;
        RECT 141.500 159.875 141.670 161.525 ;
        RECT 141.840 160.585 142.110 161.525 ;
        RECT 141.840 160.200 142.170 160.370 ;
        RECT 142.500 159.875 142.670 161.525 ;
        RECT 143.120 160.585 143.510 161.525 ;
        RECT 143.800 161.500 143.970 163.315 ;
        RECT 144.180 162.270 144.570 163.635 ;
        RECT 143.680 161.000 143.970 161.500 ;
        RECT 143.100 160.200 143.430 160.370 ;
        RECT 143.800 160.170 143.970 161.000 ;
        RECT 144.180 159.875 144.570 161.465 ;
        RECT 87.500 159.625 144.750 159.875 ;
        RECT 145.250 156.750 145.750 180.750 ;
        RECT 77.500 156.250 145.750 156.750 ;
        RECT 22.875 150.125 41.125 150.375 ;
        RECT 41.875 155.125 52.625 155.375 ;
        RECT 11.125 149.125 22.375 149.375 ;
        RECT 11.125 144.875 11.375 149.125 ;
        RECT 13.910 148.250 14.080 148.750 ;
        RECT 11.715 145.230 11.885 147.270 ;
        RECT 12.155 145.230 12.325 147.270 ;
        RECT 12.595 145.230 12.765 147.270 ;
        RECT 13.035 145.230 13.205 147.270 ;
        RECT 13.475 145.230 13.645 147.270 ;
        RECT 13.915 145.230 14.085 147.270 ;
        RECT 14.355 145.230 14.525 147.270 ;
        RECT 14.795 145.230 14.965 147.270 ;
        RECT 15.235 145.230 15.405 147.270 ;
        RECT 15.675 145.230 15.845 147.270 ;
        RECT 16.115 145.230 16.285 147.270 ;
        RECT 16.625 144.875 16.875 149.125 ;
        RECT 19.410 148.250 19.580 148.750 ;
        RECT 17.215 145.230 17.385 147.270 ;
        RECT 17.655 145.230 17.825 147.270 ;
        RECT 18.095 145.230 18.265 147.270 ;
        RECT 18.535 145.230 18.705 147.270 ;
        RECT 18.975 145.230 19.145 147.270 ;
        RECT 19.415 145.230 19.585 147.270 ;
        RECT 19.855 145.230 20.025 147.270 ;
        RECT 20.295 145.230 20.465 147.270 ;
        RECT 20.735 145.230 20.905 147.270 ;
        RECT 21.175 145.230 21.345 147.270 ;
        RECT 21.615 145.230 21.785 147.270 ;
        RECT 22.125 144.875 22.375 149.125 ;
        RECT 11.125 144.625 22.375 144.875 ;
        RECT 22.875 149.125 41.125 149.375 ;
        RECT 22.875 142.875 23.125 149.125 ;
        RECT 25.915 148.250 26.085 148.750 ;
        RECT 23.615 143.230 23.785 147.270 ;
        RECT 24.075 143.230 24.245 147.270 ;
        RECT 24.535 143.230 24.705 147.270 ;
        RECT 24.995 143.230 25.165 147.270 ;
        RECT 25.455 143.230 25.625 147.270 ;
        RECT 25.915 143.230 26.085 147.270 ;
        RECT 26.375 143.230 26.545 147.270 ;
        RECT 26.835 143.230 27.005 147.270 ;
        RECT 27.295 143.230 27.465 147.270 ;
        RECT 27.755 143.230 27.925 147.270 ;
        RECT 28.215 143.230 28.385 147.270 ;
        RECT 28.875 142.875 29.125 149.125 ;
        RECT 31.915 148.250 32.085 148.750 ;
        RECT 29.615 143.230 29.785 147.270 ;
        RECT 30.075 143.230 30.245 147.270 ;
        RECT 30.535 143.230 30.705 147.270 ;
        RECT 30.995 143.230 31.165 147.270 ;
        RECT 31.455 143.230 31.625 147.270 ;
        RECT 31.915 143.230 32.085 147.270 ;
        RECT 32.375 143.230 32.545 147.270 ;
        RECT 32.835 143.230 33.005 147.270 ;
        RECT 33.295 143.230 33.465 147.270 ;
        RECT 33.755 143.230 33.925 147.270 ;
        RECT 34.215 143.230 34.385 147.270 ;
        RECT 34.875 142.875 35.125 149.125 ;
        RECT 37.915 148.250 38.085 148.750 ;
        RECT 35.615 143.230 35.785 147.270 ;
        RECT 36.075 143.230 36.245 147.270 ;
        RECT 36.535 143.230 36.705 147.270 ;
        RECT 36.995 143.230 37.165 147.270 ;
        RECT 37.455 143.230 37.625 147.270 ;
        RECT 37.915 143.230 38.085 147.270 ;
        RECT 38.375 143.230 38.545 147.270 ;
        RECT 38.835 143.230 39.005 147.270 ;
        RECT 39.295 143.230 39.465 147.270 ;
        RECT 39.755 143.230 39.925 147.270 ;
        RECT 40.215 143.230 40.385 147.270 ;
        RECT 40.875 142.875 41.125 149.125 ;
        RECT 41.875 144.375 42.125 155.125 ;
        RECT 43.415 154.250 44.085 154.750 ;
        RECT 42.530 145.480 43.190 154.020 ;
        RECT 44.310 145.480 44.970 154.020 ;
        RECT 43.415 144.750 44.085 145.250 ;
        RECT 45.375 144.375 45.625 155.125 ;
        RECT 46.915 154.250 47.585 154.750 ;
        RECT 46.030 145.480 46.690 154.020 ;
        RECT 47.810 145.480 48.470 154.020 ;
        RECT 46.915 144.750 47.585 145.250 ;
        RECT 48.875 144.375 49.125 155.125 ;
        RECT 50.415 154.250 51.085 154.750 ;
        RECT 49.530 145.480 50.190 154.020 ;
        RECT 51.310 145.480 51.970 154.020 ;
        RECT 50.415 144.750 51.085 145.250 ;
        RECT 52.375 144.375 52.625 155.125 ;
        RECT 114.600 149.035 138.980 149.205 ;
        RECT 114.685 148.285 115.895 149.035 ;
        RECT 114.685 147.745 115.205 148.285 ;
        RECT 116.525 148.265 120.035 149.035 ;
        RECT 120.210 148.490 125.555 149.035 ;
        RECT 115.375 147.575 115.895 148.115 ;
        RECT 114.685 146.485 115.895 147.575 ;
        RECT 116.525 147.575 118.215 148.095 ;
        RECT 118.385 147.745 120.035 148.265 ;
        RECT 116.525 146.485 120.035 147.575 ;
        RECT 121.800 146.920 122.150 148.170 ;
        RECT 123.630 147.660 123.970 148.490 ;
        RECT 125.725 148.310 126.015 149.035 ;
        RECT 126.650 148.490 131.995 149.035 ;
        RECT 132.170 148.490 137.515 149.035 ;
        RECT 120.210 146.485 125.555 146.920 ;
        RECT 125.725 146.485 126.015 147.650 ;
        RECT 128.240 146.920 128.590 148.170 ;
        RECT 130.070 147.660 130.410 148.490 ;
        RECT 133.760 146.920 134.110 148.170 ;
        RECT 135.590 147.660 135.930 148.490 ;
        RECT 137.685 148.285 138.895 149.035 ;
        RECT 137.685 147.575 138.205 148.115 ;
        RECT 138.375 147.745 138.895 148.285 ;
        RECT 126.650 146.485 131.995 146.920 ;
        RECT 132.170 146.485 137.515 146.920 ;
        RECT 137.685 146.485 138.895 147.575 ;
        RECT 114.600 146.315 138.980 146.485 ;
        RECT 114.685 145.225 115.895 146.315 ;
        RECT 41.875 144.125 52.625 144.375 ;
        RECT 114.685 144.515 115.205 145.055 ;
        RECT 115.375 144.685 115.895 145.225 ;
        RECT 116.065 145.225 117.275 146.315 ;
        RECT 117.455 145.345 117.745 146.315 ;
        RECT 116.065 144.685 116.585 145.225 ;
        RECT 116.755 144.515 117.275 145.055 ;
        RECT 114.685 143.765 115.895 144.515 ;
        RECT 116.065 143.765 117.275 144.515 ;
        RECT 117.915 144.505 118.145 146.145 ;
        RECT 118.315 145.900 118.645 146.315 ;
        RECT 118.835 145.600 119.150 146.145 ;
        RECT 118.315 145.370 119.150 145.600 ;
        RECT 119.320 145.615 119.545 146.145 ;
        RECT 119.715 145.805 120.045 146.315 ;
        RECT 120.215 145.615 120.435 146.145 ;
        RECT 118.315 144.675 118.655 145.370 ;
        RECT 119.320 145.350 120.435 145.615 ;
        RECT 121.125 145.225 124.635 146.315 ;
        RECT 124.810 145.880 130.155 146.315 ;
        RECT 118.825 144.675 119.150 145.090 ;
        RECT 118.485 144.505 118.655 144.675 ;
        RECT 117.915 144.315 118.315 144.505 ;
        RECT 118.485 144.335 119.225 144.505 ;
        RECT 117.625 143.765 117.955 144.145 ;
        RECT 118.125 143.935 118.315 144.315 ;
        RECT 118.485 143.765 118.815 144.125 ;
        RECT 119.035 143.935 119.225 144.335 ;
        RECT 119.600 144.045 119.980 145.005 ;
        RECT 120.170 144.430 120.485 145.005 ;
        RECT 121.125 144.705 122.815 145.225 ;
        RECT 122.985 144.535 124.635 145.055 ;
        RECT 126.400 144.630 126.750 145.880 ;
        RECT 130.525 145.645 130.805 146.315 ;
        RECT 120.165 143.765 120.495 144.245 ;
        RECT 121.125 143.765 124.635 144.535 ;
        RECT 128.230 144.310 128.570 145.140 ;
        RECT 130.325 145.005 130.640 145.445 ;
        RECT 130.975 145.425 131.275 145.975 ;
        RECT 131.485 145.595 131.815 146.315 ;
        RECT 132.005 145.595 132.455 146.145 ;
        RECT 130.975 145.255 131.915 145.425 ;
        RECT 131.745 145.005 131.915 145.255 ;
        RECT 130.325 144.755 131.015 145.005 ;
        RECT 131.245 144.755 131.575 145.005 ;
        RECT 131.745 144.675 132.035 145.005 ;
        RECT 131.745 144.585 131.915 144.675 ;
        RECT 130.525 144.395 131.915 144.585 ;
        RECT 124.810 143.765 130.155 144.310 ;
        RECT 130.525 144.035 130.855 144.395 ;
        RECT 132.205 144.225 132.455 145.595 ;
        RECT 132.625 145.175 132.915 146.315 ;
        RECT 133.145 145.615 133.365 146.145 ;
        RECT 133.535 145.805 133.865 146.315 ;
        RECT 134.035 145.615 134.260 146.145 ;
        RECT 133.145 145.350 134.260 145.615 ;
        RECT 134.430 145.600 134.745 146.145 ;
        RECT 134.935 145.900 135.265 146.315 ;
        RECT 134.430 145.370 135.265 145.600 ;
        RECT 131.485 143.765 131.735 144.225 ;
        RECT 131.905 143.935 132.455 144.225 ;
        RECT 132.625 143.765 132.915 144.565 ;
        RECT 133.095 144.430 133.410 145.005 ;
        RECT 133.085 143.765 133.415 144.245 ;
        RECT 133.600 144.045 133.980 145.005 ;
        RECT 134.430 144.675 134.755 145.090 ;
        RECT 134.925 144.675 135.265 145.370 ;
        RECT 134.925 144.505 135.095 144.675 ;
        RECT 135.435 144.505 135.665 146.145 ;
        RECT 135.835 145.345 136.125 146.315 ;
        RECT 136.495 145.590 136.825 146.315 ;
        RECT 134.355 144.335 135.095 144.505 ;
        RECT 134.355 143.935 134.545 144.335 ;
        RECT 135.265 144.315 135.665 144.505 ;
        RECT 134.765 143.765 135.095 144.125 ;
        RECT 135.265 143.935 135.455 144.315 ;
        RECT 135.625 143.765 135.955 144.145 ;
        RECT 136.305 143.935 136.825 145.420 ;
        RECT 136.995 144.595 137.515 146.145 ;
        RECT 137.685 145.225 138.895 146.315 ;
        RECT 137.685 144.685 138.205 145.225 ;
        RECT 138.375 144.515 138.895 145.055 ;
        RECT 136.995 143.765 137.335 144.425 ;
        RECT 137.685 143.765 138.895 144.515 ;
        RECT 114.600 143.595 138.980 143.765 ;
        RECT 22.875 142.625 41.125 142.875 ;
        RECT 114.685 142.845 115.895 143.595 ;
        RECT 114.685 142.305 115.205 142.845 ;
        RECT 116.525 142.825 118.195 143.595 ;
        RECT 118.545 143.215 118.875 143.595 ;
        RECT 119.045 143.045 119.235 143.425 ;
        RECT 119.405 143.235 119.735 143.595 ;
        RECT 115.375 142.135 115.895 142.675 ;
        RECT 21.625 141.375 24.875 141.625 ;
        RECT 21.625 137.875 21.875 141.375 ;
        RECT 23.165 140.500 23.335 141.000 ;
        RECT 22.280 139.230 22.760 140.270 ;
        RECT 23.030 139.230 23.470 140.270 ;
        RECT 23.740 139.230 24.220 140.270 ;
        RECT 23.165 138.500 23.335 139.000 ;
        RECT 24.625 137.875 24.875 141.375 ;
        RECT 21.625 137.625 24.875 137.875 ;
        RECT 21.625 134.125 21.875 137.625 ;
        RECT 23.165 136.750 23.335 137.250 ;
        RECT 22.280 135.480 22.760 136.520 ;
        RECT 23.030 135.480 23.470 136.520 ;
        RECT 23.740 135.480 24.220 136.520 ;
        RECT 23.165 134.750 23.335 135.250 ;
        RECT 24.625 134.125 24.875 137.625 ;
        RECT 21.625 133.875 24.875 134.125 ;
        RECT 21.625 130.375 21.875 133.875 ;
        RECT 23.165 133.000 23.335 133.500 ;
        RECT 22.280 131.730 22.760 132.770 ;
        RECT 23.030 131.730 23.470 132.770 ;
        RECT 23.740 131.730 24.220 132.770 ;
        RECT 23.165 131.000 23.335 131.500 ;
        RECT 24.625 130.375 24.875 133.875 ;
        RECT 21.625 130.125 24.875 130.375 ;
        RECT 21.625 126.625 21.875 130.125 ;
        RECT 23.165 129.250 23.335 129.750 ;
        RECT 22.280 127.980 22.760 129.020 ;
        RECT 23.030 127.980 23.470 129.020 ;
        RECT 23.740 127.980 24.220 129.020 ;
        RECT 23.165 127.250 23.335 127.750 ;
        RECT 24.625 126.625 24.875 130.125 ;
        RECT 21.625 126.375 24.875 126.625 ;
        RECT 21.625 122.875 21.875 126.375 ;
        RECT 23.165 125.500 23.335 126.000 ;
        RECT 22.280 124.230 22.760 125.270 ;
        RECT 23.030 124.230 23.470 125.270 ;
        RECT 23.740 124.230 24.220 125.270 ;
        RECT 23.165 123.500 23.335 124.000 ;
        RECT 24.625 122.875 24.875 126.375 ;
        RECT 21.625 122.625 24.875 122.875 ;
        RECT 21.625 119.125 21.875 122.625 ;
        RECT 23.165 121.750 23.335 122.250 ;
        RECT 22.280 120.480 22.760 121.520 ;
        RECT 23.030 120.480 23.470 121.520 ;
        RECT 23.740 120.480 24.220 121.520 ;
        RECT 23.165 119.750 23.335 120.250 ;
        RECT 24.625 119.125 24.875 122.625 ;
        RECT 21.625 118.875 24.875 119.125 ;
        RECT 21.625 115.375 21.875 118.875 ;
        RECT 23.165 118.000 23.335 118.500 ;
        RECT 22.280 116.730 22.760 117.770 ;
        RECT 23.030 116.730 23.470 117.770 ;
        RECT 23.740 116.730 24.220 117.770 ;
        RECT 23.165 116.000 23.335 116.500 ;
        RECT 24.625 115.375 24.875 118.875 ;
        RECT 21.625 115.125 24.875 115.375 ;
        RECT 21.625 111.625 21.875 115.125 ;
        RECT 23.165 114.250 23.335 114.750 ;
        RECT 22.280 112.980 22.760 114.020 ;
        RECT 23.030 112.980 23.470 114.020 ;
        RECT 23.740 112.980 24.220 114.020 ;
        RECT 23.165 112.250 23.335 112.750 ;
        RECT 24.625 111.625 24.875 115.125 ;
        RECT 21.625 111.375 24.875 111.625 ;
        RECT 31.125 141.375 34.375 141.625 ;
        RECT 31.125 137.875 31.375 141.375 ;
        RECT 32.665 140.500 32.835 141.000 ;
        RECT 31.780 139.230 32.260 140.270 ;
        RECT 32.530 139.230 32.970 140.270 ;
        RECT 33.240 139.230 33.720 140.270 ;
        RECT 32.665 138.500 32.835 139.000 ;
        RECT 34.125 137.875 34.375 141.375 ;
        RECT 31.125 137.625 34.375 137.875 ;
        RECT 31.125 134.125 31.375 137.625 ;
        RECT 32.665 136.750 32.835 137.250 ;
        RECT 31.780 135.480 32.260 136.520 ;
        RECT 32.530 135.480 32.970 136.520 ;
        RECT 33.240 135.480 33.720 136.520 ;
        RECT 32.665 134.750 32.835 135.250 ;
        RECT 34.125 134.125 34.375 137.625 ;
        RECT 31.125 133.875 34.375 134.125 ;
        RECT 31.125 130.375 31.375 133.875 ;
        RECT 32.665 133.000 32.835 133.500 ;
        RECT 31.780 131.730 32.260 132.770 ;
        RECT 32.530 131.730 32.970 132.770 ;
        RECT 33.240 131.730 33.720 132.770 ;
        RECT 32.665 131.000 32.835 131.500 ;
        RECT 34.125 130.375 34.375 133.875 ;
        RECT 31.125 130.125 34.375 130.375 ;
        RECT 31.125 126.625 31.375 130.125 ;
        RECT 32.665 129.250 32.835 129.750 ;
        RECT 31.780 127.980 32.260 129.020 ;
        RECT 32.530 127.980 32.970 129.020 ;
        RECT 33.240 127.980 33.720 129.020 ;
        RECT 32.665 127.250 32.835 127.750 ;
        RECT 34.125 126.625 34.375 130.125 ;
        RECT 31.125 126.375 34.375 126.625 ;
        RECT 31.125 122.875 31.375 126.375 ;
        RECT 32.665 125.500 32.835 126.000 ;
        RECT 31.780 124.230 32.260 125.270 ;
        RECT 32.530 124.230 32.970 125.270 ;
        RECT 33.240 124.230 33.720 125.270 ;
        RECT 32.665 123.500 32.835 124.000 ;
        RECT 34.125 122.875 34.375 126.375 ;
        RECT 31.125 122.625 34.375 122.875 ;
        RECT 31.125 119.125 31.375 122.625 ;
        RECT 32.665 121.750 32.835 122.250 ;
        RECT 31.780 120.480 32.260 121.520 ;
        RECT 32.530 120.480 32.970 121.520 ;
        RECT 33.240 120.480 33.720 121.520 ;
        RECT 32.665 119.750 32.835 120.250 ;
        RECT 34.125 119.125 34.375 122.625 ;
        RECT 31.125 118.875 34.375 119.125 ;
        RECT 31.125 115.375 31.375 118.875 ;
        RECT 32.665 118.000 32.835 118.500 ;
        RECT 31.780 116.730 32.260 117.770 ;
        RECT 32.530 116.730 32.970 117.770 ;
        RECT 33.240 116.730 33.720 117.770 ;
        RECT 32.665 116.000 32.835 116.500 ;
        RECT 34.125 115.375 34.375 118.875 ;
        RECT 31.125 115.125 34.375 115.375 ;
        RECT 31.125 111.625 31.375 115.125 ;
        RECT 32.665 114.250 32.835 114.750 ;
        RECT 31.780 112.980 32.260 114.020 ;
        RECT 32.530 112.980 32.970 114.020 ;
        RECT 33.240 112.980 33.720 114.020 ;
        RECT 32.665 112.250 32.835 112.750 ;
        RECT 34.125 111.625 34.375 115.125 ;
        RECT 31.125 111.375 34.375 111.625 ;
        RECT 40.625 141.375 43.875 141.625 ;
        RECT 40.625 137.875 40.875 141.375 ;
        RECT 42.165 140.500 42.335 141.000 ;
        RECT 41.280 139.230 41.760 140.270 ;
        RECT 42.030 139.230 42.470 140.270 ;
        RECT 42.740 139.230 43.220 140.270 ;
        RECT 42.165 138.500 42.335 139.000 ;
        RECT 43.625 137.875 43.875 141.375 ;
        RECT 114.685 141.045 115.895 142.135 ;
        RECT 116.525 142.135 117.275 142.655 ;
        RECT 117.445 142.305 118.195 142.825 ;
        RECT 118.835 142.855 119.235 143.045 ;
        RECT 119.955 143.025 120.145 143.425 ;
        RECT 119.405 142.855 120.145 143.025 ;
        RECT 116.525 141.045 118.195 142.135 ;
        RECT 118.375 141.045 118.665 142.015 ;
        RECT 118.835 141.215 119.065 142.855 ;
        RECT 119.405 142.685 119.575 142.855 ;
        RECT 119.235 141.990 119.575 142.685 ;
        RECT 119.745 142.270 120.070 142.685 ;
        RECT 120.520 142.355 120.900 143.315 ;
        RECT 121.085 143.115 121.415 143.595 ;
        RECT 121.090 142.355 121.405 142.930 ;
        RECT 122.045 142.825 125.555 143.595 ;
        RECT 125.725 142.870 126.015 143.595 ;
        RECT 126.185 142.825 128.775 143.595 ;
        RECT 128.965 143.110 129.755 143.375 ;
        RECT 122.045 142.135 123.735 142.655 ;
        RECT 123.905 142.305 125.555 142.825 ;
        RECT 119.235 141.760 120.070 141.990 ;
        RECT 119.235 141.045 119.565 141.460 ;
        RECT 119.755 141.215 120.070 141.760 ;
        RECT 120.240 141.745 121.355 142.010 ;
        RECT 120.240 141.215 120.465 141.745 ;
        RECT 120.635 141.045 120.965 141.555 ;
        RECT 121.135 141.215 121.355 141.745 ;
        RECT 122.045 141.045 125.555 142.135 ;
        RECT 125.725 141.045 126.015 142.210 ;
        RECT 126.185 142.135 127.395 142.655 ;
        RECT 127.565 142.305 128.775 142.825 ;
        RECT 128.945 142.435 129.330 142.915 ;
        RECT 129.500 142.255 129.755 143.110 ;
        RECT 129.925 142.930 130.155 143.375 ;
        RECT 130.335 143.100 130.665 143.595 ;
        RECT 130.840 142.965 131.090 143.425 ;
        RECT 129.925 142.435 130.335 142.930 ;
        RECT 130.920 142.755 131.090 142.965 ;
        RECT 131.260 142.935 131.535 143.595 ;
        RECT 132.185 143.085 132.425 143.595 ;
        RECT 132.595 143.085 132.885 143.425 ;
        RECT 133.115 143.085 133.430 143.595 ;
        RECT 130.520 142.255 130.750 142.685 ;
        RECT 126.185 141.045 128.775 142.135 ;
        RECT 128.960 142.085 130.750 142.255 ;
        RECT 130.920 142.235 131.535 142.755 ;
        RECT 132.225 142.745 132.425 142.915 ;
        RECT 132.230 142.355 132.425 142.745 ;
        RECT 128.960 141.720 129.215 142.085 ;
        RECT 129.385 141.725 129.715 141.915 ;
        RECT 129.940 141.790 130.190 142.085 ;
        RECT 129.385 141.550 129.575 141.725 ;
        RECT 128.945 141.045 129.575 141.550 ;
        RECT 129.755 141.215 130.230 141.555 ;
        RECT 130.415 141.045 130.630 141.890 ;
        RECT 130.935 141.885 131.105 142.235 ;
        RECT 132.595 142.185 132.775 143.085 ;
        RECT 133.600 143.025 133.770 143.295 ;
        RECT 133.940 143.195 134.270 143.595 ;
        RECT 132.945 142.355 133.355 142.915 ;
        RECT 133.600 142.855 134.295 143.025 ;
        RECT 133.525 142.185 133.695 142.685 ;
        RECT 130.830 141.215 131.105 141.885 ;
        RECT 131.275 141.045 131.535 142.055 ;
        RECT 132.235 142.015 133.695 142.185 ;
        RECT 132.235 141.840 132.595 142.015 ;
        RECT 133.865 141.845 134.295 142.855 ;
        RECT 134.925 142.825 137.515 143.595 ;
        RECT 137.685 142.845 138.895 143.595 ;
        RECT 133.180 141.045 133.350 141.845 ;
        RECT 133.520 141.675 134.295 141.845 ;
        RECT 134.925 142.135 136.135 142.655 ;
        RECT 136.305 142.305 137.515 142.825 ;
        RECT 137.685 142.135 138.205 142.675 ;
        RECT 138.375 142.305 138.895 142.845 ;
        RECT 133.520 141.215 133.850 141.675 ;
        RECT 134.020 141.045 134.190 141.505 ;
        RECT 134.925 141.045 137.515 142.135 ;
        RECT 137.685 141.045 138.895 142.135 ;
        RECT 114.600 140.875 138.980 141.045 ;
        RECT 114.685 139.785 115.895 140.875 ;
        RECT 114.685 139.075 115.205 139.615 ;
        RECT 115.375 139.245 115.895 139.785 ;
        RECT 116.065 139.785 117.735 140.875 ;
        RECT 116.065 139.265 116.815 139.785 ;
        RECT 117.910 139.725 118.170 140.875 ;
        RECT 118.345 139.800 118.600 140.705 ;
        RECT 118.770 140.115 119.100 140.875 ;
        RECT 119.315 139.945 119.485 140.705 ;
        RECT 116.985 139.095 117.735 139.615 ;
        RECT 114.685 138.325 115.895 139.075 ;
        RECT 116.065 138.325 117.735 139.095 ;
        RECT 117.910 138.325 118.170 139.165 ;
        RECT 118.345 139.070 118.515 139.800 ;
        RECT 118.770 139.775 119.485 139.945 ;
        RECT 119.745 139.785 120.955 140.875 ;
        RECT 121.130 140.440 126.475 140.875 ;
        RECT 126.650 140.440 131.995 140.875 ;
        RECT 132.170 140.440 137.515 140.875 ;
        RECT 118.770 139.565 118.940 139.775 ;
        RECT 118.685 139.235 118.940 139.565 ;
        RECT 118.345 138.495 118.600 139.070 ;
        RECT 118.770 139.045 118.940 139.235 ;
        RECT 119.220 139.225 119.575 139.595 ;
        RECT 119.745 139.245 120.265 139.785 ;
        RECT 120.435 139.075 120.955 139.615 ;
        RECT 122.720 139.190 123.070 140.440 ;
        RECT 118.770 138.875 119.485 139.045 ;
        RECT 118.770 138.325 119.100 138.705 ;
        RECT 119.315 138.495 119.485 138.875 ;
        RECT 119.745 138.325 120.955 139.075 ;
        RECT 124.550 138.870 124.890 139.700 ;
        RECT 128.240 139.190 128.590 140.440 ;
        RECT 130.070 138.870 130.410 139.700 ;
        RECT 133.760 139.190 134.110 140.440 ;
        RECT 137.685 139.785 138.895 140.875 ;
        RECT 135.590 138.870 135.930 139.700 ;
        RECT 137.685 139.245 138.205 139.785 ;
        RECT 138.375 139.075 138.895 139.615 ;
        RECT 121.130 138.325 126.475 138.870 ;
        RECT 126.650 138.325 131.995 138.870 ;
        RECT 132.170 138.325 137.515 138.870 ;
        RECT 137.685 138.325 138.895 139.075 ;
        RECT 114.600 138.155 138.980 138.325 ;
        RECT 40.625 137.625 43.875 137.875 ;
        RECT 40.625 134.125 40.875 137.625 ;
        RECT 42.165 136.750 42.335 137.250 ;
        RECT 41.280 135.480 41.760 136.520 ;
        RECT 42.030 135.480 42.470 136.520 ;
        RECT 42.740 135.480 43.220 136.520 ;
        RECT 42.165 134.750 42.335 135.250 ;
        RECT 43.625 134.125 43.875 137.625 ;
        RECT 114.685 137.405 115.895 138.155 ;
        RECT 116.065 137.405 117.275 138.155 ;
        RECT 117.625 137.775 117.955 138.155 ;
        RECT 118.125 137.605 118.315 137.985 ;
        RECT 118.485 137.795 118.815 138.155 ;
        RECT 114.685 136.865 115.205 137.405 ;
        RECT 115.375 136.695 115.895 137.235 ;
        RECT 114.685 135.605 115.895 136.695 ;
        RECT 116.065 136.695 116.585 137.235 ;
        RECT 116.755 136.865 117.275 137.405 ;
        RECT 117.915 137.415 118.315 137.605 ;
        RECT 119.035 137.585 119.225 137.985 ;
        RECT 118.485 137.415 119.225 137.585 ;
        RECT 116.065 135.605 117.275 136.695 ;
        RECT 117.455 135.605 117.745 136.575 ;
        RECT 117.915 135.775 118.145 137.415 ;
        RECT 118.485 137.245 118.655 137.415 ;
        RECT 118.315 136.550 118.655 137.245 ;
        RECT 118.825 136.830 119.150 137.245 ;
        RECT 119.600 136.915 119.980 137.875 ;
        RECT 120.165 137.675 120.495 138.155 ;
        RECT 120.170 136.915 120.485 137.490 ;
        RECT 120.665 137.405 121.875 138.155 ;
        RECT 120.665 136.695 121.185 137.235 ;
        RECT 121.355 136.865 121.875 137.405 ;
        RECT 122.045 137.385 125.555 138.155 ;
        RECT 125.725 137.430 126.015 138.155 ;
        RECT 126.650 137.610 131.995 138.155 ;
        RECT 132.625 137.775 132.955 138.155 ;
        RECT 122.045 136.695 123.735 137.215 ;
        RECT 123.905 136.865 125.555 137.385 ;
        RECT 118.315 136.320 119.150 136.550 ;
        RECT 118.315 135.605 118.645 136.020 ;
        RECT 118.835 135.775 119.150 136.320 ;
        RECT 119.320 136.305 120.435 136.570 ;
        RECT 119.320 135.775 119.545 136.305 ;
        RECT 119.715 135.605 120.045 136.115 ;
        RECT 120.215 135.775 120.435 136.305 ;
        RECT 120.665 135.605 121.875 136.695 ;
        RECT 122.045 135.605 125.555 136.695 ;
        RECT 125.725 135.605 126.015 136.770 ;
        RECT 128.240 136.040 128.590 137.290 ;
        RECT 130.070 136.780 130.410 137.610 ;
        RECT 132.180 137.605 132.455 137.745 ;
        RECT 133.125 137.605 133.335 137.775 ;
        RECT 132.180 137.415 133.335 137.605 ;
        RECT 133.505 137.605 133.835 137.985 ;
        RECT 134.025 137.775 134.355 138.155 ;
        RECT 133.505 137.400 134.355 137.605 ;
        RECT 132.175 136.790 132.435 137.245 ;
        RECT 132.690 136.840 133.275 137.215 ;
        RECT 126.650 135.605 131.995 136.040 ;
        RECT 132.180 135.605 132.505 136.590 ;
        RECT 132.690 136.455 132.895 136.840 ;
        RECT 133.445 136.625 133.855 137.230 ;
        RECT 134.025 136.910 134.355 137.400 ;
        RECT 134.025 136.455 134.195 136.910 ;
        RECT 132.685 136.285 132.895 136.455 ;
        RECT 132.690 136.255 132.895 136.285 ;
        RECT 133.075 136.235 134.195 136.455 ;
        RECT 133.075 135.775 133.335 136.235 ;
        RECT 133.505 135.605 134.355 136.055 ;
        RECT 134.525 135.775 134.770 137.985 ;
        RECT 134.955 137.355 135.195 138.155 ;
        RECT 135.845 137.385 137.515 138.155 ;
        RECT 137.685 137.405 138.895 138.155 ;
        RECT 135.845 136.695 136.595 137.215 ;
        RECT 136.765 136.865 137.515 137.385 ;
        RECT 137.685 136.695 138.205 137.235 ;
        RECT 138.375 136.865 138.895 137.405 ;
        RECT 134.955 135.605 135.210 136.605 ;
        RECT 135.845 135.605 137.515 136.695 ;
        RECT 137.685 135.605 138.895 136.695 ;
        RECT 114.600 135.435 138.980 135.605 ;
        RECT 114.685 134.345 115.895 135.435 ;
        RECT 116.990 135.000 122.335 135.435 ;
        RECT 122.510 135.000 127.855 135.435 ;
        RECT 128.030 135.000 133.375 135.435 ;
        RECT 40.625 133.875 43.875 134.125 ;
        RECT 40.625 130.375 40.875 133.875 ;
        RECT 42.165 133.000 42.335 133.500 ;
        RECT 41.280 131.730 41.760 132.770 ;
        RECT 42.030 131.730 42.470 132.770 ;
        RECT 42.740 131.730 43.220 132.770 ;
        RECT 42.165 131.000 42.335 131.500 ;
        RECT 43.625 130.375 43.875 133.875 ;
        RECT 114.685 133.635 115.205 134.175 ;
        RECT 115.375 133.805 115.895 134.345 ;
        RECT 118.580 133.750 118.930 135.000 ;
        RECT 114.685 132.885 115.895 133.635 ;
        RECT 120.410 133.430 120.750 134.260 ;
        RECT 124.100 133.750 124.450 135.000 ;
        RECT 125.930 133.430 126.270 134.260 ;
        RECT 129.620 133.750 129.970 135.000 ;
        RECT 131.450 133.430 131.790 134.260 ;
        RECT 133.545 134.230 133.835 135.435 ;
        RECT 134.005 134.295 134.280 135.265 ;
        RECT 134.490 134.635 134.770 135.435 ;
        RECT 134.940 134.925 136.135 135.215 ;
        RECT 134.950 134.585 136.115 134.755 ;
        RECT 134.950 134.465 135.120 134.585 ;
        RECT 134.450 134.295 135.120 134.465 ;
        RECT 116.990 132.885 122.335 133.430 ;
        RECT 122.510 132.885 127.855 133.430 ;
        RECT 128.030 132.885 133.375 133.430 ;
        RECT 133.545 132.885 133.835 133.715 ;
        RECT 134.005 133.560 134.175 134.295 ;
        RECT 134.450 134.125 134.620 134.295 ;
        RECT 135.390 134.125 135.615 134.415 ;
        RECT 135.785 134.295 136.115 134.585 ;
        RECT 136.305 134.345 137.515 135.435 ;
        RECT 137.685 134.345 138.895 135.435 ;
        RECT 134.345 133.795 134.620 134.125 ;
        RECT 134.790 133.795 135.615 134.125 ;
        RECT 135.785 133.795 136.135 134.125 ;
        RECT 136.305 133.805 136.825 134.345 ;
        RECT 134.450 133.625 134.620 133.795 ;
        RECT 136.995 133.635 137.515 134.175 ;
        RECT 137.685 133.805 138.205 134.345 ;
        RECT 138.375 133.635 138.895 134.175 ;
        RECT 134.005 133.215 134.280 133.560 ;
        RECT 134.450 133.455 136.115 133.625 ;
        RECT 134.470 132.885 134.850 133.285 ;
        RECT 135.020 133.105 135.190 133.455 ;
        RECT 135.360 132.885 135.690 133.285 ;
        RECT 135.860 133.105 136.115 133.455 ;
        RECT 136.305 132.885 137.515 133.635 ;
        RECT 137.685 132.885 138.895 133.635 ;
        RECT 114.600 132.715 138.980 132.885 ;
        RECT 114.685 131.965 115.895 132.715 ;
        RECT 114.685 131.425 115.205 131.965 ;
        RECT 116.065 131.945 117.735 132.715 ;
        RECT 115.375 131.255 115.895 131.795 ;
        RECT 40.625 130.125 43.875 130.375 ;
        RECT 114.685 130.165 115.895 131.255 ;
        RECT 116.065 131.255 116.815 131.775 ;
        RECT 116.985 131.425 117.735 131.945 ;
        RECT 117.925 131.915 118.165 132.715 ;
        RECT 116.065 130.165 117.735 131.255 ;
        RECT 117.910 130.165 118.165 131.165 ;
        RECT 118.350 130.335 118.595 132.545 ;
        RECT 118.765 132.335 119.095 132.715 ;
        RECT 119.285 132.165 119.615 132.545 ;
        RECT 120.165 132.335 120.495 132.715 ;
        RECT 118.765 131.960 119.615 132.165 ;
        RECT 119.785 132.165 119.995 132.335 ;
        RECT 120.665 132.165 120.940 132.305 ;
        RECT 119.785 131.975 120.940 132.165 ;
        RECT 118.765 131.470 119.095 131.960 ;
        RECT 122.045 131.945 125.555 132.715 ;
        RECT 125.725 131.990 126.015 132.715 ;
        RECT 127.105 131.945 130.615 132.715 ;
        RECT 130.810 132.315 131.140 132.715 ;
        RECT 131.310 132.145 131.480 132.415 ;
        RECT 131.650 132.205 131.965 132.715 ;
        RECT 132.195 132.205 132.485 132.545 ;
        RECT 132.655 132.205 132.895 132.715 ;
        RECT 133.085 132.235 133.345 132.715 ;
        RECT 133.515 132.465 133.760 132.545 ;
        RECT 133.515 132.295 133.845 132.465 ;
        RECT 118.925 131.015 119.095 131.470 ;
        RECT 119.265 131.185 119.675 131.790 ;
        RECT 119.845 131.400 120.430 131.775 ;
        RECT 120.225 131.015 120.430 131.400 ;
        RECT 120.685 131.350 120.945 131.805 ;
        RECT 122.045 131.255 123.735 131.775 ;
        RECT 123.905 131.425 125.555 131.945 ;
        RECT 118.925 130.795 120.045 131.015 ;
        RECT 120.225 130.845 120.435 131.015 ;
        RECT 120.225 130.815 120.430 130.845 ;
        RECT 118.765 130.165 119.615 130.615 ;
        RECT 119.785 130.335 120.045 130.795 ;
        RECT 120.615 130.165 120.940 131.150 ;
        RECT 122.045 130.165 125.555 131.255 ;
        RECT 125.725 130.165 126.015 131.330 ;
        RECT 127.105 131.255 128.795 131.775 ;
        RECT 128.965 131.425 130.615 131.945 ;
        RECT 130.785 131.975 131.480 132.145 ;
        RECT 127.105 130.165 130.615 131.255 ;
        RECT 130.785 130.965 131.215 131.975 ;
        RECT 131.385 131.305 131.555 131.805 ;
        RECT 131.725 131.475 132.135 132.035 ;
        RECT 132.305 131.305 132.485 132.205 ;
        RECT 132.655 131.695 132.850 132.035 ;
        RECT 132.655 131.525 132.855 131.695 ;
        RECT 132.655 131.475 132.850 131.525 ;
        RECT 133.130 131.475 133.325 132.045 ;
        RECT 133.515 131.305 133.685 132.295 ;
        RECT 134.045 132.100 134.255 132.385 ;
        RECT 134.520 132.375 134.690 132.400 ;
        RECT 134.520 132.205 134.695 132.375 ;
        RECT 134.935 132.335 135.265 132.715 ;
        RECT 135.035 132.255 135.205 132.335 ;
        RECT 134.520 132.105 134.690 132.205 ;
        RECT 133.865 131.930 134.255 132.100 ;
        RECT 134.425 131.935 134.690 132.105 ;
        RECT 135.455 132.085 135.625 132.545 ;
        RECT 135.875 132.255 136.130 132.715 ;
        RECT 133.865 131.475 134.035 131.930 ;
        RECT 134.425 131.725 134.595 131.935 ;
        RECT 134.950 131.805 135.155 132.040 ;
        RECT 135.455 131.915 136.130 132.085 ;
        RECT 136.305 131.965 137.515 132.715 ;
        RECT 137.685 131.965 138.895 132.715 ;
        RECT 134.265 131.555 134.595 131.725 ;
        RECT 134.425 131.540 134.595 131.555 ;
        RECT 134.825 131.475 135.155 131.805 ;
        RECT 135.335 131.555 135.665 131.725 ;
        RECT 135.495 131.305 135.665 131.555 ;
        RECT 131.385 131.135 132.845 131.305 ;
        RECT 130.785 130.795 131.560 130.965 ;
        RECT 130.890 130.165 131.060 130.625 ;
        RECT 131.230 130.335 131.560 130.795 ;
        RECT 131.730 130.165 131.900 130.965 ;
        RECT 132.485 130.960 132.845 131.135 ;
        RECT 133.175 131.135 135.665 131.305 ;
        RECT 133.175 130.335 133.345 131.135 ;
        RECT 135.875 130.965 136.130 131.915 ;
        RECT 133.575 130.795 134.865 130.965 ;
        RECT 133.635 130.375 133.885 130.795 ;
        RECT 134.075 130.165 134.405 130.625 ;
        RECT 134.615 130.375 134.865 130.795 ;
        RECT 135.035 130.165 135.285 130.965 ;
        RECT 135.455 130.795 136.130 130.965 ;
        RECT 136.305 131.255 136.825 131.795 ;
        RECT 136.995 131.425 137.515 131.965 ;
        RECT 137.685 131.255 138.205 131.795 ;
        RECT 138.375 131.425 138.895 131.965 ;
        RECT 135.455 130.335 135.625 130.795 ;
        RECT 135.835 130.165 136.085 130.625 ;
        RECT 136.305 130.165 137.515 131.255 ;
        RECT 137.685 130.165 138.895 131.255 ;
        RECT 40.625 126.625 40.875 130.125 ;
        RECT 42.165 129.250 42.335 129.750 ;
        RECT 41.280 127.980 41.760 129.020 ;
        RECT 42.030 127.980 42.470 129.020 ;
        RECT 42.740 127.980 43.220 129.020 ;
        RECT 42.165 127.250 42.335 127.750 ;
        RECT 43.625 126.625 43.875 130.125 ;
        RECT 114.600 129.995 138.980 130.165 ;
        RECT 114.685 128.905 115.895 129.995 ;
        RECT 114.685 128.195 115.205 128.735 ;
        RECT 115.375 128.365 115.895 128.905 ;
        RECT 116.065 128.905 117.275 129.995 ;
        RECT 117.495 129.535 117.745 129.995 ;
        RECT 117.955 129.365 118.125 129.825 ;
        RECT 117.450 129.195 118.125 129.365 ;
        RECT 118.295 129.195 118.545 129.995 ;
        RECT 118.715 129.365 118.965 129.785 ;
        RECT 119.175 129.535 119.505 129.995 ;
        RECT 119.695 129.365 119.945 129.785 ;
        RECT 118.715 129.195 120.005 129.365 ;
        RECT 116.065 128.365 116.585 128.905 ;
        RECT 116.755 128.195 117.275 128.735 ;
        RECT 114.685 127.445 115.895 128.195 ;
        RECT 116.065 127.445 117.275 128.195 ;
        RECT 117.450 128.245 117.705 129.195 ;
        RECT 120.235 129.025 120.405 129.825 ;
        RECT 120.670 129.560 126.015 129.995 ;
        RECT 126.190 129.560 131.535 129.995 ;
        RECT 117.915 128.855 120.405 129.025 ;
        RECT 117.915 128.605 118.085 128.855 ;
        RECT 117.915 128.435 118.245 128.605 ;
        RECT 118.425 128.355 118.755 128.685 ;
        RECT 118.985 128.605 119.155 128.620 ;
        RECT 118.985 128.435 119.315 128.605 ;
        RECT 117.450 128.075 118.125 128.245 ;
        RECT 118.425 128.120 118.630 128.355 ;
        RECT 118.985 128.225 119.155 128.435 ;
        RECT 119.545 128.230 119.715 128.685 ;
        RECT 117.450 127.445 117.705 127.905 ;
        RECT 117.955 127.615 118.125 128.075 ;
        RECT 118.890 128.055 119.155 128.225 ;
        RECT 119.325 128.060 119.715 128.230 ;
        RECT 118.890 127.955 119.060 128.055 ;
        RECT 118.375 127.825 118.545 127.905 ;
        RECT 118.315 127.445 118.645 127.825 ;
        RECT 118.885 127.785 119.060 127.955 ;
        RECT 118.890 127.760 119.060 127.785 ;
        RECT 119.325 127.775 119.535 128.060 ;
        RECT 119.895 127.865 120.065 128.855 ;
        RECT 120.255 128.115 120.450 128.685 ;
        RECT 122.260 128.310 122.610 129.560 ;
        RECT 124.090 127.990 124.430 128.820 ;
        RECT 127.780 128.310 128.130 129.560 ;
        RECT 131.905 129.325 132.185 129.995 ;
        RECT 129.610 127.990 129.950 128.820 ;
        RECT 131.705 128.685 132.020 129.125 ;
        RECT 132.355 129.105 132.655 129.655 ;
        RECT 132.865 129.275 133.195 129.995 ;
        RECT 133.385 129.275 133.835 129.825 ;
        RECT 132.355 128.935 133.295 129.105 ;
        RECT 133.125 128.685 133.295 128.935 ;
        RECT 131.705 128.435 132.395 128.685 ;
        RECT 132.625 128.435 132.955 128.685 ;
        RECT 133.125 128.355 133.415 128.685 ;
        RECT 133.125 128.265 133.295 128.355 ;
        RECT 131.905 128.075 133.295 128.265 ;
        RECT 119.735 127.695 120.065 127.865 ;
        RECT 119.820 127.615 120.065 127.695 ;
        RECT 120.235 127.445 120.495 127.925 ;
        RECT 120.670 127.445 126.015 127.990 ;
        RECT 126.190 127.445 131.535 127.990 ;
        RECT 131.905 127.715 132.235 128.075 ;
        RECT 133.585 127.905 133.835 129.275 ;
        RECT 134.005 128.855 134.295 129.995 ;
        RECT 134.925 128.905 137.515 129.995 ;
        RECT 137.685 128.905 138.895 129.995 ;
        RECT 134.925 128.385 136.135 128.905 ;
        RECT 132.865 127.445 133.115 127.905 ;
        RECT 133.285 127.615 133.835 127.905 ;
        RECT 134.005 127.445 134.295 128.245 ;
        RECT 136.305 128.215 137.515 128.735 ;
        RECT 137.685 128.365 138.205 128.905 ;
        RECT 134.925 127.445 137.515 128.215 ;
        RECT 138.375 128.195 138.895 128.735 ;
        RECT 137.685 127.445 138.895 128.195 ;
        RECT 114.600 127.275 138.980 127.445 ;
        RECT 40.625 126.375 43.875 126.625 ;
        RECT 40.625 122.875 40.875 126.375 ;
        RECT 42.165 125.500 42.335 126.000 ;
        RECT 41.280 124.230 41.760 125.270 ;
        RECT 42.030 124.230 42.470 125.270 ;
        RECT 42.740 124.230 43.220 125.270 ;
        RECT 42.165 123.500 42.335 124.000 ;
        RECT 43.625 122.875 43.875 126.375 ;
        RECT 114.685 126.525 115.895 127.275 ;
        RECT 114.685 125.985 115.205 126.525 ;
        RECT 116.525 126.505 120.035 127.275 ;
        RECT 120.210 126.730 125.555 127.275 ;
        RECT 115.375 125.815 115.895 126.355 ;
        RECT 114.685 124.725 115.895 125.815 ;
        RECT 116.525 125.815 118.215 126.335 ;
        RECT 118.385 125.985 120.035 126.505 ;
        RECT 116.525 124.725 120.035 125.815 ;
        RECT 121.800 125.160 122.150 126.410 ;
        RECT 123.630 125.900 123.970 126.730 ;
        RECT 125.725 126.550 126.015 127.275 ;
        RECT 126.650 126.730 131.995 127.275 ;
        RECT 132.170 126.730 137.515 127.275 ;
        RECT 120.210 124.725 125.555 125.160 ;
        RECT 125.725 124.725 126.015 125.890 ;
        RECT 128.240 125.160 128.590 126.410 ;
        RECT 130.070 125.900 130.410 126.730 ;
        RECT 133.760 125.160 134.110 126.410 ;
        RECT 135.590 125.900 135.930 126.730 ;
        RECT 137.685 126.525 138.895 127.275 ;
        RECT 137.685 125.815 138.205 126.355 ;
        RECT 138.375 125.985 138.895 126.525 ;
        RECT 126.650 124.725 131.995 125.160 ;
        RECT 132.170 124.725 137.515 125.160 ;
        RECT 137.685 124.725 138.895 125.815 ;
        RECT 114.600 124.555 138.980 124.725 ;
        RECT 40.625 122.625 43.875 122.875 ;
        RECT 40.625 119.125 40.875 122.625 ;
        RECT 42.165 121.750 42.335 122.250 ;
        RECT 41.280 120.480 41.760 121.520 ;
        RECT 42.030 120.480 42.470 121.520 ;
        RECT 42.740 120.480 43.220 121.520 ;
        RECT 42.165 119.750 42.335 120.250 ;
        RECT 43.625 119.125 43.875 122.625 ;
        RECT 40.625 118.875 43.875 119.125 ;
        RECT 88.375 123.375 106.125 123.625 ;
        RECT 88.375 119.125 88.625 123.375 ;
        RECT 89.055 120.870 89.225 121.910 ;
        RECT 89.495 120.870 89.665 121.910 ;
        RECT 89.935 120.870 90.105 121.910 ;
        RECT 90.375 120.870 90.545 121.910 ;
        RECT 90.815 120.870 90.985 121.910 ;
        RECT 91.465 120.870 91.635 121.910 ;
        RECT 91.905 120.870 92.075 121.910 ;
        RECT 92.345 120.870 92.515 121.910 ;
        RECT 92.785 120.870 92.955 121.910 ;
        RECT 93.225 120.870 93.395 121.910 ;
        RECT 93.875 120.870 94.045 121.910 ;
        RECT 94.315 120.870 94.485 121.910 ;
        RECT 94.755 120.870 94.925 121.910 ;
        RECT 95.195 120.870 95.365 121.910 ;
        RECT 95.635 120.870 95.805 121.910 ;
        RECT 96.285 120.870 96.455 121.910 ;
        RECT 96.725 120.870 96.895 121.910 ;
        RECT 97.165 120.870 97.335 121.910 ;
        RECT 97.605 120.870 97.775 121.910 ;
        RECT 98.045 120.870 98.215 121.910 ;
        RECT 98.695 120.870 98.865 121.910 ;
        RECT 99.135 120.870 99.305 121.910 ;
        RECT 99.575 120.870 99.745 121.910 ;
        RECT 100.015 120.870 100.185 121.910 ;
        RECT 100.455 120.870 100.625 121.910 ;
        RECT 101.105 120.870 101.275 121.910 ;
        RECT 101.545 120.870 101.715 121.910 ;
        RECT 101.985 120.870 102.155 121.910 ;
        RECT 102.425 120.870 102.595 121.910 ;
        RECT 102.865 120.870 103.035 121.910 ;
        RECT 103.515 120.870 103.685 121.910 ;
        RECT 103.955 120.870 104.125 121.910 ;
        RECT 104.395 120.870 104.565 121.910 ;
        RECT 104.835 120.870 105.005 121.910 ;
        RECT 105.275 120.870 105.445 121.910 ;
        RECT 89.855 119.560 90.185 119.940 ;
        RECT 92.265 119.560 92.595 119.940 ;
        RECT 94.675 119.560 95.005 119.940 ;
        RECT 97.085 119.560 97.415 119.940 ;
        RECT 99.495 119.560 99.825 119.940 ;
        RECT 101.905 119.560 102.235 119.940 ;
        RECT 104.315 119.560 104.645 119.940 ;
        RECT 105.875 119.125 106.125 123.375 ;
        RECT 88.375 118.875 106.125 119.125 ;
        RECT 40.625 115.375 40.875 118.875 ;
        RECT 42.165 118.000 42.335 118.500 ;
        RECT 41.280 116.730 41.760 117.770 ;
        RECT 42.030 116.730 42.470 117.770 ;
        RECT 42.740 116.730 43.220 117.770 ;
        RECT 42.165 116.000 42.335 116.500 ;
        RECT 43.625 115.375 43.875 118.875 ;
        RECT 40.625 115.125 43.875 115.375 ;
        RECT 40.625 111.625 40.875 115.125 ;
        RECT 42.165 114.250 42.335 114.750 ;
        RECT 41.280 112.980 41.760 114.020 ;
        RECT 42.030 112.980 42.470 114.020 ;
        RECT 42.740 112.980 43.220 114.020 ;
        RECT 42.165 112.250 42.335 112.750 ;
        RECT 43.625 111.625 43.875 115.125 ;
        RECT 76.375 118.375 82.625 118.625 ;
        RECT 76.375 115.125 76.625 118.375 ;
        RECT 77.835 117.530 78.165 117.970 ;
        RECT 77.425 116.230 77.865 117.270 ;
        RECT 78.135 116.230 78.575 117.270 ;
        RECT 77.835 115.530 78.165 115.970 ;
        RECT 79.375 115.125 79.625 118.375 ;
        RECT 80.835 117.530 81.165 117.970 ;
        RECT 80.425 116.230 80.865 117.270 ;
        RECT 81.135 116.230 81.575 117.270 ;
        RECT 80.835 115.530 81.165 115.970 ;
        RECT 82.375 115.125 82.625 118.375 ;
        RECT 76.375 114.875 82.625 115.125 ;
        RECT 88.375 115.125 106.125 115.375 ;
        RECT 40.625 111.375 43.875 111.625 ;
        RECT 88.375 110.125 88.625 115.125 ;
        RECT 89.855 114.310 90.185 114.690 ;
        RECT 92.265 114.310 92.595 114.690 ;
        RECT 94.675 114.310 95.005 114.690 ;
        RECT 97.085 114.310 97.415 114.690 ;
        RECT 99.495 114.310 99.825 114.690 ;
        RECT 101.905 114.310 102.235 114.690 ;
        RECT 104.315 114.310 104.645 114.690 ;
        RECT 89.055 111.340 89.225 113.380 ;
        RECT 89.495 111.340 89.665 113.380 ;
        RECT 89.935 111.340 90.105 113.380 ;
        RECT 90.375 111.340 90.545 113.380 ;
        RECT 90.815 111.340 90.985 113.380 ;
        RECT 91.465 111.340 91.635 113.380 ;
        RECT 91.905 111.340 92.075 113.380 ;
        RECT 92.345 111.340 92.515 113.380 ;
        RECT 92.785 111.340 92.955 113.380 ;
        RECT 93.225 111.340 93.395 113.380 ;
        RECT 93.875 111.340 94.045 113.380 ;
        RECT 94.315 111.340 94.485 113.380 ;
        RECT 94.755 111.340 94.925 113.380 ;
        RECT 95.195 111.340 95.365 113.380 ;
        RECT 95.635 111.340 95.805 113.380 ;
        RECT 96.285 111.340 96.455 113.380 ;
        RECT 96.725 111.340 96.895 113.380 ;
        RECT 97.165 111.340 97.335 113.380 ;
        RECT 97.605 111.340 97.775 113.380 ;
        RECT 98.045 111.340 98.215 113.380 ;
        RECT 98.695 111.340 98.865 113.380 ;
        RECT 99.135 111.340 99.305 113.380 ;
        RECT 99.575 111.340 99.745 113.380 ;
        RECT 100.015 111.340 100.185 113.380 ;
        RECT 100.455 111.340 100.625 113.380 ;
        RECT 101.105 111.340 101.275 113.380 ;
        RECT 101.545 111.340 101.715 113.380 ;
        RECT 101.985 111.340 102.155 113.380 ;
        RECT 102.425 111.340 102.595 113.380 ;
        RECT 102.865 111.340 103.035 113.380 ;
        RECT 103.515 111.340 103.685 113.380 ;
        RECT 103.955 111.340 104.125 113.380 ;
        RECT 104.395 111.340 104.565 113.380 ;
        RECT 104.835 111.340 105.005 113.380 ;
        RECT 105.275 111.340 105.445 113.380 ;
        RECT 105.875 110.125 106.125 115.125 ;
        RECT 88.375 109.875 106.125 110.125 ;
      LAYER met1 ;
        RECT 0.000 200.000 147.500 204.000 ;
        RECT 5.000 195.000 147.500 199.000 ;
        RECT 81.500 194.500 82.500 195.000 ;
        RECT 137.000 194.500 138.000 195.000 ;
        RECT 81.500 194.000 138.000 194.500 ;
        RECT 20.750 188.500 49.250 189.500 ;
        RECT 21.000 187.750 25.500 188.500 ;
        RECT 21.000 184.500 22.000 187.750 ;
        RECT 22.250 186.500 22.750 187.000 ;
        RECT 23.000 186.750 23.500 187.250 ;
        RECT 23.750 186.500 24.250 187.000 ;
        RECT 22.250 185.500 22.790 186.500 ;
        RECT 23.000 185.500 23.500 186.500 ;
        RECT 23.710 185.500 24.250 186.500 ;
        RECT 23.000 184.750 23.500 185.250 ;
        RECT 24.500 184.500 25.500 187.750 ;
        RECT 21.000 184.000 25.500 184.500 ;
        RECT 21.000 180.750 22.000 184.000 ;
        RECT 22.250 182.750 22.750 183.250 ;
        RECT 23.000 183.000 23.500 183.500 ;
        RECT 23.750 182.750 24.250 183.250 ;
        RECT 22.250 181.750 22.790 182.750 ;
        RECT 23.000 181.750 23.500 182.750 ;
        RECT 23.710 181.750 24.250 182.750 ;
        RECT 23.000 181.000 23.500 181.500 ;
        RECT 24.500 180.750 25.500 184.000 ;
        RECT 21.000 180.250 25.500 180.750 ;
        RECT 21.000 177.000 22.000 180.250 ;
        RECT 22.250 179.000 22.750 179.500 ;
        RECT 23.000 179.250 23.500 179.750 ;
        RECT 23.750 179.000 24.250 179.500 ;
        RECT 22.250 178.000 22.790 179.000 ;
        RECT 23.000 178.000 23.500 179.000 ;
        RECT 23.710 178.000 24.250 179.000 ;
        RECT 23.000 177.250 23.500 177.750 ;
        RECT 24.500 177.000 25.500 180.250 ;
        RECT 21.000 176.500 25.500 177.000 ;
        RECT 21.000 173.250 22.000 176.500 ;
        RECT 22.250 175.250 22.750 175.750 ;
        RECT 23.000 175.500 23.500 176.000 ;
        RECT 23.750 175.250 24.250 175.750 ;
        RECT 22.250 174.250 22.790 175.250 ;
        RECT 23.000 174.250 23.500 175.250 ;
        RECT 23.710 174.250 24.250 175.250 ;
        RECT 23.000 173.500 23.500 174.000 ;
        RECT 24.500 173.250 25.500 176.500 ;
        RECT 21.000 172.750 25.500 173.250 ;
        RECT 21.000 169.500 22.000 172.750 ;
        RECT 22.250 171.500 22.750 172.000 ;
        RECT 23.000 171.750 23.500 172.250 ;
        RECT 23.750 171.500 24.250 172.000 ;
        RECT 22.250 170.500 22.790 171.500 ;
        RECT 23.000 170.500 23.500 171.500 ;
        RECT 23.710 170.500 24.250 171.500 ;
        RECT 23.000 169.750 23.500 170.250 ;
        RECT 24.500 169.500 25.500 172.750 ;
        RECT 21.000 169.000 25.500 169.500 ;
        RECT 21.000 165.750 22.000 169.000 ;
        RECT 22.250 167.750 22.750 168.250 ;
        RECT 23.000 168.000 23.500 168.500 ;
        RECT 23.750 167.750 24.250 168.250 ;
        RECT 22.250 166.750 22.790 167.750 ;
        RECT 23.000 166.750 23.500 167.750 ;
        RECT 23.710 166.750 24.250 167.750 ;
        RECT 23.000 166.000 23.500 166.500 ;
        RECT 24.500 165.750 25.500 169.000 ;
        RECT 21.000 165.250 25.500 165.750 ;
        RECT 21.000 162.000 22.000 165.250 ;
        RECT 22.250 164.000 22.750 164.500 ;
        RECT 23.000 164.250 23.500 164.750 ;
        RECT 23.750 164.000 24.250 164.500 ;
        RECT 22.250 163.000 22.790 164.000 ;
        RECT 23.000 163.000 23.500 164.000 ;
        RECT 23.710 163.000 24.250 164.000 ;
        RECT 23.000 162.250 23.500 162.750 ;
        RECT 24.500 162.000 25.500 165.250 ;
        RECT 21.000 161.500 25.500 162.000 ;
        RECT 21.000 158.250 22.000 161.500 ;
        RECT 22.250 160.250 22.750 160.750 ;
        RECT 23.000 160.500 23.500 161.000 ;
        RECT 23.750 160.250 24.250 160.750 ;
        RECT 22.250 159.250 22.790 160.250 ;
        RECT 23.000 159.250 23.500 160.250 ;
        RECT 23.710 159.250 24.250 160.250 ;
        RECT 23.000 158.500 23.500 159.000 ;
        RECT 24.500 158.250 25.500 161.500 ;
        RECT 21.000 157.500 25.500 158.250 ;
        RECT 30.500 187.750 35.000 188.500 ;
        RECT 30.500 184.500 31.500 187.750 ;
        RECT 31.750 186.500 32.250 187.000 ;
        RECT 32.500 186.750 33.000 187.250 ;
        RECT 33.250 186.500 33.750 187.000 ;
        RECT 31.750 185.500 32.290 186.500 ;
        RECT 32.500 185.500 33.000 186.500 ;
        RECT 33.210 185.500 33.750 186.500 ;
        RECT 32.500 184.750 33.000 185.250 ;
        RECT 34.000 184.500 35.000 187.750 ;
        RECT 30.500 184.000 35.000 184.500 ;
        RECT 30.500 180.750 31.500 184.000 ;
        RECT 31.750 182.750 32.250 183.250 ;
        RECT 32.500 183.000 33.000 183.500 ;
        RECT 33.250 182.750 33.750 183.250 ;
        RECT 31.750 181.750 32.290 182.750 ;
        RECT 32.500 181.750 33.000 182.750 ;
        RECT 33.210 181.750 33.750 182.750 ;
        RECT 32.500 181.000 33.000 181.500 ;
        RECT 34.000 180.750 35.000 184.000 ;
        RECT 30.500 180.250 35.000 180.750 ;
        RECT 30.500 177.000 31.500 180.250 ;
        RECT 31.750 179.000 32.250 179.500 ;
        RECT 32.500 179.250 33.000 179.750 ;
        RECT 33.250 179.000 33.750 179.500 ;
        RECT 31.750 178.000 32.290 179.000 ;
        RECT 32.500 178.000 33.000 179.000 ;
        RECT 33.210 178.000 33.750 179.000 ;
        RECT 32.500 177.250 33.000 177.750 ;
        RECT 34.000 177.000 35.000 180.250 ;
        RECT 30.500 176.500 35.000 177.000 ;
        RECT 30.500 173.250 31.500 176.500 ;
        RECT 31.750 175.250 32.250 175.750 ;
        RECT 32.500 175.500 33.000 176.000 ;
        RECT 33.250 175.250 33.750 175.750 ;
        RECT 31.750 174.250 32.290 175.250 ;
        RECT 32.500 174.250 33.000 175.250 ;
        RECT 33.210 174.250 33.750 175.250 ;
        RECT 32.500 173.500 33.000 174.000 ;
        RECT 34.000 173.250 35.000 176.500 ;
        RECT 30.500 172.750 35.000 173.250 ;
        RECT 30.500 169.500 31.500 172.750 ;
        RECT 31.750 171.500 32.250 172.000 ;
        RECT 32.500 171.750 33.000 172.250 ;
        RECT 33.250 171.500 33.750 172.000 ;
        RECT 31.750 170.500 32.290 171.500 ;
        RECT 32.500 170.500 33.000 171.500 ;
        RECT 33.210 170.500 33.750 171.500 ;
        RECT 32.500 169.750 33.000 170.250 ;
        RECT 34.000 169.500 35.000 172.750 ;
        RECT 30.500 169.000 35.000 169.500 ;
        RECT 30.500 165.750 31.500 169.000 ;
        RECT 31.750 167.750 32.250 168.250 ;
        RECT 32.500 168.000 33.000 168.500 ;
        RECT 33.250 167.750 33.750 168.250 ;
        RECT 31.750 166.750 32.290 167.750 ;
        RECT 32.500 166.750 33.000 167.750 ;
        RECT 33.210 166.750 33.750 167.750 ;
        RECT 32.500 166.000 33.000 166.500 ;
        RECT 34.000 165.750 35.000 169.000 ;
        RECT 30.500 165.250 35.000 165.750 ;
        RECT 30.500 162.000 31.500 165.250 ;
        RECT 31.750 164.000 32.250 164.500 ;
        RECT 32.500 164.250 33.000 164.750 ;
        RECT 33.250 164.000 33.750 164.500 ;
        RECT 31.750 163.000 32.290 164.000 ;
        RECT 32.500 163.000 33.000 164.000 ;
        RECT 33.210 163.000 33.750 164.000 ;
        RECT 32.500 162.250 33.000 162.750 ;
        RECT 34.000 162.000 35.000 165.250 ;
        RECT 30.500 161.500 35.000 162.000 ;
        RECT 30.500 158.250 31.500 161.500 ;
        RECT 31.750 160.250 32.250 160.750 ;
        RECT 32.500 160.500 33.000 161.000 ;
        RECT 33.250 160.250 33.750 160.750 ;
        RECT 31.750 159.250 32.290 160.250 ;
        RECT 32.500 159.250 33.000 160.250 ;
        RECT 33.210 159.250 33.750 160.250 ;
        RECT 32.500 158.500 33.000 159.000 ;
        RECT 34.000 158.250 35.000 161.500 ;
        RECT 30.500 157.500 35.000 158.250 ;
        RECT 40.000 187.750 44.500 188.500 ;
        RECT 40.000 184.500 41.000 187.750 ;
        RECT 41.250 186.500 41.750 187.000 ;
        RECT 42.000 186.750 42.500 187.250 ;
        RECT 42.750 186.500 43.250 187.000 ;
        RECT 41.250 185.500 41.790 186.500 ;
        RECT 42.000 185.500 42.500 186.500 ;
        RECT 42.710 185.500 43.250 186.500 ;
        RECT 42.000 184.750 42.500 185.250 ;
        RECT 43.500 184.500 44.500 187.750 ;
        RECT 81.500 188.250 82.500 194.000 ;
        RECT 89.370 193.585 92.280 193.815 ;
        RECT 95.870 193.585 98.780 193.815 ;
        RECT 107.120 193.585 110.030 193.815 ;
        RECT 111.870 193.585 114.780 193.815 ;
        RECT 120.870 193.585 123.780 193.815 ;
        RECT 127.870 193.585 130.780 193.815 ;
        RECT 88.280 192.750 88.510 193.405 ;
        RECT 88.720 192.955 88.950 193.405 ;
        RECT 94.780 192.750 95.010 193.405 ;
        RECT 95.220 192.955 95.450 193.405 ;
        RECT 100.270 192.955 100.725 193.405 ;
        RECT 101.770 192.955 102.225 193.405 ;
        RECT 103.270 192.955 103.725 193.405 ;
        RECT 100.270 192.750 100.500 192.955 ;
        RECT 101.770 192.750 102.000 192.955 ;
        RECT 103.270 192.750 103.500 192.955 ;
        RECT 106.030 192.750 106.260 193.405 ;
        RECT 106.470 192.955 106.700 193.405 ;
        RECT 110.780 192.750 111.010 193.405 ;
        RECT 111.220 192.955 111.450 193.405 ;
        RECT 116.270 192.955 116.725 193.405 ;
        RECT 116.270 192.750 116.500 192.955 ;
        RECT 119.780 192.750 120.010 193.405 ;
        RECT 120.220 192.955 120.450 193.405 ;
        RECT 126.780 192.750 127.010 193.405 ;
        RECT 127.220 192.955 127.450 193.405 ;
        RECT 132.270 192.955 132.725 193.405 ;
        RECT 132.270 192.750 132.500 192.955 ;
        RECT 88.000 192.250 88.510 192.750 ;
        RECT 88.650 192.365 91.940 192.595 ;
        RECT 88.280 191.105 88.510 192.250 ;
        RECT 94.250 192.000 95.010 192.750 ;
        RECT 98.000 192.250 100.500 192.750 ;
        RECT 100.750 192.250 101.250 192.750 ;
        RECT 101.500 192.250 102.000 192.750 ;
        RECT 102.250 192.250 103.500 192.750 ;
        RECT 103.750 192.250 106.260 192.750 ;
        RECT 106.400 192.365 109.690 192.595 ;
        RECT 100.270 192.005 100.500 192.250 ;
        RECT 101.770 192.005 102.000 192.250 ;
        RECT 103.270 192.005 103.500 192.250 ;
        RECT 91.500 191.500 95.010 192.000 ;
        RECT 98.000 191.500 98.660 192.000 ;
        RECT 94.780 191.105 95.010 191.500 ;
        RECT 100.270 191.105 100.725 192.005 ;
        RECT 101.770 191.105 102.225 192.005 ;
        RECT 103.270 191.105 103.725 192.005 ;
        RECT 106.030 191.105 106.260 192.250 ;
        RECT 110.250 192.000 111.010 192.750 ;
        RECT 114.000 192.250 116.500 192.750 ;
        RECT 116.750 192.250 117.250 192.750 ;
        RECT 119.500 192.250 120.010 192.750 ;
        RECT 120.150 192.365 123.440 192.595 ;
        RECT 126.250 192.250 127.010 192.750 ;
        RECT 130.000 192.250 132.500 192.750 ;
        RECT 132.750 192.250 133.250 192.750 ;
        RECT 116.270 192.005 116.500 192.250 ;
        RECT 109.250 191.500 111.010 192.000 ;
        RECT 114.000 191.500 114.660 192.000 ;
        RECT 110.780 191.105 111.010 191.500 ;
        RECT 116.270 191.105 116.725 192.005 ;
        RECT 119.780 191.105 120.010 192.250 ;
        RECT 123.750 192.000 124.750 192.250 ;
        RECT 122.500 191.500 124.750 192.000 ;
        RECT 123.750 191.250 124.750 191.500 ;
        RECT 126.780 191.105 127.010 192.250 ;
        RECT 132.270 192.005 132.500 192.250 ;
        RECT 130.000 191.500 130.660 192.000 ;
        RECT 132.270 191.105 132.725 192.005 ;
        RECT 90.090 190.670 92.280 190.900 ;
        RECT 96.590 190.670 98.780 190.900 ;
        RECT 107.840 190.670 110.030 190.900 ;
        RECT 112.590 190.670 114.780 190.900 ;
        RECT 121.590 190.670 123.780 190.900 ;
        RECT 128.590 190.670 130.780 190.900 ;
        RECT 84.500 190.000 136.500 190.500 ;
        RECT 88.000 189.250 94.000 189.750 ;
        RECT 94.250 189.250 101.250 189.750 ;
        RECT 101.500 189.250 110.000 189.750 ;
        RECT 110.250 189.250 117.250 189.750 ;
        RECT 118.750 189.250 133.250 189.750 ;
        RECT 86.000 188.500 100.500 189.000 ;
        RECT 102.000 188.500 116.500 189.000 ;
        RECT 118.000 188.500 132.500 189.000 ;
        RECT 137.000 188.250 138.000 194.000 ;
        RECT 81.500 187.750 138.000 188.250 ;
        RECT 40.000 184.000 44.500 184.500 ;
        RECT 50.250 184.000 58.500 184.500 ;
        RECT 40.000 180.750 41.000 184.000 ;
        RECT 41.250 182.750 41.750 183.250 ;
        RECT 42.000 183.000 42.500 183.500 ;
        RECT 42.750 182.750 43.250 183.250 ;
        RECT 41.250 181.750 41.790 182.750 ;
        RECT 42.000 181.750 42.500 182.750 ;
        RECT 42.710 181.750 43.250 182.750 ;
        RECT 42.000 181.000 42.500 181.500 ;
        RECT 43.500 180.750 44.500 184.000 ;
        RECT 81.500 182.500 82.500 187.750 ;
        RECT 87.370 187.335 90.280 187.565 ;
        RECT 98.370 187.335 101.280 187.565 ;
        RECT 103.370 187.335 106.280 187.565 ;
        RECT 114.370 187.335 117.280 187.565 ;
        RECT 119.370 187.335 122.280 187.565 ;
        RECT 130.370 187.335 133.280 187.565 ;
        RECT 86.280 186.500 86.510 187.155 ;
        RECT 86.720 186.705 86.950 187.155 ;
        RECT 86.000 186.000 86.510 186.500 ;
        RECT 86.280 184.855 86.510 186.000 ;
        RECT 88.250 185.750 88.750 187.335 ;
        RECT 91.500 186.545 93.000 187.000 ;
        RECT 94.000 186.545 94.750 187.000 ;
        RECT 90.850 186.500 93.000 186.545 ;
        RECT 89.500 186.175 90.000 186.500 ;
        RECT 90.850 186.315 92.000 186.500 ;
        RECT 89.500 185.945 91.250 186.175 ;
        RECT 88.250 185.250 90.500 185.750 ;
        RECT 90.750 185.500 91.250 185.945 ;
        RECT 91.500 185.500 92.000 186.145 ;
        RECT 92.500 186.000 93.000 186.500 ;
        RECT 93.350 186.500 94.750 186.545 ;
        RECT 95.270 186.705 95.725 187.155 ;
        RECT 95.270 186.500 95.500 186.705 ;
        RECT 97.280 186.500 97.510 187.155 ;
        RECT 97.720 186.705 97.950 187.155 ;
        RECT 93.350 186.315 94.500 186.500 ;
        RECT 93.250 186.000 93.750 186.145 ;
        RECT 92.500 185.500 93.750 186.000 ;
        RECT 94.000 186.000 94.500 186.145 ;
        RECT 95.000 186.000 95.500 186.500 ;
        RECT 95.750 186.000 97.510 186.500 ;
        RECT 94.000 185.755 95.500 186.000 ;
        RECT 94.000 185.500 95.725 185.755 ;
        RECT 88.250 184.650 88.750 185.250 ;
        RECT 90.860 184.855 91.090 185.500 ;
        RECT 93.360 184.855 93.590 185.500 ;
        RECT 95.270 184.855 95.725 185.500 ;
        RECT 97.280 184.855 97.510 186.000 ;
        RECT 99.250 185.750 99.750 187.335 ;
        RECT 102.280 186.500 102.510 187.155 ;
        RECT 102.720 186.705 102.950 187.155 ;
        RECT 100.000 186.000 101.000 186.500 ;
        RECT 102.000 186.000 102.510 186.500 ;
        RECT 97.750 185.250 101.160 185.750 ;
        RECT 99.250 184.650 99.750 185.250 ;
        RECT 102.280 184.855 102.510 186.000 ;
        RECT 104.250 185.750 104.750 187.335 ;
        RECT 107.500 186.545 109.000 187.000 ;
        RECT 110.000 186.545 110.750 187.000 ;
        RECT 106.850 186.500 109.000 186.545 ;
        RECT 105.500 186.175 106.000 186.500 ;
        RECT 106.850 186.315 108.000 186.500 ;
        RECT 105.500 185.945 107.250 186.175 ;
        RECT 104.250 185.250 106.500 185.750 ;
        RECT 106.750 185.500 107.250 185.945 ;
        RECT 107.500 185.500 108.000 186.145 ;
        RECT 108.500 186.000 109.000 186.500 ;
        RECT 109.350 186.500 110.750 186.545 ;
        RECT 111.270 186.705 111.725 187.155 ;
        RECT 111.270 186.500 111.500 186.705 ;
        RECT 113.280 186.500 113.510 187.155 ;
        RECT 113.720 186.705 113.950 187.155 ;
        RECT 109.350 186.315 110.500 186.500 ;
        RECT 109.250 186.000 109.750 186.145 ;
        RECT 108.500 185.500 109.750 186.000 ;
        RECT 110.000 186.000 110.500 186.145 ;
        RECT 111.000 186.000 111.500 186.500 ;
        RECT 111.750 186.000 113.510 186.500 ;
        RECT 110.000 185.755 111.500 186.000 ;
        RECT 110.000 185.500 111.725 185.755 ;
        RECT 104.250 184.650 104.750 185.250 ;
        RECT 106.860 184.855 107.090 185.500 ;
        RECT 109.360 184.855 109.590 185.500 ;
        RECT 111.270 184.855 111.725 185.500 ;
        RECT 113.280 184.855 113.510 186.000 ;
        RECT 115.250 185.750 115.750 187.335 ;
        RECT 118.280 186.500 118.510 187.155 ;
        RECT 118.720 186.705 118.950 187.155 ;
        RECT 116.000 186.000 117.000 186.500 ;
        RECT 118.000 186.000 118.510 186.500 ;
        RECT 113.750 185.250 117.160 185.750 ;
        RECT 115.250 184.650 115.750 185.250 ;
        RECT 118.280 184.855 118.510 186.000 ;
        RECT 120.250 185.750 120.750 187.335 ;
        RECT 123.500 186.545 125.000 187.000 ;
        RECT 126.000 186.545 126.750 187.000 ;
        RECT 122.850 186.500 125.000 186.545 ;
        RECT 121.500 186.175 122.000 186.500 ;
        RECT 122.850 186.315 124.000 186.500 ;
        RECT 121.500 185.945 123.250 186.175 ;
        RECT 120.250 185.250 122.500 185.750 ;
        RECT 122.750 185.500 123.250 185.945 ;
        RECT 123.500 185.500 124.000 186.145 ;
        RECT 124.500 186.000 125.000 186.500 ;
        RECT 125.350 186.500 126.750 186.545 ;
        RECT 127.270 186.705 127.725 187.155 ;
        RECT 127.270 186.500 127.500 186.705 ;
        RECT 129.280 186.500 129.510 187.155 ;
        RECT 129.720 186.705 129.950 187.155 ;
        RECT 125.350 186.315 126.500 186.500 ;
        RECT 125.250 186.000 125.750 186.145 ;
        RECT 124.500 185.500 125.750 186.000 ;
        RECT 126.000 186.000 126.500 186.145 ;
        RECT 127.000 186.000 127.500 186.500 ;
        RECT 127.750 186.000 129.510 186.500 ;
        RECT 126.000 185.755 127.500 186.000 ;
        RECT 126.000 185.500 127.725 185.755 ;
        RECT 120.250 184.650 120.750 185.250 ;
        RECT 122.860 184.855 123.090 185.500 ;
        RECT 125.360 184.855 125.590 185.500 ;
        RECT 127.270 184.855 127.725 185.500 ;
        RECT 129.280 184.855 129.510 186.000 ;
        RECT 131.250 185.750 131.750 187.335 ;
        RECT 132.000 186.000 133.000 186.500 ;
        RECT 129.750 185.250 133.160 185.750 ;
        RECT 131.250 184.650 131.750 185.250 ;
        RECT 88.090 184.420 90.280 184.650 ;
        RECT 99.090 184.420 101.280 184.650 ;
        RECT 104.090 184.420 106.280 184.650 ;
        RECT 115.090 184.420 117.280 184.650 ;
        RECT 120.090 184.420 122.280 184.650 ;
        RECT 131.090 184.420 133.280 184.650 ;
        RECT 84.500 183.750 136.500 184.250 ;
        RECT 90.000 183.000 104.250 183.500 ;
        RECT 106.000 183.000 119.250 183.500 ;
        RECT 119.500 183.000 130.250 183.500 ;
        RECT 137.000 182.500 138.000 187.750 ;
        RECT 81.500 181.500 138.000 182.500 ;
        RECT 40.000 180.250 44.500 180.750 ;
        RECT 50.250 180.250 60.500 180.750 ;
        RECT 77.250 180.500 146.000 181.500 ;
        RECT 40.000 177.000 41.000 180.250 ;
        RECT 41.250 179.000 41.750 179.500 ;
        RECT 42.000 179.250 42.500 179.750 ;
        RECT 42.750 179.000 43.250 179.500 ;
        RECT 41.250 178.000 41.790 179.000 ;
        RECT 42.000 178.000 42.500 179.000 ;
        RECT 42.710 178.000 43.250 179.000 ;
        RECT 42.000 177.250 42.500 177.750 ;
        RECT 43.500 177.000 44.500 180.250 ;
        RECT 77.250 178.000 78.250 180.500 ;
        RECT 103.500 179.750 116.250 180.250 ;
        RECT 95.000 179.000 105.500 179.500 ;
        RECT 108.000 179.000 115.500 179.500 ;
        RECT 91.250 178.250 99.250 178.750 ;
        RECT 104.250 178.250 112.250 178.750 ;
        RECT 145.000 178.000 146.000 180.500 ;
        RECT 77.250 177.500 146.000 178.000 ;
        RECT 40.000 176.500 44.500 177.000 ;
        RECT 50.250 176.500 62.500 177.000 ;
        RECT 40.000 173.250 41.000 176.500 ;
        RECT 41.250 175.250 41.750 175.750 ;
        RECT 42.000 175.500 42.500 176.000 ;
        RECT 42.750 175.250 43.250 175.750 ;
        RECT 41.250 174.250 41.790 175.250 ;
        RECT 42.000 174.250 42.500 175.250 ;
        RECT 42.710 174.250 43.250 175.250 ;
        RECT 42.000 173.500 42.500 174.000 ;
        RECT 43.500 173.250 44.500 176.500 ;
        RECT 40.000 172.750 44.500 173.250 ;
        RECT 50.250 172.750 64.500 173.250 ;
        RECT 40.000 169.500 41.000 172.750 ;
        RECT 41.250 171.500 41.750 172.000 ;
        RECT 42.000 171.750 42.500 172.250 ;
        RECT 42.750 171.500 43.250 172.000 ;
        RECT 41.250 170.500 41.790 171.500 ;
        RECT 42.000 170.500 42.500 171.500 ;
        RECT 42.710 170.500 43.250 171.500 ;
        RECT 42.000 169.750 42.500 170.250 ;
        RECT 43.500 169.500 44.500 172.750 ;
        RECT 77.250 171.000 78.250 177.500 ;
        RECT 90.500 177.130 94.400 177.360 ;
        RECT 99.435 177.130 101.175 177.360 ;
        RECT 104.100 177.130 107.400 177.360 ;
        RECT 112.435 177.130 114.175 177.360 ;
        RECT 81.520 176.455 81.975 176.905 ;
        RECT 84.020 176.455 84.475 176.905 ;
        RECT 85.520 176.455 85.975 176.905 ;
        RECT 81.520 176.250 81.750 176.455 ;
        RECT 84.020 176.250 84.250 176.455 ;
        RECT 85.520 176.250 85.750 176.455 ;
        RECT 86.970 176.250 87.250 176.905 ;
        RECT 88.770 176.750 89.225 176.905 ;
        RECT 81.250 175.750 81.750 176.250 ;
        RECT 82.000 175.750 84.250 176.250 ;
        RECT 84.500 175.750 85.750 176.250 ;
        RECT 86.000 175.750 87.250 176.250 ;
        RECT 87.600 176.455 89.225 176.750 ;
        RECT 90.500 176.750 91.250 177.130 ;
        RECT 92.470 177.100 93.030 177.130 ;
        RECT 87.600 176.065 89.000 176.455 ;
        RECT 81.520 175.505 81.750 175.750 ;
        RECT 84.020 175.505 84.250 175.750 ;
        RECT 85.520 175.505 85.750 175.750 ;
        RECT 87.020 175.505 87.250 175.750 ;
        RECT 81.520 175.500 81.975 175.505 ;
        RECT 81.250 174.500 82.250 175.500 ;
        RECT 84.020 174.605 84.475 175.505 ;
        RECT 85.520 174.605 85.975 175.505 ;
        RECT 87.020 174.605 87.600 175.505 ;
        RECT 87.750 175.250 88.250 175.925 ;
        RECT 88.500 175.750 89.000 176.065 ;
        RECT 89.250 175.750 89.750 176.250 ;
        RECT 88.770 175.505 89.000 175.750 ;
        RECT 88.770 174.605 89.225 175.505 ;
        RECT 90.500 175.500 91.000 176.750 ;
        RECT 91.480 176.685 91.710 176.905 ;
        RECT 92.760 176.685 92.990 176.905 ;
        RECT 91.480 176.455 92.520 176.685 ;
        RECT 92.760 176.455 94.480 176.685 ;
        RECT 91.250 175.750 91.750 176.250 ;
        RECT 92.750 176.080 93.980 176.310 ;
        RECT 95.000 176.250 95.230 176.905 ;
        RECT 97.525 176.455 97.980 176.905 ;
        RECT 97.750 176.250 97.980 176.455 ;
        RECT 98.750 176.265 99.250 176.750 ;
        RECT 99.435 176.455 99.665 177.130 ;
        RECT 100.345 176.760 102.225 176.990 ;
        RECT 101.995 176.455 102.225 176.760 ;
        RECT 104.480 176.685 104.710 176.905 ;
        RECT 105.760 176.685 105.990 176.905 ;
        RECT 104.480 176.455 105.520 176.685 ;
        RECT 105.760 176.455 107.480 176.685 ;
        RECT 92.750 175.680 92.980 176.080 ;
        RECT 95.000 175.980 95.500 176.250 ;
        RECT 97.000 175.980 97.500 176.250 ;
        RECT 93.190 175.710 94.860 175.940 ;
        RECT 95.000 175.750 97.500 175.980 ;
        RECT 97.750 175.895 98.250 176.250 ;
        RECT 98.750 176.035 101.915 176.265 ;
        RECT 90.500 175.230 93.000 175.500 ;
        RECT 90.500 175.000 94.210 175.230 ;
        RECT 91.000 174.370 91.750 174.750 ;
        RECT 92.340 174.370 92.570 174.800 ;
        RECT 91.000 174.250 93.360 174.370 ;
        RECT 91.250 174.140 93.360 174.250 ;
        RECT 93.980 174.140 94.210 175.000 ;
        RECT 95.000 174.605 95.230 175.750 ;
        RECT 97.730 175.665 100.545 175.895 ;
        RECT 100.750 175.750 101.250 176.035 ;
        RECT 102.250 175.895 104.000 176.250 ;
        RECT 101.435 175.750 104.000 175.895 ;
        RECT 104.250 175.750 104.750 176.250 ;
        RECT 105.750 176.080 106.980 176.310 ;
        RECT 108.000 176.250 108.230 176.905 ;
        RECT 110.525 176.455 110.980 176.905 ;
        RECT 110.750 176.250 110.980 176.455 ;
        RECT 111.750 176.265 112.250 176.750 ;
        RECT 112.435 176.455 112.665 177.130 ;
        RECT 113.345 176.760 115.225 176.990 ;
        RECT 114.995 176.455 115.225 176.760 ;
        RECT 117.500 176.730 118.000 177.000 ;
        RECT 118.170 176.925 119.450 177.155 ;
        RECT 133.600 177.130 136.900 177.360 ;
        RECT 117.500 176.500 118.650 176.730 ;
        RECT 101.435 175.665 102.750 175.750 ;
        RECT 105.750 175.680 105.980 176.080 ;
        RECT 108.000 175.980 108.500 176.250 ;
        RECT 110.000 175.980 110.500 176.250 ;
        RECT 106.190 175.710 107.860 175.940 ;
        RECT 108.000 175.750 110.500 175.980 ;
        RECT 110.750 175.895 111.250 176.250 ;
        RECT 111.750 176.035 114.915 176.265 ;
        RECT 97.750 175.505 97.980 175.665 ;
        RECT 97.525 174.605 97.980 175.505 ;
        RECT 98.750 175.250 99.250 175.665 ;
        RECT 99.395 174.370 99.625 175.505 ;
        RECT 101.435 175.340 101.895 175.665 ;
        RECT 100.685 174.880 101.895 175.340 ;
        RECT 100.245 174.510 101.415 174.740 ;
        RECT 102.035 174.370 102.265 175.505 ;
        RECT 104.100 175.230 105.500 175.500 ;
        RECT 104.100 175.000 107.210 175.230 ;
        RECT 99.395 174.140 100.515 174.370 ;
        RECT 100.965 174.140 102.265 174.370 ;
        RECT 104.000 174.370 104.750 174.750 ;
        RECT 105.340 174.370 105.570 174.800 ;
        RECT 104.000 174.250 106.360 174.370 ;
        RECT 104.250 174.140 106.360 174.250 ;
        RECT 106.980 174.140 107.210 175.000 ;
        RECT 108.000 174.605 108.230 175.750 ;
        RECT 110.730 175.665 113.545 175.895 ;
        RECT 113.750 175.750 114.250 176.035 ;
        RECT 115.250 175.895 116.000 176.250 ;
        RECT 114.435 175.665 116.000 175.895 ;
        RECT 116.500 175.750 118.000 176.250 ;
        RECT 117.480 175.695 118.000 175.750 ;
        RECT 110.750 175.505 110.980 175.665 ;
        RECT 110.525 174.605 110.980 175.505 ;
        RECT 111.750 175.250 112.250 175.665 ;
        RECT 112.395 174.370 112.625 175.505 ;
        RECT 114.435 175.340 114.895 175.665 ;
        RECT 113.685 174.880 114.895 175.340 ;
        RECT 113.245 174.510 114.415 174.740 ;
        RECT 115.035 174.370 115.265 175.505 ;
        RECT 115.500 175.500 116.000 175.665 ;
        RECT 115.500 175.230 118.000 175.500 ;
        RECT 118.790 175.230 119.020 176.665 ;
        RECT 119.220 175.635 119.450 176.925 ;
        RECT 119.590 176.250 119.820 176.905 ;
        RECT 122.025 176.455 122.480 176.905 ;
        RECT 123.775 176.455 124.230 176.905 ;
        RECT 125.525 176.455 125.980 176.905 ;
        RECT 127.275 176.455 127.730 176.905 ;
        RECT 129.775 176.750 130.230 176.905 ;
        RECT 129.775 176.455 131.500 176.750 ;
        RECT 122.250 176.250 122.480 176.455 ;
        RECT 124.000 176.250 124.230 176.455 ;
        RECT 125.750 176.250 125.980 176.455 ;
        RECT 127.500 176.250 127.730 176.455 ;
        RECT 130.000 176.250 131.500 176.455 ;
        RECT 119.590 175.750 122.000 176.250 ;
        RECT 122.250 175.750 123.750 176.250 ;
        RECT 124.000 175.750 125.500 176.250 ;
        RECT 125.750 175.750 127.250 176.250 ;
        RECT 127.500 175.750 129.750 176.250 ;
        RECT 130.000 175.750 130.500 176.250 ;
        RECT 131.000 176.065 131.500 176.250 ;
        RECT 131.640 175.935 131.870 176.905 ;
        RECT 132.420 176.250 132.650 176.905 ;
        RECT 133.980 176.685 134.210 176.905 ;
        RECT 135.260 176.685 135.490 176.905 ;
        RECT 133.980 176.455 135.020 176.685 ;
        RECT 135.260 176.455 136.980 176.685 ;
        RECT 115.500 175.000 119.020 175.230 ;
        RECT 112.395 174.140 113.515 174.370 ;
        RECT 113.965 174.140 115.265 174.370 ;
        RECT 115.750 174.250 118.110 174.750 ;
        RECT 118.790 174.370 119.020 175.000 ;
        RECT 119.590 174.605 119.820 175.750 ;
        RECT 122.250 175.505 122.480 175.750 ;
        RECT 124.000 175.505 124.500 175.750 ;
        RECT 125.750 175.505 125.980 175.750 ;
        RECT 127.500 175.505 127.730 175.750 ;
        RECT 130.000 175.505 130.230 175.750 ;
        RECT 122.025 174.605 122.480 175.505 ;
        RECT 123.775 174.605 124.500 175.505 ;
        RECT 125.525 174.605 125.980 175.505 ;
        RECT 127.275 174.605 127.730 175.505 ;
        RECT 129.775 174.605 130.230 175.505 ;
        RECT 117.500 174.140 118.110 174.250 ;
        RECT 118.660 174.140 119.020 174.370 ;
        RECT 124.000 174.465 124.500 174.605 ;
        RECT 131.000 174.465 131.500 175.910 ;
        RECT 131.640 175.705 132.110 175.935 ;
        RECT 132.250 175.750 133.500 176.250 ;
        RECT 133.750 175.750 134.250 176.250 ;
        RECT 135.250 176.080 136.480 176.310 ;
        RECT 137.500 176.250 137.730 176.905 ;
        RECT 131.640 174.605 131.870 175.705 ;
        RECT 132.420 174.605 132.650 175.750 ;
        RECT 135.250 175.680 135.480 176.080 ;
        RECT 135.690 175.710 137.360 175.940 ;
        RECT 137.500 175.750 138.500 176.250 ;
        RECT 133.600 175.230 136.250 175.500 ;
        RECT 133.600 175.000 136.710 175.230 ;
        RECT 134.840 174.750 135.070 174.800 ;
        RECT 124.000 174.235 131.500 174.465 ;
        RECT 133.750 174.370 135.070 174.750 ;
        RECT 133.750 174.140 135.860 174.370 ;
        RECT 136.480 174.140 136.710 175.000 ;
        RECT 137.500 174.605 137.730 175.750 ;
        RECT 78.500 173.500 139.750 174.000 ;
        RECT 83.750 172.750 88.250 173.250 ;
        RECT 88.500 172.750 89.750 173.250 ;
        RECT 91.000 172.750 104.500 173.250 ;
        RECT 104.750 172.750 117.000 173.250 ;
        RECT 122.750 172.750 135.000 173.250 ;
        RECT 97.000 172.000 99.500 172.500 ;
        RECT 102.000 172.000 112.500 172.500 ;
        RECT 124.000 172.000 134.250 172.500 ;
        RECT 83.000 171.250 88.000 171.750 ;
        RECT 95.250 171.250 103.250 171.750 ;
        RECT 108.250 171.250 116.250 171.750 ;
        RECT 116.750 171.250 138.000 171.750 ;
        RECT 145.000 171.000 146.000 177.500 ;
        RECT 77.250 170.500 146.000 171.000 ;
        RECT 40.000 169.000 44.500 169.500 ;
        RECT 50.250 169.000 66.500 169.500 ;
        RECT 40.000 165.750 41.000 169.000 ;
        RECT 41.250 167.750 41.750 168.250 ;
        RECT 42.000 168.000 42.500 168.500 ;
        RECT 42.750 167.750 43.250 168.250 ;
        RECT 41.250 166.750 41.790 167.750 ;
        RECT 42.000 166.750 42.500 167.750 ;
        RECT 42.710 166.750 43.250 167.750 ;
        RECT 42.000 166.000 42.500 166.500 ;
        RECT 43.500 165.750 44.500 169.000 ;
        RECT 40.000 165.250 44.500 165.750 ;
        RECT 50.250 165.250 68.500 165.750 ;
        RECT 40.000 162.000 41.000 165.250 ;
        RECT 41.250 164.000 41.750 164.500 ;
        RECT 42.000 164.250 42.500 164.750 ;
        RECT 42.750 164.000 43.250 164.500 ;
        RECT 41.250 163.000 41.790 164.000 ;
        RECT 42.000 163.000 42.500 164.000 ;
        RECT 42.710 163.000 43.250 164.000 ;
        RECT 42.000 162.250 42.500 162.750 ;
        RECT 43.500 162.000 44.500 165.250 ;
        RECT 77.250 164.000 78.250 170.500 ;
        RECT 93.325 170.130 95.065 170.360 ;
        RECT 100.100 170.130 103.400 170.360 ;
        RECT 106.325 170.130 108.065 170.360 ;
        RECT 113.100 170.130 116.400 170.360 ;
        RECT 81.520 169.455 81.975 169.905 ;
        RECT 84.020 169.455 84.475 169.905 ;
        RECT 85.520 169.455 85.975 169.905 ;
        RECT 81.520 169.250 81.750 169.455 ;
        RECT 84.020 169.250 84.250 169.455 ;
        RECT 85.520 169.250 85.750 169.455 ;
        RECT 86.970 169.250 87.250 169.905 ;
        RECT 92.275 169.760 94.155 169.990 ;
        RECT 87.500 169.250 88.250 169.750 ;
        RECT 92.275 169.455 92.505 169.760 ;
        RECT 94.835 169.455 95.065 170.130 ;
        RECT 95.250 169.265 95.750 169.750 ;
        RECT 81.250 168.750 81.750 169.250 ;
        RECT 82.000 168.750 84.250 169.250 ;
        RECT 84.500 168.750 85.750 169.250 ;
        RECT 86.000 168.750 87.250 169.250 ;
        RECT 87.600 169.065 88.250 169.250 ;
        RECT 81.520 168.505 81.750 168.750 ;
        RECT 84.020 168.505 84.250 168.750 ;
        RECT 85.520 168.505 85.750 168.750 ;
        RECT 87.020 168.505 87.250 168.750 ;
        RECT 87.750 168.750 88.250 168.925 ;
        RECT 91.750 168.895 92.250 169.250 ;
        RECT 92.585 169.035 95.750 169.265 ;
        RECT 96.520 169.455 96.975 169.905 ;
        RECT 96.520 169.250 96.750 169.455 ;
        RECT 99.270 169.250 99.500 169.905 ;
        RECT 101.510 169.685 101.740 169.905 ;
        RECT 102.790 169.685 103.020 169.905 ;
        RECT 100.020 169.455 101.740 169.685 ;
        RECT 101.980 169.455 103.020 169.685 ;
        RECT 105.275 169.760 107.155 169.990 ;
        RECT 105.275 169.455 105.505 169.760 ;
        RECT 107.835 169.455 108.065 170.130 ;
        RECT 81.520 168.500 81.975 168.505 ;
        RECT 81.520 167.605 83.750 168.500 ;
        RECT 84.020 167.605 84.475 168.505 ;
        RECT 85.520 167.605 85.975 168.505 ;
        RECT 87.020 167.605 87.600 168.505 ;
        RECT 87.750 168.250 89.750 168.750 ;
        RECT 91.750 168.665 93.065 168.895 ;
        RECT 93.250 168.750 93.750 169.035 ;
        RECT 96.250 168.895 96.750 169.250 ;
        RECT 97.000 168.980 97.500 169.250 ;
        RECT 99.000 168.980 99.500 169.250 ;
        RECT 100.520 169.080 101.750 169.310 ;
        RECT 108.250 169.265 108.750 169.750 ;
        RECT 93.955 168.665 96.770 168.895 ;
        RECT 97.000 168.750 99.500 168.980 ;
        RECT 82.750 167.500 83.750 167.605 ;
        RECT 92.235 167.370 92.465 168.505 ;
        RECT 92.605 168.340 93.065 168.665 ;
        RECT 92.605 167.880 93.815 168.340 ;
        RECT 93.085 167.510 94.255 167.740 ;
        RECT 94.875 167.370 95.105 168.505 ;
        RECT 95.250 168.250 95.750 168.665 ;
        RECT 96.520 168.505 96.750 168.665 ;
        RECT 96.520 167.605 96.975 168.505 ;
        RECT 99.270 167.605 99.500 168.750 ;
        RECT 99.640 168.710 101.310 168.940 ;
        RECT 101.520 168.680 101.750 169.080 ;
        RECT 102.750 168.750 103.250 169.250 ;
        RECT 104.750 168.895 105.250 169.250 ;
        RECT 105.585 169.035 108.750 169.265 ;
        RECT 109.520 169.455 109.975 169.905 ;
        RECT 109.520 169.250 109.750 169.455 ;
        RECT 112.270 169.250 112.500 169.905 ;
        RECT 114.510 169.685 114.740 169.905 ;
        RECT 115.790 169.685 116.020 169.905 ;
        RECT 113.020 169.455 114.740 169.685 ;
        RECT 114.980 169.455 116.020 169.685 ;
        RECT 122.025 169.455 122.480 169.905 ;
        RECT 123.775 169.455 124.230 169.905 ;
        RECT 125.525 169.455 125.980 169.905 ;
        RECT 127.275 169.455 127.730 169.905 ;
        RECT 129.775 169.750 130.230 169.905 ;
        RECT 129.775 169.455 131.500 169.750 ;
        RECT 104.750 168.665 106.065 168.895 ;
        RECT 106.250 168.750 106.750 169.035 ;
        RECT 109.250 168.895 109.750 169.250 ;
        RECT 110.000 168.980 110.500 169.250 ;
        RECT 112.000 168.980 112.500 169.250 ;
        RECT 113.520 169.080 114.750 169.310 ;
        RECT 122.250 169.250 122.480 169.455 ;
        RECT 124.000 169.250 124.230 169.455 ;
        RECT 125.750 169.250 125.980 169.455 ;
        RECT 127.500 169.250 127.730 169.455 ;
        RECT 130.000 169.250 131.500 169.455 ;
        RECT 106.955 168.665 109.770 168.895 ;
        RECT 110.000 168.750 112.500 168.980 ;
        RECT 102.000 168.230 103.400 168.500 ;
        RECT 100.290 168.000 103.400 168.230 ;
        RECT 92.235 167.140 93.535 167.370 ;
        RECT 93.985 167.140 95.105 167.370 ;
        RECT 100.290 167.140 100.520 168.000 ;
        RECT 101.930 167.370 102.160 167.800 ;
        RECT 102.750 167.370 103.500 167.750 ;
        RECT 101.140 167.250 103.500 167.370 ;
        RECT 105.235 167.370 105.465 168.505 ;
        RECT 105.605 168.340 106.065 168.665 ;
        RECT 105.605 167.880 106.815 168.340 ;
        RECT 106.085 167.510 107.255 167.740 ;
        RECT 107.875 167.370 108.105 168.505 ;
        RECT 108.250 168.250 108.750 168.665 ;
        RECT 109.520 168.505 109.750 168.665 ;
        RECT 109.520 167.605 109.975 168.505 ;
        RECT 112.270 167.605 112.500 168.750 ;
        RECT 112.640 168.710 114.310 168.940 ;
        RECT 114.520 168.680 114.750 169.080 ;
        RECT 115.750 168.750 116.250 169.250 ;
        RECT 120.000 168.750 122.000 169.250 ;
        RECT 122.250 168.750 123.750 169.250 ;
        RECT 124.000 168.750 125.500 169.250 ;
        RECT 125.750 168.750 127.250 169.250 ;
        RECT 127.500 168.750 129.750 169.250 ;
        RECT 130.000 168.750 130.500 169.250 ;
        RECT 131.000 169.065 131.500 169.250 ;
        RECT 131.640 168.935 131.870 169.905 ;
        RECT 132.420 169.750 132.650 169.905 ;
        RECT 134.690 169.890 135.460 170.120 ;
        RECT 132.420 169.250 134.750 169.750 ;
        RECT 122.250 168.505 122.480 168.750 ;
        RECT 124.000 168.505 124.500 168.750 ;
        RECT 125.750 168.505 125.980 168.750 ;
        RECT 127.500 168.505 127.730 168.750 ;
        RECT 130.000 168.505 130.230 168.750 ;
        RECT 115.000 168.230 116.400 168.500 ;
        RECT 113.290 168.000 116.400 168.230 ;
        RECT 101.140 167.140 103.250 167.250 ;
        RECT 105.235 167.140 106.535 167.370 ;
        RECT 106.985 167.140 108.105 167.370 ;
        RECT 113.290 167.140 113.520 168.000 ;
        RECT 114.930 167.370 115.160 167.800 ;
        RECT 115.750 167.370 116.500 167.750 ;
        RECT 122.025 167.605 122.480 168.505 ;
        RECT 123.775 167.605 124.500 168.505 ;
        RECT 125.525 167.605 125.980 168.505 ;
        RECT 127.275 167.605 127.730 168.505 ;
        RECT 129.775 167.605 130.230 168.505 ;
        RECT 114.140 167.250 116.500 167.370 ;
        RECT 124.000 167.465 124.500 167.605 ;
        RECT 131.000 167.465 131.500 168.910 ;
        RECT 131.640 168.705 132.110 168.935 ;
        RECT 132.250 168.750 132.750 169.250 ;
        RECT 134.250 169.065 134.750 169.250 ;
        RECT 135.230 169.025 135.460 169.890 ;
        RECT 135.600 169.455 135.980 169.905 ;
        RECT 137.275 169.455 137.730 169.905 ;
        RECT 135.750 169.250 135.980 169.455 ;
        RECT 137.500 169.250 137.730 169.455 ;
        RECT 134.250 168.750 134.750 168.895 ;
        RECT 131.640 167.605 131.870 168.705 ;
        RECT 132.420 167.605 132.650 168.750 ;
        RECT 133.000 168.250 134.750 168.750 ;
        RECT 135.230 168.710 135.610 169.025 ;
        RECT 135.750 168.750 136.250 169.250 ;
        RECT 136.500 168.750 137.250 169.250 ;
        RECT 137.500 168.750 138.000 169.250 ;
        RECT 135.230 168.110 135.460 168.710 ;
        RECT 135.750 168.505 135.980 168.750 ;
        RECT 137.500 168.505 137.730 168.750 ;
        RECT 134.290 167.880 135.460 168.110 ;
        RECT 135.600 167.605 135.980 168.505 ;
        RECT 137.275 167.605 137.730 168.505 ;
        RECT 114.140 167.140 116.250 167.250 ;
        RECT 124.000 167.235 131.500 167.465 ;
        RECT 78.500 166.500 139.750 167.000 ;
        RECT 103.000 165.750 117.250 166.250 ;
        RECT 91.750 165.000 118.000 165.500 ;
        RECT 131.750 165.000 138.000 165.500 ;
        RECT 108.500 164.250 122.000 164.750 ;
        RECT 123.750 164.250 138.250 164.750 ;
        RECT 145.000 164.000 146.000 170.500 ;
        RECT 77.250 163.500 146.000 164.000 ;
        RECT 40.000 161.500 44.500 162.000 ;
        RECT 50.250 161.500 70.500 162.000 ;
        RECT 40.000 158.250 41.000 161.500 ;
        RECT 41.250 160.250 41.750 160.750 ;
        RECT 42.000 160.500 42.500 161.000 ;
        RECT 42.750 160.250 43.250 160.750 ;
        RECT 41.250 159.250 41.790 160.250 ;
        RECT 42.000 159.250 42.500 160.250 ;
        RECT 42.710 159.250 43.250 160.250 ;
        RECT 42.000 158.500 42.500 159.000 ;
        RECT 43.500 158.250 44.500 161.500 ;
        RECT 40.000 157.500 44.500 158.250 ;
        RECT 50.250 157.750 72.500 158.250 ;
        RECT 20.750 156.500 53.000 157.500 ;
        RECT 77.250 157.000 78.250 163.500 ;
        RECT 93.620 163.085 96.530 163.315 ;
        RECT 99.370 163.085 102.280 163.315 ;
        RECT 104.370 163.085 107.280 163.315 ;
        RECT 111.870 163.085 114.780 163.315 ;
        RECT 120.120 163.085 123.030 163.315 ;
        RECT 125.120 163.085 128.030 163.315 ;
        RECT 136.120 163.085 139.030 163.315 ;
        RECT 141.120 163.085 144.030 163.315 ;
        RECT 86.750 162.905 89.000 163.000 ;
        RECT 86.750 162.455 89.225 162.905 ;
        RECT 90.520 162.455 90.975 162.905 ;
        RECT 86.750 161.505 89.000 162.455 ;
        RECT 90.520 162.250 90.750 162.455 ;
        RECT 92.530 162.250 92.760 162.905 ;
        RECT 92.970 162.455 93.200 162.905 ;
        RECT 98.280 162.250 98.510 162.905 ;
        RECT 98.720 162.455 98.950 162.905 ;
        RECT 103.280 162.250 103.510 162.905 ;
        RECT 103.720 162.455 103.950 162.905 ;
        RECT 108.770 162.455 109.225 162.905 ;
        RECT 108.770 162.250 109.000 162.455 ;
        RECT 110.780 162.250 111.010 162.905 ;
        RECT 111.220 162.455 111.450 162.905 ;
        RECT 89.250 161.750 90.750 162.250 ;
        RECT 91.000 161.750 92.760 162.250 ;
        RECT 92.900 161.865 96.190 162.095 ;
        RECT 90.520 161.505 90.750 161.750 ;
        RECT 86.750 160.605 89.225 161.505 ;
        RECT 90.520 160.605 90.975 161.505 ;
        RECT 91.250 161.000 92.760 161.750 ;
        RECT 98.000 161.500 98.510 162.250 ;
        RECT 98.650 161.865 101.940 162.095 ;
        RECT 103.000 161.500 103.510 162.250 ;
        RECT 103.650 161.865 106.940 162.095 ;
        RECT 108.500 161.505 109.000 162.250 ;
        RECT 109.250 161.750 111.010 162.250 ;
        RECT 108.500 161.500 109.225 161.505 ;
        RECT 95.750 161.000 98.510 161.500 ;
        RECT 101.500 161.000 103.510 161.500 ;
        RECT 106.500 161.000 109.225 161.500 ;
        RECT 92.530 160.605 92.760 161.000 ;
        RECT 98.280 160.605 98.510 161.000 ;
        RECT 103.280 160.605 103.510 161.000 ;
        RECT 108.770 160.605 109.225 161.000 ;
        RECT 110.780 160.605 111.010 161.750 ;
        RECT 112.500 161.500 113.000 163.085 ;
        RECT 115.600 162.250 115.830 162.905 ;
        RECT 114.000 161.750 116.000 162.250 ;
        RECT 116.380 161.935 116.610 162.905 ;
        RECT 119.030 162.750 119.260 162.905 ;
        RECT 116.750 162.250 119.260 162.750 ;
        RECT 119.470 162.455 119.700 162.905 ;
        RECT 116.750 162.065 117.250 162.250 ;
        RECT 112.500 161.000 114.660 161.500 ;
        RECT 86.750 160.500 89.000 160.605 ;
        RECT 112.500 160.400 113.000 161.000 ;
        RECT 115.600 160.605 115.830 161.750 ;
        RECT 116.140 161.705 116.610 161.935 ;
        RECT 116.380 160.605 116.610 161.705 ;
        RECT 116.750 161.250 117.250 161.910 ;
        RECT 118.750 161.750 119.260 162.250 ;
        RECT 119.030 160.605 119.260 161.750 ;
        RECT 120.750 161.500 121.250 163.085 ;
        RECT 124.030 162.250 124.260 162.905 ;
        RECT 124.470 162.455 124.700 162.905 ;
        RECT 121.500 161.750 122.750 162.250 ;
        RECT 123.750 161.500 124.260 162.250 ;
        RECT 120.750 161.000 124.260 161.500 ;
        RECT 120.750 160.400 121.250 161.000 ;
        RECT 124.030 160.605 124.260 161.000 ;
        RECT 126.000 161.500 126.500 163.085 ;
        RECT 129.250 162.295 130.750 162.750 ;
        RECT 131.750 162.295 132.250 162.750 ;
        RECT 128.600 162.250 130.750 162.295 ;
        RECT 127.250 161.925 127.750 162.250 ;
        RECT 128.600 162.065 129.750 162.250 ;
        RECT 127.250 161.695 129.000 161.925 ;
        RECT 126.000 161.000 128.250 161.500 ;
        RECT 128.500 161.250 129.000 161.695 ;
        RECT 129.250 161.250 129.750 161.895 ;
        RECT 130.250 161.750 130.750 162.250 ;
        RECT 131.100 162.065 132.250 162.295 ;
        RECT 133.020 162.455 133.475 162.905 ;
        RECT 133.020 162.250 133.250 162.455 ;
        RECT 135.030 162.250 135.260 162.905 ;
        RECT 135.470 162.455 135.700 162.905 ;
        RECT 131.000 161.750 131.500 161.895 ;
        RECT 130.250 161.250 131.500 161.750 ;
        RECT 131.750 161.750 132.250 161.895 ;
        RECT 132.750 161.750 133.250 162.250 ;
        RECT 133.500 161.750 135.260 162.250 ;
        RECT 131.750 161.505 133.250 161.750 ;
        RECT 131.750 161.250 133.475 161.505 ;
        RECT 126.000 160.400 126.500 161.000 ;
        RECT 128.610 160.605 128.840 161.250 ;
        RECT 131.110 160.605 131.340 161.250 ;
        RECT 133.020 160.605 133.475 161.250 ;
        RECT 135.030 160.605 135.260 161.750 ;
        RECT 137.000 161.500 137.500 163.085 ;
        RECT 139.750 162.905 140.250 163.000 ;
        RECT 137.750 161.750 138.750 162.250 ;
        RECT 139.750 161.500 140.260 162.905 ;
        RECT 140.470 162.455 140.700 162.905 ;
        RECT 140.400 161.865 143.690 162.095 ;
        RECT 135.500 161.000 140.260 161.500 ;
        RECT 137.000 160.750 140.260 161.000 ;
        RECT 137.000 160.400 137.500 160.750 ;
        RECT 139.750 160.605 140.260 160.750 ;
        RECT 141.250 161.000 144.250 161.500 ;
        RECT 139.750 160.500 140.250 160.605 ;
        RECT 141.250 160.400 142.500 161.000 ;
        RECT 94.340 160.170 96.530 160.400 ;
        RECT 100.090 160.170 102.280 160.400 ;
        RECT 105.090 160.170 107.280 160.400 ;
        RECT 112.500 160.250 114.780 160.400 ;
        RECT 120.750 160.250 123.030 160.400 ;
        RECT 112.590 160.170 114.780 160.250 ;
        RECT 120.840 160.170 123.030 160.250 ;
        RECT 125.840 160.170 128.030 160.400 ;
        RECT 136.840 160.170 139.030 160.400 ;
        RECT 141.250 160.250 144.030 160.400 ;
        RECT 141.840 160.170 144.030 160.250 ;
        RECT 78.500 159.500 144.750 160.000 ;
        RECT 112.500 158.750 121.250 159.250 ;
        RECT 127.750 158.750 136.000 159.250 ;
        RECT 91.750 158.000 120.500 158.500 ;
        RECT 92.500 157.250 124.250 157.750 ;
        RECT 130.750 157.250 142.500 158.500 ;
        RECT 145.000 157.000 146.000 163.500 ;
        RECT 22.250 155.500 23.250 156.500 ;
        RECT 11.000 154.500 23.250 155.500 ;
        RECT 11.000 150.500 11.500 154.500 ;
        RECT 11.685 152.175 11.915 154.500 ;
        RECT 12.125 152.000 12.355 154.175 ;
        RECT 12.565 152.175 12.795 154.500 ;
        RECT 13.005 152.000 13.235 154.175 ;
        RECT 13.445 152.175 13.675 154.500 ;
        RECT 13.885 152.000 14.115 154.175 ;
        RECT 14.325 152.175 14.555 154.500 ;
        RECT 14.765 152.000 14.995 154.175 ;
        RECT 15.205 152.175 15.435 154.500 ;
        RECT 15.645 152.000 15.875 154.175 ;
        RECT 16.085 152.175 16.315 154.500 ;
        RECT 12.125 151.500 15.875 152.000 ;
        RECT 13.750 150.750 14.250 151.250 ;
        RECT 16.500 150.500 17.000 154.500 ;
        RECT 17.185 152.175 17.415 154.500 ;
        RECT 17.625 152.000 17.855 154.175 ;
        RECT 18.065 152.175 18.295 154.500 ;
        RECT 18.505 152.000 18.735 154.175 ;
        RECT 18.945 152.175 19.175 154.500 ;
        RECT 19.385 152.000 19.615 154.175 ;
        RECT 19.825 152.175 20.055 154.500 ;
        RECT 20.265 152.000 20.495 154.175 ;
        RECT 20.705 152.175 20.935 154.500 ;
        RECT 21.145 152.000 21.375 154.175 ;
        RECT 21.585 152.175 21.815 154.500 ;
        RECT 17.625 151.500 21.375 152.000 ;
        RECT 19.250 150.750 19.750 151.250 ;
        RECT 22.000 150.500 22.500 154.500 ;
        RECT 11.000 150.000 22.500 150.500 ;
        RECT 22.750 150.500 23.250 154.500 ;
        RECT 23.585 152.250 23.815 156.500 ;
        RECT 24.045 152.000 24.275 156.250 ;
        RECT 24.505 152.250 24.735 156.500 ;
        RECT 24.965 152.000 25.195 156.250 ;
        RECT 25.425 152.250 25.655 156.500 ;
        RECT 25.885 152.000 26.115 156.250 ;
        RECT 26.345 152.250 26.575 156.500 ;
        RECT 26.805 152.000 27.035 156.250 ;
        RECT 27.265 152.250 27.495 156.500 ;
        RECT 27.725 152.000 27.955 156.250 ;
        RECT 28.185 152.250 28.415 156.500 ;
        RECT 24.045 151.500 27.955 152.000 ;
        RECT 25.750 150.750 26.250 151.250 ;
        RECT 28.750 150.500 29.250 156.500 ;
        RECT 29.585 152.250 29.815 156.500 ;
        RECT 30.045 152.000 30.275 156.250 ;
        RECT 30.505 152.250 30.735 156.500 ;
        RECT 30.965 152.000 31.195 156.250 ;
        RECT 31.425 152.250 31.655 156.500 ;
        RECT 31.885 152.000 32.115 156.250 ;
        RECT 32.345 152.250 32.575 156.500 ;
        RECT 32.805 152.000 33.035 156.250 ;
        RECT 33.265 152.250 33.495 156.500 ;
        RECT 33.725 152.000 33.955 156.250 ;
        RECT 34.185 152.250 34.415 156.500 ;
        RECT 30.045 151.500 33.955 152.000 ;
        RECT 31.750 150.750 32.250 151.250 ;
        RECT 34.750 150.500 35.250 156.500 ;
        RECT 35.585 152.250 35.815 156.500 ;
        RECT 36.045 152.000 36.275 156.250 ;
        RECT 36.505 152.250 36.735 156.500 ;
        RECT 36.965 152.000 37.195 156.250 ;
        RECT 37.425 152.250 37.655 156.500 ;
        RECT 37.885 152.000 38.115 156.250 ;
        RECT 38.345 152.250 38.575 156.500 ;
        RECT 38.805 152.000 39.035 156.250 ;
        RECT 39.265 152.250 39.495 156.500 ;
        RECT 39.725 152.000 39.955 156.250 ;
        RECT 40.185 152.250 40.415 156.500 ;
        RECT 40.750 155.500 42.250 156.500 ;
        RECT 45.250 155.500 45.750 156.500 ;
        RECT 48.750 155.500 49.250 156.500 ;
        RECT 52.250 155.500 52.750 156.500 ;
        RECT 40.750 155.000 52.750 155.500 ;
        RECT 77.250 155.000 146.500 157.000 ;
        RECT 36.045 151.500 39.955 152.000 ;
        RECT 37.750 150.750 38.250 151.250 ;
        RECT 40.750 150.500 42.250 155.000 ;
        RECT 43.250 154.250 44.250 154.750 ;
        RECT 22.750 150.000 42.250 150.500 ;
        RECT 11.000 149.000 22.500 149.500 ;
        RECT 11.000 145.000 11.500 149.000 ;
        RECT 13.750 148.250 14.250 148.750 ;
        RECT 12.125 147.500 15.875 148.000 ;
        RECT 11.685 145.000 11.915 147.250 ;
        RECT 12.125 145.250 12.355 147.500 ;
        RECT 12.565 145.000 12.795 147.250 ;
        RECT 13.005 145.250 13.235 147.500 ;
        RECT 13.445 145.000 13.675 147.250 ;
        RECT 13.885 145.250 14.115 147.500 ;
        RECT 14.325 145.000 14.555 147.250 ;
        RECT 14.765 145.250 14.995 147.500 ;
        RECT 15.205 145.000 15.435 147.250 ;
        RECT 15.645 145.250 15.875 147.500 ;
        RECT 16.085 145.000 16.315 147.250 ;
        RECT 16.500 145.000 17.000 149.000 ;
        RECT 19.250 148.250 19.750 148.750 ;
        RECT 17.625 147.500 21.375 148.000 ;
        RECT 17.185 145.000 17.415 147.250 ;
        RECT 17.625 145.250 17.855 147.500 ;
        RECT 18.065 145.000 18.295 147.250 ;
        RECT 18.505 145.250 18.735 147.500 ;
        RECT 18.945 145.000 19.175 147.250 ;
        RECT 19.385 145.250 19.615 147.500 ;
        RECT 19.825 145.000 20.055 147.250 ;
        RECT 20.265 145.250 20.495 147.500 ;
        RECT 20.705 145.000 20.935 147.250 ;
        RECT 21.145 145.250 21.375 147.500 ;
        RECT 21.585 145.000 21.815 147.250 ;
        RECT 22.000 145.000 22.500 149.000 ;
        RECT 22.750 149.000 41.250 149.500 ;
        RECT 22.750 145.000 23.250 149.000 ;
        RECT 25.750 148.250 26.250 148.750 ;
        RECT 24.045 147.500 27.955 148.000 ;
        RECT 11.000 144.000 23.250 145.000 ;
        RECT 22.250 143.000 23.250 144.000 ;
        RECT 23.585 143.000 23.815 147.250 ;
        RECT 24.045 143.250 24.275 147.500 ;
        RECT 24.505 143.000 24.735 147.250 ;
        RECT 24.965 143.250 25.195 147.500 ;
        RECT 25.425 143.000 25.655 147.250 ;
        RECT 25.885 143.250 26.115 147.500 ;
        RECT 26.345 143.000 26.575 147.250 ;
        RECT 26.805 143.250 27.035 147.500 ;
        RECT 27.265 143.000 27.495 147.250 ;
        RECT 27.725 143.250 27.955 147.500 ;
        RECT 28.185 143.000 28.415 147.250 ;
        RECT 28.750 143.000 29.250 149.000 ;
        RECT 31.750 148.250 32.250 148.750 ;
        RECT 30.045 147.500 33.955 148.000 ;
        RECT 29.585 143.000 29.815 147.250 ;
        RECT 30.045 143.250 30.275 147.500 ;
        RECT 30.505 143.000 30.735 147.250 ;
        RECT 30.965 143.250 31.195 147.500 ;
        RECT 31.425 143.000 31.655 147.250 ;
        RECT 31.885 143.250 32.115 147.500 ;
        RECT 32.345 143.000 32.575 147.250 ;
        RECT 32.805 143.250 33.035 147.500 ;
        RECT 33.265 143.000 33.495 147.250 ;
        RECT 33.725 143.250 33.955 147.500 ;
        RECT 34.185 143.000 34.415 147.250 ;
        RECT 34.750 143.000 35.250 149.000 ;
        RECT 37.750 148.250 38.250 148.750 ;
        RECT 36.045 147.500 39.955 148.000 ;
        RECT 35.585 143.000 35.815 147.250 ;
        RECT 36.045 143.250 36.275 147.500 ;
        RECT 36.505 143.000 36.735 147.250 ;
        RECT 36.965 143.250 37.195 147.500 ;
        RECT 37.425 143.000 37.655 147.250 ;
        RECT 37.885 143.250 38.115 147.500 ;
        RECT 38.345 143.000 38.575 147.250 ;
        RECT 38.805 143.250 39.035 147.500 ;
        RECT 39.265 143.000 39.495 147.250 ;
        RECT 39.725 143.250 39.955 147.500 ;
        RECT 40.185 143.000 40.415 147.250 ;
        RECT 40.750 143.000 41.250 149.000 ;
        RECT 41.750 144.500 42.250 150.000 ;
        RECT 42.500 145.500 43.220 154.000 ;
        RECT 44.280 145.500 45.000 154.000 ;
        RECT 43.250 144.750 44.250 145.250 ;
        RECT 45.250 144.500 45.750 155.000 ;
        RECT 46.750 154.250 47.750 154.750 ;
        RECT 46.000 145.500 46.720 154.000 ;
        RECT 47.780 145.500 48.500 154.000 ;
        RECT 46.750 144.750 47.750 145.250 ;
        RECT 48.750 144.500 49.250 155.000 ;
        RECT 50.250 154.250 51.250 154.750 ;
        RECT 49.500 145.500 50.220 154.000 ;
        RECT 51.280 145.500 52.000 154.000 ;
        RECT 50.250 144.750 51.250 145.250 ;
        RECT 52.250 144.500 52.750 155.000 ;
        RECT 77.250 152.500 146.500 154.500 ;
        RECT 54.000 150.000 132.750 152.000 ;
        RECT 111.500 148.880 140.500 149.360 ;
        RECT 111.500 146.160 142.000 146.640 ;
        RECT 130.740 145.960 131.060 146.020 ;
        RECT 135.370 145.960 135.690 146.020 ;
        RECT 130.740 145.820 135.690 145.960 ;
        RECT 130.740 145.760 131.060 145.820 ;
        RECT 135.370 145.760 135.690 145.820 ;
        RECT 137.210 145.760 137.530 146.020 ;
        RECT 117.890 145.420 118.210 145.680 ;
        RECT 132.150 145.420 132.470 145.680 ;
        RECT 117.430 144.940 117.750 145.000 ;
        RECT 118.825 144.940 119.115 144.985 ;
        RECT 117.430 144.800 119.115 144.940 ;
        RECT 117.430 144.740 117.750 144.800 ;
        RECT 118.825 144.755 119.115 144.800 ;
        RECT 120.205 144.940 120.495 144.985 ;
        RECT 121.110 144.940 121.430 145.000 ;
        RECT 130.785 144.940 131.075 144.985 ;
        RECT 120.205 144.800 131.075 144.940 ;
        RECT 120.205 144.755 120.495 144.800 ;
        RECT 121.110 144.740 121.430 144.800 ;
        RECT 130.785 144.755 131.075 144.800 ;
        RECT 41.750 144.000 52.750 144.500 ;
        RECT 130.860 144.600 131.000 144.755 ;
        RECT 131.230 144.740 131.550 145.000 ;
        RECT 134.450 144.740 134.770 145.000 ;
        RECT 133.085 144.600 133.375 144.645 ;
        RECT 134.910 144.600 135.230 144.660 ;
        RECT 130.860 144.460 135.230 144.600 ;
        RECT 133.085 144.415 133.375 144.460 ;
        RECT 134.910 144.400 135.230 144.460 ;
        RECT 119.745 144.260 120.035 144.305 ;
        RECT 120.190 144.260 120.510 144.320 ;
        RECT 119.745 144.120 120.510 144.260 ;
        RECT 119.745 144.075 120.035 144.120 ;
        RECT 120.190 144.060 120.510 144.120 ;
        RECT 133.530 144.060 133.850 144.320 ;
        RECT 111.500 143.440 140.500 143.920 ;
        RECT 120.665 143.240 120.955 143.285 ;
        RECT 133.530 143.240 133.850 143.300 ;
        RECT 120.665 143.100 133.850 143.240 ;
        RECT 120.665 143.055 120.955 143.100 ;
        RECT 20.750 142.000 53.000 143.000 ;
        RECT 120.190 142.900 120.510 142.960 ;
        RECT 129.020 142.945 129.160 143.100 ;
        RECT 133.530 143.040 133.850 143.100 ;
        RECT 121.125 142.900 121.415 142.945 ;
        RECT 119.360 142.760 121.415 142.900 ;
        RECT 119.360 142.220 119.500 142.760 ;
        RECT 120.190 142.700 120.510 142.760 ;
        RECT 121.125 142.715 121.415 142.760 ;
        RECT 128.945 142.715 129.235 142.945 ;
        RECT 129.865 142.900 130.155 142.945 ;
        RECT 132.150 142.900 132.470 142.960 ;
        RECT 129.865 142.760 132.470 142.900 ;
        RECT 129.865 142.715 130.155 142.760 ;
        RECT 119.745 142.560 120.035 142.605 ;
        RECT 129.940 142.560 130.080 142.715 ;
        RECT 132.150 142.700 132.470 142.760 ;
        RECT 133.070 142.700 133.390 142.960 ;
        RECT 119.745 142.420 130.080 142.560 ;
        RECT 119.745 142.375 120.035 142.420 ;
        RECT 131.230 142.360 131.550 142.620 ;
        RECT 130.265 142.220 130.585 142.280 ;
        RECT 134.005 142.220 134.295 142.265 ;
        RECT 134.450 142.220 134.770 142.280 ;
        RECT 119.360 142.080 130.080 142.220 ;
        RECT 21.000 141.250 25.500 141.750 ;
        RECT 21.000 138.000 22.000 141.250 ;
        RECT 23.000 140.500 23.500 141.000 ;
        RECT 22.250 139.250 22.790 140.250 ;
        RECT 23.000 139.250 23.500 140.250 ;
        RECT 23.710 139.250 24.250 140.250 ;
        RECT 22.250 138.750 22.750 139.250 ;
        RECT 23.000 138.500 23.500 139.000 ;
        RECT 23.750 138.750 24.250 139.250 ;
        RECT 24.500 138.000 25.500 141.250 ;
        RECT 21.000 137.500 25.500 138.000 ;
        RECT 21.000 134.250 22.000 137.500 ;
        RECT 23.000 136.750 23.500 137.250 ;
        RECT 22.250 135.500 22.790 136.500 ;
        RECT 23.000 135.500 23.500 136.500 ;
        RECT 23.710 135.500 24.250 136.500 ;
        RECT 22.250 135.000 22.750 135.500 ;
        RECT 23.000 134.750 23.500 135.250 ;
        RECT 23.750 135.000 24.250 135.500 ;
        RECT 24.500 134.250 25.500 137.500 ;
        RECT 21.000 133.750 25.500 134.250 ;
        RECT 21.000 130.500 22.000 133.750 ;
        RECT 23.000 133.000 23.500 133.500 ;
        RECT 22.250 131.750 22.790 132.750 ;
        RECT 23.000 131.750 23.500 132.750 ;
        RECT 23.710 131.750 24.250 132.750 ;
        RECT 22.250 131.250 22.750 131.750 ;
        RECT 23.000 131.000 23.500 131.500 ;
        RECT 23.750 131.250 24.250 131.750 ;
        RECT 24.500 130.500 25.500 133.750 ;
        RECT 21.000 130.000 25.500 130.500 ;
        RECT 21.000 126.750 22.000 130.000 ;
        RECT 23.000 129.250 23.500 129.750 ;
        RECT 22.250 128.000 22.790 129.000 ;
        RECT 23.000 128.000 23.500 129.000 ;
        RECT 23.710 128.000 24.250 129.000 ;
        RECT 22.250 127.500 22.750 128.000 ;
        RECT 23.000 127.250 23.500 127.750 ;
        RECT 23.750 127.500 24.250 128.000 ;
        RECT 24.500 126.750 25.500 130.000 ;
        RECT 21.000 126.250 25.500 126.750 ;
        RECT 21.000 123.000 22.000 126.250 ;
        RECT 23.000 125.500 23.500 126.000 ;
        RECT 22.250 124.250 22.790 125.250 ;
        RECT 23.000 124.250 23.500 125.250 ;
        RECT 23.710 124.250 24.250 125.250 ;
        RECT 22.250 123.750 22.750 124.250 ;
        RECT 23.000 123.500 23.500 124.000 ;
        RECT 23.750 123.750 24.250 124.250 ;
        RECT 24.500 123.000 25.500 126.250 ;
        RECT 21.000 122.500 25.500 123.000 ;
        RECT 21.000 119.250 22.000 122.500 ;
        RECT 23.000 121.750 23.500 122.250 ;
        RECT 22.250 120.500 22.790 121.500 ;
        RECT 23.000 120.500 23.500 121.500 ;
        RECT 23.710 120.500 24.250 121.500 ;
        RECT 22.250 120.000 22.750 120.500 ;
        RECT 23.000 119.750 23.500 120.250 ;
        RECT 23.750 120.000 24.250 120.500 ;
        RECT 24.500 119.250 25.500 122.500 ;
        RECT 21.000 118.750 25.500 119.250 ;
        RECT 21.000 115.500 22.000 118.750 ;
        RECT 23.000 118.000 23.500 118.500 ;
        RECT 22.250 116.750 22.790 117.750 ;
        RECT 23.000 116.750 23.500 117.750 ;
        RECT 23.710 116.750 24.250 117.750 ;
        RECT 22.250 116.250 22.750 116.750 ;
        RECT 23.000 116.000 23.500 116.500 ;
        RECT 23.750 116.250 24.250 116.750 ;
        RECT 24.500 115.500 25.500 118.750 ;
        RECT 21.000 115.000 25.500 115.500 ;
        RECT 21.000 111.750 22.000 115.000 ;
        RECT 23.000 114.250 23.500 114.750 ;
        RECT 22.250 113.000 22.790 114.000 ;
        RECT 23.000 113.000 23.500 114.000 ;
        RECT 23.710 113.000 24.250 114.000 ;
        RECT 22.250 112.500 22.750 113.000 ;
        RECT 23.000 112.250 23.500 112.750 ;
        RECT 23.750 112.500 24.250 113.000 ;
        RECT 24.500 111.750 25.500 115.000 ;
        RECT 21.000 111.000 25.500 111.750 ;
        RECT 30.500 141.250 35.000 141.750 ;
        RECT 30.500 138.000 31.500 141.250 ;
        RECT 32.500 140.500 33.000 141.000 ;
        RECT 31.750 139.250 32.290 140.250 ;
        RECT 32.500 139.250 33.000 140.250 ;
        RECT 33.210 139.250 33.750 140.250 ;
        RECT 31.750 138.750 32.250 139.250 ;
        RECT 32.500 138.500 33.000 139.000 ;
        RECT 33.250 138.750 33.750 139.250 ;
        RECT 34.000 138.000 35.000 141.250 ;
        RECT 30.500 137.500 35.000 138.000 ;
        RECT 30.500 134.250 31.500 137.500 ;
        RECT 32.500 136.750 33.000 137.250 ;
        RECT 31.750 135.500 32.290 136.500 ;
        RECT 32.500 135.500 33.000 136.500 ;
        RECT 33.210 135.500 33.750 136.500 ;
        RECT 31.750 135.000 32.250 135.500 ;
        RECT 32.500 134.750 33.000 135.250 ;
        RECT 33.250 135.000 33.750 135.500 ;
        RECT 34.000 134.250 35.000 137.500 ;
        RECT 30.500 133.750 35.000 134.250 ;
        RECT 30.500 130.500 31.500 133.750 ;
        RECT 32.500 133.000 33.000 133.500 ;
        RECT 31.750 131.750 32.290 132.750 ;
        RECT 32.500 131.750 33.000 132.750 ;
        RECT 33.210 131.750 33.750 132.750 ;
        RECT 31.750 131.250 32.250 131.750 ;
        RECT 32.500 131.000 33.000 131.500 ;
        RECT 33.250 131.250 33.750 131.750 ;
        RECT 34.000 130.500 35.000 133.750 ;
        RECT 30.500 130.000 35.000 130.500 ;
        RECT 30.500 126.750 31.500 130.000 ;
        RECT 32.500 129.250 33.000 129.750 ;
        RECT 31.750 128.000 32.290 129.000 ;
        RECT 32.500 128.000 33.000 129.000 ;
        RECT 33.210 128.000 33.750 129.000 ;
        RECT 31.750 127.500 32.250 128.000 ;
        RECT 32.500 127.250 33.000 127.750 ;
        RECT 33.250 127.500 33.750 128.000 ;
        RECT 34.000 126.750 35.000 130.000 ;
        RECT 30.500 126.250 35.000 126.750 ;
        RECT 30.500 123.000 31.500 126.250 ;
        RECT 32.500 125.500 33.000 126.000 ;
        RECT 31.750 124.250 32.290 125.250 ;
        RECT 32.500 124.250 33.000 125.250 ;
        RECT 33.210 124.250 33.750 125.250 ;
        RECT 31.750 123.750 32.250 124.250 ;
        RECT 32.500 123.500 33.000 124.000 ;
        RECT 33.250 123.750 33.750 124.250 ;
        RECT 34.000 123.000 35.000 126.250 ;
        RECT 30.500 122.500 35.000 123.000 ;
        RECT 30.500 119.250 31.500 122.500 ;
        RECT 32.500 121.750 33.000 122.250 ;
        RECT 31.750 120.500 32.290 121.500 ;
        RECT 32.500 120.500 33.000 121.500 ;
        RECT 33.210 120.500 33.750 121.500 ;
        RECT 31.750 120.000 32.250 120.500 ;
        RECT 32.500 119.750 33.000 120.250 ;
        RECT 33.250 120.000 33.750 120.500 ;
        RECT 34.000 119.250 35.000 122.500 ;
        RECT 30.500 118.750 35.000 119.250 ;
        RECT 30.500 115.500 31.500 118.750 ;
        RECT 32.500 118.000 33.000 118.500 ;
        RECT 31.750 116.750 32.290 117.750 ;
        RECT 32.500 116.750 33.000 117.750 ;
        RECT 33.210 116.750 33.750 117.750 ;
        RECT 31.750 116.250 32.250 116.750 ;
        RECT 32.500 116.000 33.000 116.500 ;
        RECT 33.250 116.250 33.750 116.750 ;
        RECT 34.000 115.500 35.000 118.750 ;
        RECT 30.500 115.000 35.000 115.500 ;
        RECT 30.500 111.750 31.500 115.000 ;
        RECT 32.500 114.250 33.000 114.750 ;
        RECT 31.750 113.000 32.290 114.000 ;
        RECT 32.500 113.000 33.000 114.000 ;
        RECT 33.210 113.000 33.750 114.000 ;
        RECT 31.750 112.500 32.250 113.000 ;
        RECT 32.500 112.250 33.000 112.750 ;
        RECT 33.250 112.500 33.750 113.000 ;
        RECT 34.000 111.750 35.000 115.000 ;
        RECT 30.500 111.000 35.000 111.750 ;
        RECT 40.000 141.250 44.500 141.750 ;
        RECT 50.250 141.250 71.500 141.750 ;
        RECT 117.430 141.540 117.750 141.600 ;
        RECT 129.940 141.585 130.080 142.080 ;
        RECT 130.265 142.080 134.770 142.220 ;
        RECT 130.265 142.020 130.585 142.080 ;
        RECT 134.005 142.035 134.295 142.080 ;
        RECT 134.450 142.020 134.770 142.080 ;
        RECT 118.825 141.540 119.115 141.585 ;
        RECT 117.430 141.400 119.115 141.540 ;
        RECT 117.430 141.340 117.750 141.400 ;
        RECT 118.825 141.355 119.115 141.400 ;
        RECT 129.865 141.540 130.155 141.585 ;
        RECT 133.070 141.540 133.390 141.600 ;
        RECT 129.865 141.400 133.390 141.540 ;
        RECT 129.865 141.355 130.155 141.400 ;
        RECT 133.070 141.340 133.390 141.400 ;
        RECT 40.000 138.000 41.000 141.250 ;
        RECT 42.000 140.500 42.500 141.000 ;
        RECT 41.250 139.250 41.790 140.250 ;
        RECT 42.000 139.250 42.500 140.250 ;
        RECT 42.710 139.250 43.250 140.250 ;
        RECT 41.250 138.750 41.750 139.250 ;
        RECT 42.000 138.500 42.500 139.000 ;
        RECT 42.750 138.750 43.250 139.250 ;
        RECT 43.500 138.000 44.500 141.250 ;
        RECT 111.500 140.720 142.000 141.200 ;
        RECT 118.350 139.980 118.670 140.240 ;
        RECT 119.285 139.500 119.575 139.545 ;
        RECT 120.650 139.500 120.970 139.560 ;
        RECT 119.285 139.360 120.970 139.500 ;
        RECT 119.285 139.315 119.575 139.360 ;
        RECT 120.650 139.300 120.970 139.360 ;
        RECT 111.500 138.000 140.500 138.480 ;
        RECT 40.000 137.500 44.500 138.000 ;
        RECT 50.250 137.500 69.500 138.000 ;
        RECT 134.465 137.800 134.755 137.845 ;
        RECT 136.290 137.800 136.610 137.860 ;
        RECT 134.465 137.660 136.610 137.800 ;
        RECT 134.465 137.615 134.755 137.660 ;
        RECT 136.290 137.600 136.610 137.660 ;
        RECT 40.000 134.250 41.000 137.500 ;
        RECT 42.000 136.750 42.500 137.250 ;
        RECT 41.250 135.500 41.790 136.500 ;
        RECT 42.000 135.500 42.500 136.500 ;
        RECT 42.710 135.500 43.250 136.500 ;
        RECT 41.250 135.000 41.750 135.500 ;
        RECT 42.000 134.750 42.500 135.250 ;
        RECT 42.750 135.000 43.250 135.500 ;
        RECT 43.500 134.250 44.500 137.500 ;
        RECT 114.670 137.460 114.990 137.520 ;
        RECT 117.905 137.460 118.195 137.505 ;
        RECT 114.670 137.320 118.195 137.460 ;
        RECT 114.670 137.260 114.990 137.320 ;
        RECT 117.905 137.275 118.195 137.320 ;
        RECT 120.205 137.460 120.495 137.505 ;
        RECT 121.110 137.460 121.430 137.520 ;
        RECT 133.530 137.460 133.850 137.520 ;
        RECT 135.370 137.460 135.690 137.520 ;
        RECT 120.205 137.320 121.430 137.460 ;
        RECT 120.205 137.275 120.495 137.320 ;
        RECT 121.110 137.260 121.430 137.320 ;
        RECT 132.240 137.320 135.690 137.460 ;
        RECT 118.810 136.920 119.130 137.180 ;
        RECT 119.745 137.120 120.035 137.165 ;
        RECT 120.650 137.120 120.970 137.180 ;
        RECT 132.240 137.165 132.380 137.320 ;
        RECT 133.530 137.260 133.850 137.320 ;
        RECT 135.370 137.260 135.690 137.320 ;
        RECT 119.745 136.980 120.970 137.120 ;
        RECT 119.745 136.935 120.035 136.980 ;
        RECT 120.650 136.920 120.970 136.980 ;
        RECT 132.165 136.935 132.455 137.165 ;
        RECT 133.530 136.780 133.850 136.840 ;
        RECT 133.990 136.780 134.310 136.840 ;
        RECT 133.530 136.640 134.310 136.780 ;
        RECT 133.530 136.580 133.850 136.640 ;
        RECT 133.990 136.580 134.310 136.640 ;
        RECT 132.625 136.440 132.915 136.485 ;
        RECT 134.910 136.440 135.230 136.500 ;
        RECT 132.625 136.300 135.230 136.440 ;
        RECT 132.625 136.255 132.915 136.300 ;
        RECT 134.910 136.240 135.230 136.300 ;
        RECT 111.500 135.280 142.000 135.760 ;
        RECT 133.990 134.880 134.310 135.140 ;
        RECT 134.925 134.895 135.215 135.125 ;
        RECT 131.690 134.740 132.010 134.800 ;
        RECT 133.070 134.740 133.390 134.800 ;
        RECT 135.000 134.740 135.140 134.895 ;
        RECT 131.690 134.600 135.140 134.740 ;
        RECT 131.690 134.540 132.010 134.600 ;
        RECT 133.070 134.540 133.390 134.600 ;
        RECT 40.000 133.750 44.500 134.250 ;
        RECT 50.250 133.750 67.500 134.250 ;
        RECT 135.370 134.200 135.690 134.460 ;
        RECT 132.150 134.060 132.470 134.120 ;
        RECT 134.450 134.060 134.770 134.120 ;
        RECT 135.845 134.060 136.135 134.105 ;
        RECT 132.150 133.920 136.135 134.060 ;
        RECT 132.150 133.860 132.470 133.920 ;
        RECT 134.450 133.860 134.770 133.920 ;
        RECT 135.845 133.875 136.135 133.920 ;
        RECT 40.000 130.500 41.000 133.750 ;
        RECT 42.000 133.000 42.500 133.500 ;
        RECT 41.250 131.750 41.790 132.750 ;
        RECT 42.000 131.750 42.500 132.750 ;
        RECT 42.710 131.750 43.250 132.750 ;
        RECT 41.250 131.250 41.750 131.750 ;
        RECT 42.000 131.000 42.500 131.500 ;
        RECT 42.750 131.250 43.250 131.750 ;
        RECT 43.500 130.500 44.500 133.750 ;
        RECT 134.770 133.240 135.730 133.380 ;
        RECT 111.500 132.560 140.500 133.040 ;
        RECT 118.350 132.360 118.670 132.420 ;
        RECT 118.810 132.360 119.130 132.420 ;
        RECT 134.005 132.360 134.295 132.405 ;
        RECT 118.350 132.220 119.130 132.360 ;
        RECT 118.350 132.160 118.670 132.220 ;
        RECT 118.810 132.160 119.130 132.220 ;
        RECT 120.740 132.220 134.295 132.360 ;
        RECT 119.270 132.020 119.590 132.080 ;
        RECT 120.740 132.020 120.880 132.220 ;
        RECT 134.005 132.175 134.295 132.220 ;
        RECT 119.270 131.880 120.880 132.020 ;
        RECT 119.270 131.820 119.590 131.880 ;
        RECT 120.740 131.725 120.880 131.880 ;
        RECT 133.085 132.020 133.375 132.065 ;
        RECT 133.530 132.020 133.850 132.080 ;
        RECT 133.085 131.880 133.850 132.020 ;
        RECT 134.080 132.020 134.220 132.175 ;
        RECT 134.450 132.160 134.770 132.420 ;
        RECT 134.080 131.880 134.680 132.020 ;
        RECT 133.085 131.835 133.375 131.880 ;
        RECT 133.530 131.820 133.850 131.880 ;
        RECT 120.665 131.495 120.955 131.725 ;
        RECT 131.705 131.495 131.995 131.725 ;
        RECT 132.625 131.680 132.915 131.725 ;
        RECT 133.990 131.680 134.310 131.740 ;
        RECT 132.625 131.540 134.310 131.680 ;
        RECT 134.540 131.680 134.680 131.880 ;
        RECT 134.910 131.820 135.230 132.080 ;
        RECT 135.830 131.820 136.150 132.080 ;
        RECT 135.370 131.680 135.690 131.740 ;
        RECT 134.540 131.540 135.690 131.680 ;
        RECT 132.625 131.495 132.915 131.540 ;
        RECT 119.285 131.340 119.575 131.385 ;
        RECT 131.780 131.340 131.920 131.495 ;
        RECT 133.990 131.480 134.310 131.540 ;
        RECT 135.370 131.480 135.690 131.540 ;
        RECT 134.910 131.340 135.230 131.400 ;
        RECT 119.285 131.200 120.880 131.340 ;
        RECT 131.780 131.200 135.230 131.340 ;
        RECT 119.285 131.155 119.575 131.200 ;
        RECT 120.740 131.060 120.880 131.200 ;
        RECT 134.910 131.140 135.230 131.200 ;
        RECT 120.205 130.815 120.495 131.045 ;
        RECT 118.810 130.660 119.130 130.720 ;
        RECT 120.280 130.660 120.420 130.815 ;
        RECT 120.650 130.800 120.970 131.060 ;
        RECT 131.690 131.000 132.010 131.060 ;
        RECT 121.200 130.860 132.010 131.000 ;
        RECT 121.200 130.660 121.340 130.860 ;
        RECT 131.690 130.800 132.010 130.860 ;
        RECT 118.810 130.520 121.340 130.660 ;
        RECT 40.000 130.000 44.500 130.500 ;
        RECT 50.250 130.000 65.500 130.500 ;
        RECT 118.810 130.460 119.130 130.520 ;
        RECT 131.215 130.460 131.535 130.720 ;
        RECT 40.000 126.750 41.000 130.000 ;
        RECT 42.000 129.250 42.500 129.750 ;
        RECT 41.250 128.000 41.790 129.000 ;
        RECT 42.000 128.000 42.500 129.000 ;
        RECT 42.710 128.000 43.250 129.000 ;
        RECT 41.250 127.500 41.750 128.000 ;
        RECT 42.000 127.250 42.500 127.750 ;
        RECT 42.750 127.500 43.250 128.000 ;
        RECT 43.500 126.750 44.500 130.000 ;
        RECT 111.500 129.840 142.000 130.320 ;
        RECT 133.530 129.440 133.850 129.700 ;
        RECT 116.970 129.300 117.290 129.360 ;
        RECT 117.430 129.300 117.750 129.360 ;
        RECT 116.970 129.160 117.750 129.300 ;
        RECT 116.970 129.100 117.290 129.160 ;
        RECT 117.430 129.100 117.750 129.160 ;
        RECT 131.690 128.760 132.010 129.020 ;
        RECT 120.205 128.620 120.495 128.665 ;
        RECT 120.650 128.620 120.970 128.680 ;
        RECT 132.610 128.620 132.930 128.680 ;
        RECT 134.450 128.620 134.770 128.680 ;
        RECT 120.205 128.480 134.770 128.620 ;
        RECT 120.205 128.435 120.495 128.480 ;
        RECT 120.650 128.420 120.970 128.480 ;
        RECT 132.610 128.420 132.930 128.480 ;
        RECT 134.450 128.420 134.770 128.480 ;
        RECT 118.365 128.280 118.655 128.325 ;
        RECT 121.110 128.280 121.430 128.340 ;
        RECT 118.365 128.140 121.430 128.280 ;
        RECT 118.365 128.095 118.655 128.140 ;
        RECT 121.110 128.080 121.430 128.140 ;
        RECT 118.810 127.740 119.130 128.000 ;
        RECT 119.270 127.740 119.590 128.000 ;
        RECT 111.500 127.120 140.500 127.600 ;
        RECT 40.000 126.250 44.500 126.750 ;
        RECT 50.250 126.250 63.500 126.750 ;
        RECT 40.000 123.000 41.000 126.250 ;
        RECT 42.000 125.500 42.500 126.000 ;
        RECT 41.250 124.250 41.790 125.250 ;
        RECT 42.000 124.250 42.500 125.250 ;
        RECT 42.710 124.250 43.250 125.250 ;
        RECT 41.250 123.750 41.750 124.250 ;
        RECT 42.000 123.500 42.500 124.000 ;
        RECT 42.750 123.750 43.250 124.250 ;
        RECT 43.500 123.000 44.500 126.250 ;
        RECT 85.250 123.250 110.750 124.500 ;
        RECT 111.500 124.400 142.000 124.880 ;
        RECT 40.000 122.500 44.500 123.000 ;
        RECT 50.250 122.500 61.500 123.000 ;
        RECT 40.000 119.250 41.000 122.500 ;
        RECT 42.000 121.750 42.500 122.250 ;
        RECT 41.250 120.500 41.790 121.500 ;
        RECT 42.000 120.500 42.500 121.500 ;
        RECT 42.710 120.500 43.250 121.500 ;
        RECT 41.250 120.000 41.750 120.500 ;
        RECT 42.000 119.750 42.500 120.250 ;
        RECT 42.750 120.000 43.250 120.500 ;
        RECT 43.500 119.250 44.500 122.500 ;
        RECT 88.250 119.250 88.750 123.250 ;
        RECT 89.025 122.500 91.015 123.250 ;
        RECT 89.025 120.890 89.255 122.500 ;
        RECT 89.465 120.750 89.695 121.890 ;
        RECT 89.905 120.890 90.135 122.500 ;
        RECT 90.345 120.750 90.575 121.890 ;
        RECT 90.785 120.890 91.015 122.500 ;
        RECT 91.435 122.500 93.425 123.250 ;
        RECT 91.435 120.890 91.665 122.500 ;
        RECT 91.875 120.750 92.105 121.890 ;
        RECT 92.315 120.890 92.545 122.500 ;
        RECT 92.755 120.750 92.985 121.890 ;
        RECT 93.195 120.890 93.425 122.500 ;
        RECT 93.845 122.500 95.835 123.250 ;
        RECT 93.845 120.890 94.075 122.500 ;
        RECT 94.285 120.750 94.515 121.890 ;
        RECT 94.725 120.890 94.955 122.500 ;
        RECT 95.165 120.750 95.395 121.890 ;
        RECT 95.605 120.890 95.835 122.500 ;
        RECT 96.255 122.500 98.245 123.250 ;
        RECT 96.255 120.890 96.485 122.500 ;
        RECT 96.695 120.750 96.925 121.890 ;
        RECT 97.135 120.890 97.365 122.500 ;
        RECT 97.575 120.750 97.805 121.890 ;
        RECT 98.015 120.890 98.245 122.500 ;
        RECT 98.665 122.500 100.660 123.000 ;
        RECT 101.075 122.500 103.065 123.250 ;
        RECT 103.480 122.500 105.475 123.000 ;
        RECT 98.665 120.890 98.895 122.500 ;
        RECT 99.105 120.750 99.335 121.890 ;
        RECT 99.545 120.890 99.775 122.500 ;
        RECT 99.985 120.750 100.215 121.890 ;
        RECT 100.425 120.890 100.655 122.500 ;
        RECT 101.075 120.890 101.305 122.500 ;
        RECT 101.515 120.750 101.745 121.890 ;
        RECT 101.955 120.890 102.185 122.500 ;
        RECT 102.395 120.750 102.625 121.890 ;
        RECT 102.835 120.890 103.065 122.500 ;
        RECT 103.485 120.890 103.715 122.500 ;
        RECT 89.465 120.250 91.020 120.750 ;
        RECT 91.875 120.250 93.430 120.750 ;
        RECT 93.840 120.250 95.395 120.750 ;
        RECT 96.250 120.250 98.250 120.750 ;
        RECT 98.660 120.250 100.215 120.750 ;
        RECT 101.070 120.250 102.625 120.750 ;
        RECT 103.925 120.750 104.155 121.890 ;
        RECT 104.365 120.890 104.595 122.500 ;
        RECT 104.805 120.750 105.035 121.890 ;
        RECT 105.245 120.890 105.475 122.500 ;
        RECT 103.925 120.250 105.480 120.750 ;
        RECT 89.770 119.500 92.680 120.000 ;
        RECT 92.930 119.500 95.090 120.000 ;
        RECT 97.000 119.500 97.500 120.000 ;
        RECT 99.410 119.500 101.570 120.000 ;
        RECT 101.820 119.500 104.730 120.000 ;
        RECT 105.750 119.250 106.250 123.250 ;
        RECT 40.000 118.750 44.500 119.250 ;
        RECT 50.250 118.750 59.500 119.250 ;
        RECT 85.250 118.750 110.750 119.250 ;
        RECT 40.000 115.500 41.000 118.750 ;
        RECT 42.000 118.000 42.500 118.500 ;
        RECT 41.250 116.750 41.790 117.750 ;
        RECT 42.000 116.750 42.500 117.750 ;
        RECT 42.710 116.750 43.250 117.750 ;
        RECT 41.250 116.250 41.750 116.750 ;
        RECT 42.000 116.000 42.500 116.500 ;
        RECT 42.750 116.250 43.250 116.750 ;
        RECT 43.500 115.500 44.500 118.750 ;
        RECT 76.250 118.250 82.750 118.750 ;
        RECT 40.000 115.000 44.500 115.500 ;
        RECT 50.250 115.000 57.500 115.500 ;
        RECT 76.250 115.250 76.750 118.250 ;
        RECT 77.750 117.500 78.250 118.000 ;
        RECT 77.000 116.250 77.895 117.250 ;
        RECT 78.105 116.250 79.000 117.250 ;
        RECT 77.750 115.500 78.250 116.000 ;
        RECT 79.250 115.250 79.750 118.250 ;
        RECT 80.750 117.500 81.250 118.000 ;
        RECT 80.000 116.250 80.895 117.250 ;
        RECT 81.105 116.250 82.000 117.250 ;
        RECT 80.750 115.500 81.250 116.000 ;
        RECT 82.250 115.250 82.750 118.250 ;
        RECT 93.840 118.000 103.980 118.500 ;
        RECT 86.750 117.250 90.270 117.750 ;
        RECT 90.520 117.250 100.660 117.750 ;
        RECT 104.230 117.250 107.750 117.750 ;
        RECT 95.340 116.500 105.480 117.000 ;
        RECT 86.750 115.750 90.270 116.250 ;
        RECT 90.520 115.750 103.980 116.250 ;
        RECT 104.230 115.750 107.750 116.250 ;
        RECT 40.000 111.750 41.000 115.000 ;
        RECT 42.000 114.250 42.500 114.750 ;
        RECT 41.250 113.000 41.790 114.000 ;
        RECT 42.000 113.000 42.500 114.000 ;
        RECT 42.710 113.000 43.250 114.000 ;
        RECT 41.250 112.500 41.750 113.000 ;
        RECT 42.000 112.250 42.500 112.750 ;
        RECT 42.750 112.500 43.250 113.000 ;
        RECT 43.500 111.750 44.500 115.000 ;
        RECT 76.250 114.000 82.750 115.250 ;
        RECT 83.750 115.000 109.250 115.500 ;
        RECT 40.000 111.000 44.500 111.750 ;
        RECT 20.750 110.000 49.250 111.000 ;
        RECT 88.250 110.250 88.750 115.000 ;
        RECT 89.770 114.250 92.680 114.750 ;
        RECT 92.930 114.250 95.090 114.750 ;
        RECT 97.000 114.250 97.500 114.750 ;
        RECT 99.410 114.250 101.570 114.750 ;
        RECT 101.820 114.250 104.730 114.750 ;
        RECT 89.465 113.500 91.020 114.000 ;
        RECT 91.875 113.500 93.430 114.000 ;
        RECT 94.285 113.500 95.840 114.000 ;
        RECT 96.250 113.500 98.250 114.000 ;
        RECT 99.105 113.500 100.660 114.000 ;
        RECT 101.070 113.500 102.625 114.000 ;
        RECT 89.025 111.000 89.255 113.360 ;
        RECT 89.465 111.360 89.695 113.500 ;
        RECT 89.905 111.000 90.135 113.360 ;
        RECT 90.345 111.360 90.575 113.500 ;
        RECT 90.785 111.000 91.015 113.360 ;
        RECT 89.025 110.250 91.015 111.000 ;
        RECT 91.435 111.000 91.665 113.360 ;
        RECT 91.875 111.360 92.105 113.500 ;
        RECT 92.315 111.000 92.545 113.360 ;
        RECT 92.755 111.360 92.985 113.500 ;
        RECT 93.195 111.000 93.425 113.360 ;
        RECT 93.845 111.000 94.075 113.360 ;
        RECT 94.285 111.360 94.515 113.500 ;
        RECT 94.725 111.000 94.955 113.360 ;
        RECT 95.165 111.360 95.395 113.500 ;
        RECT 95.605 111.000 95.835 113.360 ;
        RECT 91.435 110.250 93.425 111.000 ;
        RECT 93.840 110.500 95.835 111.000 ;
        RECT 96.255 111.000 96.485 113.360 ;
        RECT 96.695 111.360 96.925 113.500 ;
        RECT 97.135 111.000 97.365 113.360 ;
        RECT 97.575 111.360 97.805 113.500 ;
        RECT 98.015 111.000 98.245 113.360 ;
        RECT 96.255 110.250 98.245 111.000 ;
        RECT 98.665 111.000 98.895 113.360 ;
        RECT 99.105 111.360 99.335 113.500 ;
        RECT 99.545 111.000 99.775 113.360 ;
        RECT 99.985 111.360 100.215 113.500 ;
        RECT 100.425 111.000 100.655 113.360 ;
        RECT 98.665 110.250 100.655 111.000 ;
        RECT 101.075 111.000 101.305 113.360 ;
        RECT 101.515 111.360 101.745 113.500 ;
        RECT 101.955 111.000 102.185 113.360 ;
        RECT 102.395 111.360 102.625 113.500 ;
        RECT 103.925 113.500 105.480 114.000 ;
        RECT 102.835 111.000 103.065 113.360 ;
        RECT 103.485 111.000 103.715 113.360 ;
        RECT 103.925 111.360 104.155 113.500 ;
        RECT 104.365 111.000 104.595 113.360 ;
        RECT 104.805 111.360 105.035 113.500 ;
        RECT 105.245 111.000 105.475 113.360 ;
        RECT 101.075 110.250 103.065 111.000 ;
        RECT 103.480 110.500 105.475 111.000 ;
        RECT 105.750 110.250 106.250 115.000 ;
        RECT 83.750 109.000 109.250 110.250 ;
        RECT 0.000 104.000 147.500 108.000 ;
        RECT 5.000 99.000 147.500 103.000 ;
      LAYER met2 ;
        RECT 0.000 200.000 4.000 204.000 ;
        RECT 5.000 195.000 9.000 199.000 ;
        RECT 12.250 143.500 13.250 156.000 ;
        RECT 13.750 148.250 14.250 151.250 ;
        RECT 0.000 104.000 4.000 108.000 ;
        RECT 15.500 104.000 16.750 204.000 ;
        RECT 18.750 154.500 19.750 199.000 ;
        RECT 21.000 188.500 22.000 199.000 ;
        RECT 24.500 188.500 25.500 199.000 ;
        RECT 29.250 188.500 29.750 189.500 ;
        RECT 30.500 188.500 31.500 199.000 ;
        RECT 34.000 188.500 35.000 199.000 ;
        RECT 38.750 188.500 39.250 189.500 ;
        RECT 40.000 188.500 41.000 199.000 ;
        RECT 43.500 188.500 44.500 199.000 ;
        RECT 48.250 188.500 49.250 199.000 ;
        RECT 22.250 186.500 22.750 187.000 ;
        RECT 23.750 186.500 24.250 187.000 ;
        RECT 31.750 186.500 32.250 187.000 ;
        RECT 33.250 186.500 33.750 187.000 ;
        RECT 41.250 186.500 41.750 187.000 ;
        RECT 42.750 186.500 43.250 187.000 ;
        RECT 23.000 185.500 23.500 186.000 ;
        RECT 32.500 185.500 33.000 186.000 ;
        RECT 42.000 185.500 42.500 186.000 ;
        RECT 23.000 184.500 23.500 185.250 ;
        RECT 32.500 184.500 33.000 185.250 ;
        RECT 42.000 184.500 42.500 185.250 ;
        RECT 20.750 184.000 50.750 184.500 ;
        RECT 22.250 182.750 22.750 183.250 ;
        RECT 23.750 182.750 24.250 183.250 ;
        RECT 31.750 182.750 32.250 183.250 ;
        RECT 33.250 182.750 33.750 183.250 ;
        RECT 41.250 182.750 41.750 183.250 ;
        RECT 42.750 182.750 43.250 183.250 ;
        RECT 23.000 181.750 23.500 182.250 ;
        RECT 32.500 181.750 33.000 182.250 ;
        RECT 42.000 181.750 42.500 182.250 ;
        RECT 23.000 180.750 23.500 181.500 ;
        RECT 32.500 180.750 33.000 181.500 ;
        RECT 42.000 180.750 42.500 181.500 ;
        RECT 20.750 180.250 50.750 180.750 ;
        RECT 22.250 179.000 22.750 179.500 ;
        RECT 23.750 179.000 24.250 179.500 ;
        RECT 31.750 179.000 32.250 179.500 ;
        RECT 33.250 179.000 33.750 179.500 ;
        RECT 41.250 179.000 41.750 179.500 ;
        RECT 42.750 179.000 43.250 179.500 ;
        RECT 23.000 178.000 23.500 178.500 ;
        RECT 32.500 178.000 33.000 178.500 ;
        RECT 42.000 178.000 42.500 178.500 ;
        RECT 23.000 177.000 23.500 177.750 ;
        RECT 32.500 177.000 33.000 177.750 ;
        RECT 42.000 177.000 42.500 177.750 ;
        RECT 20.750 176.500 50.750 177.000 ;
        RECT 22.250 175.250 22.750 175.750 ;
        RECT 23.750 175.250 24.250 175.750 ;
        RECT 31.750 175.250 32.250 175.750 ;
        RECT 33.250 175.250 33.750 175.750 ;
        RECT 41.250 175.250 41.750 175.750 ;
        RECT 42.750 175.250 43.250 175.750 ;
        RECT 23.000 174.250 23.500 174.750 ;
        RECT 32.500 174.250 33.000 174.750 ;
        RECT 42.000 174.250 42.500 174.750 ;
        RECT 23.000 173.250 23.500 174.000 ;
        RECT 32.500 173.250 33.000 174.000 ;
        RECT 42.000 173.250 42.500 174.000 ;
        RECT 20.750 172.750 50.750 173.250 ;
        RECT 22.250 171.500 22.750 172.000 ;
        RECT 23.750 171.500 24.250 172.000 ;
        RECT 31.750 171.500 32.250 172.000 ;
        RECT 33.250 171.500 33.750 172.000 ;
        RECT 41.250 171.500 41.750 172.000 ;
        RECT 42.750 171.500 43.250 172.000 ;
        RECT 23.000 170.500 23.500 171.000 ;
        RECT 32.500 170.500 33.000 171.000 ;
        RECT 42.000 170.500 42.500 171.000 ;
        RECT 23.000 169.500 23.500 170.250 ;
        RECT 32.500 169.500 33.000 170.250 ;
        RECT 42.000 169.500 42.500 170.250 ;
        RECT 20.750 169.000 50.750 169.500 ;
        RECT 22.250 167.750 22.750 168.250 ;
        RECT 23.750 167.750 24.250 168.250 ;
        RECT 31.750 167.750 32.250 168.250 ;
        RECT 33.250 167.750 33.750 168.250 ;
        RECT 41.250 167.750 41.750 168.250 ;
        RECT 42.750 167.750 43.250 168.250 ;
        RECT 23.000 166.750 23.500 167.250 ;
        RECT 32.500 166.750 33.000 167.250 ;
        RECT 42.000 166.750 42.500 167.250 ;
        RECT 23.000 165.750 23.500 166.500 ;
        RECT 32.500 165.750 33.000 166.500 ;
        RECT 42.000 165.750 42.500 166.500 ;
        RECT 20.750 165.250 50.750 165.750 ;
        RECT 22.250 164.000 22.750 164.500 ;
        RECT 23.750 164.000 24.250 164.500 ;
        RECT 31.750 164.000 32.250 164.500 ;
        RECT 33.250 164.000 33.750 164.500 ;
        RECT 41.250 164.000 41.750 164.500 ;
        RECT 42.750 164.000 43.250 164.500 ;
        RECT 23.000 163.000 23.500 163.500 ;
        RECT 32.500 163.000 33.000 163.500 ;
        RECT 42.000 163.000 42.500 163.500 ;
        RECT 23.000 162.000 23.500 162.750 ;
        RECT 32.500 162.000 33.000 162.750 ;
        RECT 42.000 162.000 42.500 162.750 ;
        RECT 20.750 161.500 50.750 162.000 ;
        RECT 22.250 160.250 22.750 160.750 ;
        RECT 23.750 160.250 24.250 160.750 ;
        RECT 31.750 160.250 32.250 160.750 ;
        RECT 33.250 160.250 33.750 160.750 ;
        RECT 41.250 160.250 41.750 160.750 ;
        RECT 42.750 160.250 43.250 160.750 ;
        RECT 23.000 159.250 23.500 159.750 ;
        RECT 32.500 159.250 33.000 159.750 ;
        RECT 42.000 159.250 42.500 159.750 ;
        RECT 23.000 158.250 23.500 159.000 ;
        RECT 32.500 158.250 33.000 159.000 ;
        RECT 42.000 158.250 42.500 159.000 ;
        RECT 20.750 157.750 50.750 158.250 ;
        RECT 17.750 147.500 18.250 152.000 ;
        RECT 19.250 148.250 19.750 151.250 ;
        RECT 18.750 104.000 19.750 145.000 ;
        RECT 24.250 142.000 25.250 157.500 ;
        RECT 25.750 148.250 26.250 151.250 ;
        RECT 30.250 142.000 31.250 157.500 ;
        RECT 31.750 148.250 32.250 151.250 ;
        RECT 36.250 142.000 37.250 157.500 ;
        RECT 48.250 156.500 49.250 157.500 ;
        RECT 52.000 156.500 53.000 199.000 ;
        RECT 37.750 148.250 38.250 151.250 ;
        RECT 42.500 149.250 43.000 150.250 ;
        RECT 43.250 144.750 44.250 154.750 ;
        RECT 44.500 149.250 45.000 150.250 ;
        RECT 46.000 149.250 46.500 150.250 ;
        RECT 46.750 144.750 47.750 154.750 ;
        RECT 48.000 149.250 48.500 150.250 ;
        RECT 49.500 149.250 50.000 150.250 ;
        RECT 50.250 144.750 51.250 154.750 ;
        RECT 51.500 149.250 52.000 150.250 ;
        RECT 54.000 143.500 56.000 156.000 ;
        RECT 20.750 141.250 50.750 141.750 ;
        RECT 23.000 140.500 23.500 141.250 ;
        RECT 32.500 140.500 33.000 141.250 ;
        RECT 42.000 140.500 42.500 141.250 ;
        RECT 23.000 139.750 23.500 140.250 ;
        RECT 32.500 139.750 33.000 140.250 ;
        RECT 42.000 139.750 42.500 140.250 ;
        RECT 22.250 138.750 22.750 139.250 ;
        RECT 23.750 138.750 24.250 139.250 ;
        RECT 31.750 138.750 32.250 139.250 ;
        RECT 33.250 138.750 33.750 139.250 ;
        RECT 41.250 138.750 41.750 139.250 ;
        RECT 42.750 138.750 43.250 139.250 ;
        RECT 20.750 137.500 50.750 138.000 ;
        RECT 23.000 136.750 23.500 137.500 ;
        RECT 32.500 136.750 33.000 137.500 ;
        RECT 42.000 136.750 42.500 137.500 ;
        RECT 23.000 136.000 23.500 136.500 ;
        RECT 32.500 136.000 33.000 136.500 ;
        RECT 42.000 136.000 42.500 136.500 ;
        RECT 22.250 135.000 22.750 135.500 ;
        RECT 23.750 135.000 24.250 135.500 ;
        RECT 31.750 135.000 32.250 135.500 ;
        RECT 33.250 135.000 33.750 135.500 ;
        RECT 41.250 135.000 41.750 135.500 ;
        RECT 42.750 135.000 43.250 135.500 ;
        RECT 20.750 133.750 50.750 134.250 ;
        RECT 23.000 133.000 23.500 133.750 ;
        RECT 32.500 133.000 33.000 133.750 ;
        RECT 42.000 133.000 42.500 133.750 ;
        RECT 23.000 132.250 23.500 132.750 ;
        RECT 32.500 132.250 33.000 132.750 ;
        RECT 42.000 132.250 42.500 132.750 ;
        RECT 22.250 131.250 22.750 131.750 ;
        RECT 23.750 131.250 24.250 131.750 ;
        RECT 31.750 131.250 32.250 131.750 ;
        RECT 33.250 131.250 33.750 131.750 ;
        RECT 41.250 131.250 41.750 131.750 ;
        RECT 42.750 131.250 43.250 131.750 ;
        RECT 20.750 130.000 50.750 130.500 ;
        RECT 23.000 129.250 23.500 130.000 ;
        RECT 32.500 129.250 33.000 130.000 ;
        RECT 42.000 129.250 42.500 130.000 ;
        RECT 23.000 128.500 23.500 129.000 ;
        RECT 32.500 128.500 33.000 129.000 ;
        RECT 42.000 128.500 42.500 129.000 ;
        RECT 22.250 127.500 22.750 128.000 ;
        RECT 23.750 127.500 24.250 128.000 ;
        RECT 31.750 127.500 32.250 128.000 ;
        RECT 33.250 127.500 33.750 128.000 ;
        RECT 41.250 127.500 41.750 128.000 ;
        RECT 42.750 127.500 43.250 128.000 ;
        RECT 20.750 126.250 50.750 126.750 ;
        RECT 23.000 125.500 23.500 126.250 ;
        RECT 32.500 125.500 33.000 126.250 ;
        RECT 42.000 125.500 42.500 126.250 ;
        RECT 23.000 124.750 23.500 125.250 ;
        RECT 32.500 124.750 33.000 125.250 ;
        RECT 42.000 124.750 42.500 125.250 ;
        RECT 22.250 123.750 22.750 124.250 ;
        RECT 23.750 123.750 24.250 124.250 ;
        RECT 31.750 123.750 32.250 124.250 ;
        RECT 33.250 123.750 33.750 124.250 ;
        RECT 41.250 123.750 41.750 124.250 ;
        RECT 42.750 123.750 43.250 124.250 ;
        RECT 20.750 122.500 50.750 123.000 ;
        RECT 23.000 121.750 23.500 122.500 ;
        RECT 32.500 121.750 33.000 122.500 ;
        RECT 42.000 121.750 42.500 122.500 ;
        RECT 23.000 121.000 23.500 121.500 ;
        RECT 32.500 121.000 33.000 121.500 ;
        RECT 42.000 121.000 42.500 121.500 ;
        RECT 22.250 120.000 22.750 120.500 ;
        RECT 23.750 120.000 24.250 120.500 ;
        RECT 31.750 120.000 32.250 120.500 ;
        RECT 33.250 120.000 33.750 120.500 ;
        RECT 41.250 120.000 41.750 120.500 ;
        RECT 42.750 120.000 43.250 120.500 ;
        RECT 20.750 118.750 50.750 119.250 ;
        RECT 23.000 118.000 23.500 118.750 ;
        RECT 32.500 118.000 33.000 118.750 ;
        RECT 42.000 118.000 42.500 118.750 ;
        RECT 23.000 117.250 23.500 117.750 ;
        RECT 32.500 117.250 33.000 117.750 ;
        RECT 42.000 117.250 42.500 117.750 ;
        RECT 22.250 116.250 22.750 116.750 ;
        RECT 23.750 116.250 24.250 116.750 ;
        RECT 31.750 116.250 32.250 116.750 ;
        RECT 33.250 116.250 33.750 116.750 ;
        RECT 41.250 116.250 41.750 116.750 ;
        RECT 42.750 116.250 43.250 116.750 ;
        RECT 20.750 115.000 50.750 115.500 ;
        RECT 23.000 114.250 23.500 115.000 ;
        RECT 32.500 114.250 33.000 115.000 ;
        RECT 42.000 114.250 42.500 115.000 ;
        RECT 23.000 113.500 23.500 114.000 ;
        RECT 32.500 113.500 33.000 114.000 ;
        RECT 42.000 113.500 42.500 114.000 ;
        RECT 22.250 112.500 22.750 113.000 ;
        RECT 23.750 112.500 24.250 113.000 ;
        RECT 31.750 112.500 32.250 113.000 ;
        RECT 33.250 112.500 33.750 113.000 ;
        RECT 41.250 112.500 41.750 113.000 ;
        RECT 42.750 112.500 43.250 113.000 ;
        RECT 5.000 99.000 9.000 103.000 ;
        RECT 21.000 99.000 22.000 111.000 ;
        RECT 24.500 99.000 25.500 111.000 ;
        RECT 29.250 110.000 29.750 111.000 ;
        RECT 30.500 99.000 31.500 111.000 ;
        RECT 34.000 99.000 35.000 111.000 ;
        RECT 38.750 110.000 39.250 111.000 ;
        RECT 40.000 99.000 41.000 111.000 ;
        RECT 43.500 99.000 44.500 111.000 ;
        RECT 48.250 99.000 49.250 111.000 ;
        RECT 52.000 104.000 53.000 143.000 ;
        RECT 57.000 115.000 57.500 148.000 ;
        RECT 58.000 145.500 58.500 184.500 ;
        RECT 59.000 118.750 59.500 145.000 ;
        RECT 60.000 142.500 60.500 180.750 ;
        RECT 61.000 122.500 61.500 142.000 ;
        RECT 62.000 139.500 62.500 177.000 ;
        RECT 63.000 126.250 63.500 139.000 ;
        RECT 64.000 136.500 64.500 173.250 ;
        RECT 65.000 130.000 65.500 136.000 ;
        RECT 66.000 133.500 66.500 169.500 ;
        RECT 67.000 132.000 67.500 134.250 ;
        RECT 68.000 130.500 68.500 165.750 ;
        RECT 69.000 129.000 69.500 138.000 ;
        RECT 70.000 127.500 70.500 162.000 ;
        RECT 71.000 126.000 71.500 141.750 ;
        RECT 72.000 124.500 72.500 158.250 ;
        RECT 78.500 152.500 79.500 204.000 ;
        RECT 79.750 155.000 80.750 199.000 ;
        RECT 83.000 181.500 84.000 199.000 ;
        RECT 84.500 181.500 85.500 204.000 ;
        RECT 86.000 186.000 86.500 189.000 ;
        RECT 88.000 187.250 88.500 192.750 ;
        RECT 90.000 183.000 90.500 185.750 ;
        RECT 91.500 185.500 92.000 189.000 ;
        RECT 94.250 186.500 94.750 192.750 ;
        RECT 98.000 188.500 98.500 192.000 ;
        RECT 100.750 189.250 101.250 192.750 ;
        RECT 101.500 189.250 102.000 192.750 ;
        RECT 100.000 186.000 100.500 189.000 ;
        RECT 102.000 186.000 102.500 189.000 ;
        RECT 97.750 183.000 98.250 185.750 ;
        RECT 103.750 183.000 104.250 192.750 ;
        RECT 106.000 183.000 106.500 185.750 ;
        RECT 107.500 185.500 108.000 189.000 ;
        RECT 110.250 186.500 110.750 192.750 ;
        RECT 114.000 188.500 114.500 192.000 ;
        RECT 116.750 189.250 117.250 192.750 ;
        RECT 116.000 186.000 116.500 189.000 ;
        RECT 118.000 186.000 118.500 189.000 ;
        RECT 113.750 183.000 114.250 185.750 ;
        RECT 118.750 183.000 119.250 189.750 ;
        RECT 119.500 183.000 120.000 192.750 ;
        RECT 123.750 191.250 124.750 192.250 ;
        RECT 122.000 183.000 122.500 185.750 ;
        RECT 123.500 185.500 124.000 189.000 ;
        RECT 126.250 186.500 126.750 192.750 ;
        RECT 130.000 188.500 130.500 192.000 ;
        RECT 132.750 189.250 133.250 192.750 ;
        RECT 132.000 186.000 132.500 189.000 ;
        RECT 129.750 183.000 130.250 185.750 ;
        RECT 134.000 181.500 135.000 199.000 ;
        RECT 135.500 182.500 136.500 204.000 ;
        RECT 135.500 181.500 139.750 182.500 ;
        RECT 81.250 128.500 82.250 175.500 ;
        RECT 83.000 171.250 83.500 176.250 ;
        RECT 83.750 168.750 84.250 173.250 ;
        RECT 87.750 172.750 88.250 175.750 ;
        RECT 87.500 169.250 88.000 171.750 ;
        RECT 77.500 127.500 82.250 128.500 ;
        RECT 77.500 119.250 78.500 127.500 ;
        RECT 82.750 126.500 83.750 168.500 ;
        RECT 89.250 164.750 89.750 176.250 ;
        RECT 91.250 175.750 91.750 178.750 ;
        RECT 91.000 172.750 91.500 174.750 ;
        RECT 91.750 165.000 92.250 169.250 ;
        RECT 87.500 164.250 89.750 164.750 ;
        RECT 87.500 163.000 88.000 164.250 ;
        RECT 80.500 125.500 83.750 126.500 ;
        RECT 80.500 119.250 81.500 125.500 ;
        RECT 77.000 116.250 77.500 117.250 ;
        RECT 77.750 115.500 78.250 119.250 ;
        RECT 78.500 116.250 79.000 117.250 ;
        RECT 80.000 116.250 80.500 117.250 ;
        RECT 80.750 115.500 81.250 119.250 ;
        RECT 81.500 116.250 82.000 117.250 ;
        RECT 76.250 99.000 77.500 115.250 ;
        RECT 81.500 99.000 82.750 115.250 ;
        RECT 83.750 104.000 85.000 124.500 ;
        RECT 85.250 99.000 86.500 124.500 ;
        RECT 86.750 109.000 88.000 163.000 ;
        RECT 91.750 158.000 92.250 161.500 ;
        RECT 92.500 157.250 93.000 177.390 ;
        RECT 95.000 175.750 95.500 179.500 ;
        RECT 97.000 175.750 97.500 179.500 ;
        RECT 97.750 175.750 98.250 178.750 ;
        RECT 98.750 175.250 99.250 178.750 ;
        RECT 100.750 175.750 101.250 176.250 ;
        RECT 103.500 175.750 104.000 180.250 ;
        RECT 104.250 175.750 104.750 178.750 ;
        RECT 105.000 175.000 105.500 179.500 ;
        RECT 108.000 175.750 108.500 179.500 ;
        RECT 110.000 175.750 110.500 179.500 ;
        RECT 110.750 175.750 111.250 178.750 ;
        RECT 111.750 175.250 112.250 178.750 ;
        RECT 113.750 175.750 114.250 176.250 ;
        RECT 93.250 168.750 93.750 169.250 ;
        RECT 95.250 168.250 95.750 171.750 ;
        RECT 96.250 168.750 96.750 171.750 ;
        RECT 97.000 168.750 97.500 172.500 ;
        RECT 99.000 168.750 99.500 172.500 ;
        RECT 102.000 168.000 102.500 172.500 ;
        RECT 102.750 168.750 103.250 171.750 ;
        RECT 103.000 165.750 103.500 167.750 ;
        RECT 104.000 165.750 104.500 174.750 ;
        RECT 104.750 168.750 105.250 173.250 ;
        RECT 106.250 168.750 106.750 169.250 ;
        RECT 108.250 168.250 108.750 171.750 ;
        RECT 109.250 168.750 109.750 171.750 ;
        RECT 110.000 168.750 110.500 172.500 ;
        RECT 112.000 168.750 112.500 172.500 ;
        RECT 115.000 168.000 115.500 179.500 ;
        RECT 115.750 174.250 116.250 180.250 ;
        RECT 116.500 172.750 117.000 176.250 ;
        RECT 115.750 168.750 116.250 171.750 ;
        RECT 116.000 165.750 116.500 167.750 ;
        RECT 116.750 165.750 117.250 171.750 ;
        RECT 117.500 165.000 118.000 177.000 ;
        RECT 108.500 161.750 109.000 164.750 ;
        RECT 112.500 158.750 113.000 161.500 ;
        RECT 116.750 161.250 117.250 164.750 ;
        RECT 118.250 159.500 118.750 174.000 ;
        RECT 119.000 163.500 119.500 178.000 ;
        RECT 119.750 175.750 120.250 176.250 ;
        RECT 122.750 172.750 123.250 176.250 ;
        RECT 120.500 170.500 121.000 171.000 ;
        RECT 120.000 158.000 120.500 169.250 ;
        RECT 124.000 168.750 124.500 172.500 ;
        RECT 121.500 161.750 122.000 164.750 ;
        RECT 120.750 158.750 121.250 161.500 ;
        RECT 123.750 157.250 124.250 164.750 ;
        RECT 125.250 159.500 125.750 174.000 ;
        RECT 126.000 163.500 126.500 178.000 ;
        RECT 127.000 177.500 127.500 178.000 ;
        RECT 128.000 175.750 128.500 176.250 ;
        RECT 127.000 170.500 127.500 171.000 ;
        RECT 128.000 168.750 128.500 169.250 ;
        RECT 133.000 168.250 133.500 176.250 ;
        RECT 133.750 172.000 134.250 176.250 ;
        RECT 134.500 172.750 135.000 174.750 ;
        RECT 135.750 168.750 136.250 175.500 ;
        RECT 136.500 168.750 137.000 171.750 ;
        RECT 137.500 171.250 138.000 176.250 ;
        RECT 127.750 158.750 128.250 161.500 ;
        RECT 129.250 161.250 129.750 164.750 ;
        RECT 131.750 162.250 132.250 165.500 ;
        RECT 137.500 165.000 138.000 169.250 ;
        RECT 137.750 161.750 138.250 164.750 ;
        RECT 135.500 158.750 136.000 161.500 ;
        RECT 130.750 150.000 132.750 158.500 ;
        RECT 138.750 152.500 139.750 181.500 ;
        RECT 140.000 155.000 141.000 181.500 ;
        RECT 141.250 157.250 142.500 161.500 ;
        RECT 89.770 114.250 90.270 120.000 ;
        RECT 90.520 117.250 91.020 120.750 ;
        RECT 90.520 113.500 91.020 116.250 ;
        RECT 92.180 114.250 92.680 120.000 ;
        RECT 92.930 113.500 93.430 120.750 ;
        RECT 93.840 118.000 94.340 120.750 ;
        RECT 93.840 110.500 94.340 116.250 ;
        RECT 94.590 114.250 95.090 120.000 ;
        RECT 95.340 113.500 95.840 117.000 ;
        RECT 96.250 113.500 96.750 120.750 ;
        RECT 97.000 114.250 97.500 120.000 ;
        RECT 97.750 113.500 98.250 120.750 ;
        RECT 98.660 116.500 99.160 120.750 ;
        RECT 99.410 114.250 99.910 120.000 ;
        RECT 100.160 117.250 100.660 123.000 ;
        RECT 100.160 113.500 100.660 116.250 ;
        RECT 101.070 113.500 101.570 120.750 ;
        RECT 101.820 114.250 102.320 120.000 ;
        RECT 103.480 118.000 103.980 123.000 ;
        RECT 103.480 110.500 103.980 116.250 ;
        RECT 104.230 114.250 104.730 120.000 ;
        RECT 104.980 113.500 105.480 120.750 ;
        RECT 106.500 109.000 107.750 124.500 ;
        RECT 108.000 104.000 109.250 124.500 ;
        RECT 109.500 99.000 110.750 124.500 ;
        RECT 111.500 99.000 112.500 149.500 ;
        RECT 113.000 104.000 114.000 149.500 ;
        RECT 137.230 147.365 137.510 147.735 ;
        RECT 130.770 145.730 131.030 146.050 ;
        RECT 132.170 145.865 132.450 146.235 ;
        RECT 137.300 146.050 137.440 147.365 ;
        RECT 117.920 145.390 118.180 145.710 ;
        RECT 117.460 144.710 117.720 145.030 ;
        RECT 117.520 141.630 117.660 144.710 ;
        RECT 117.460 141.310 117.720 141.630 ;
        RECT 114.700 137.235 114.960 137.550 ;
        RECT 114.690 136.865 114.970 137.235 ;
        RECT 116.990 133.865 117.270 134.235 ;
        RECT 117.060 129.390 117.200 133.865 ;
        RECT 117.520 132.735 117.660 141.310 ;
        RECT 117.450 132.365 117.730 132.735 ;
        RECT 117.980 131.235 118.120 145.390 ;
        RECT 121.140 144.710 121.400 145.030 ;
        RECT 120.220 144.030 120.480 144.350 ;
        RECT 120.280 142.990 120.420 144.030 ;
        RECT 120.220 142.670 120.480 142.990 ;
        RECT 118.380 139.950 118.640 140.270 ;
        RECT 118.440 135.735 118.580 139.950 ;
        RECT 120.680 139.270 120.940 139.590 ;
        RECT 118.830 138.365 119.110 138.735 ;
        RECT 118.900 137.210 119.040 138.365 ;
        RECT 120.740 137.210 120.880 139.270 ;
        RECT 121.200 137.550 121.340 144.710 ;
        RECT 130.295 141.990 130.555 142.310 ;
        RECT 121.140 137.230 121.400 137.550 ;
        RECT 118.840 136.890 119.100 137.210 ;
        RECT 120.680 136.890 120.940 137.210 ;
        RECT 118.370 135.365 118.650 135.735 ;
        RECT 118.900 132.450 119.040 136.890 ;
        RECT 118.840 132.130 119.100 132.450 ;
        RECT 119.300 131.790 119.560 132.110 ;
        RECT 117.910 130.865 118.190 131.235 ;
        RECT 118.840 130.430 119.100 130.750 ;
        RECT 117.000 129.070 117.260 129.390 ;
        RECT 118.900 128.030 119.040 130.430 ;
        RECT 119.360 128.030 119.500 131.790 ;
        RECT 120.740 131.090 120.880 136.890 ;
        RECT 120.680 130.770 120.940 131.090 ;
        RECT 120.740 128.710 120.880 130.770 ;
        RECT 120.680 128.390 120.940 128.710 ;
        RECT 121.200 128.370 121.340 137.230 ;
        RECT 130.355 129.735 130.495 141.990 ;
        RECT 130.285 129.365 130.565 129.735 ;
        RECT 121.140 128.050 121.400 128.370 ;
        RECT 130.830 128.235 130.970 145.730 ;
        RECT 132.240 145.710 132.380 145.865 ;
        RECT 135.400 145.730 135.660 146.050 ;
        RECT 137.240 145.730 137.500 146.050 ;
        RECT 132.180 145.390 132.440 145.710 ;
        RECT 131.260 144.635 131.520 145.030 ;
        RECT 134.480 144.710 134.740 145.030 ;
        RECT 131.250 144.265 131.530 144.635 ;
        RECT 131.320 142.650 131.460 144.265 ;
        RECT 133.560 144.030 133.820 144.350 ;
        RECT 133.620 143.330 133.760 144.030 ;
        RECT 133.560 143.010 133.820 143.330 ;
        RECT 132.180 142.670 132.440 142.990 ;
        RECT 133.100 142.670 133.360 142.990 ;
        RECT 131.260 142.330 131.520 142.650 ;
        RECT 131.720 134.510 131.980 134.830 ;
        RECT 131.780 131.090 131.920 134.510 ;
        RECT 132.240 134.150 132.380 142.670 ;
        RECT 133.160 141.630 133.300 142.670 ;
        RECT 133.100 141.310 133.360 141.630 ;
        RECT 133.160 134.830 133.300 141.310 ;
        RECT 133.620 137.550 133.760 143.010 ;
        RECT 134.540 142.310 134.680 144.710 ;
        RECT 134.940 144.370 135.200 144.690 ;
        RECT 134.480 141.990 134.740 142.310 ;
        RECT 134.010 141.365 134.290 141.735 ;
        RECT 133.560 137.230 133.820 137.550 ;
        RECT 134.080 136.870 134.220 141.365 ;
        RECT 133.560 136.550 133.820 136.870 ;
        RECT 134.020 136.550 134.280 136.870 ;
        RECT 133.100 134.510 133.360 134.830 ;
        RECT 132.180 133.830 132.440 134.150 ;
        RECT 133.620 132.110 133.760 136.550 ;
        RECT 135.000 136.530 135.140 144.370 ;
        RECT 136.310 142.865 136.590 143.235 ;
        RECT 135.850 139.865 136.130 140.235 ;
        RECT 135.400 137.230 135.660 137.550 ;
        RECT 134.940 136.210 135.200 136.530 ;
        RECT 134.020 134.850 134.280 135.170 ;
        RECT 133.560 131.790 133.820 132.110 ;
        RECT 131.720 130.770 131.980 131.090 ;
        RECT 131.245 130.430 131.505 130.750 ;
        RECT 118.840 127.710 119.100 128.030 ;
        RECT 119.300 127.710 119.560 128.030 ;
        RECT 130.760 127.865 131.040 128.235 ;
        RECT 118.590 127.175 120.130 127.545 ;
        RECT 131.305 125.235 131.445 130.430 ;
        RECT 131.780 129.050 131.920 130.770 ;
        RECT 133.620 129.730 133.760 131.790 ;
        RECT 134.080 131.770 134.220 134.850 ;
        RECT 134.480 133.830 134.740 134.150 ;
        RECT 134.540 132.450 134.680 133.830 ;
        RECT 134.480 132.130 134.740 132.450 ;
        RECT 134.020 131.450 134.280 131.770 ;
        RECT 133.560 129.410 133.820 129.730 ;
        RECT 131.720 128.730 131.980 129.050 ;
        RECT 131.780 128.235 131.920 128.730 ;
        RECT 132.640 128.390 132.900 128.710 ;
        RECT 131.710 127.865 131.990 128.235 ;
        RECT 134.080 126.735 134.220 131.450 ;
        RECT 134.540 129.735 134.680 132.130 ;
        RECT 135.000 132.110 135.140 136.210 ;
        RECT 135.460 134.490 135.600 137.230 ;
        RECT 135.400 134.170 135.660 134.490 ;
        RECT 134.940 131.790 135.200 132.110 ;
        RECT 135.000 131.430 135.140 131.790 ;
        RECT 135.460 131.770 135.600 134.170 ;
        RECT 135.920 132.110 136.060 139.865 ;
        RECT 136.380 137.890 136.520 142.865 ;
        RECT 136.320 137.570 136.580 137.890 ;
        RECT 135.860 131.790 136.120 132.110 ;
        RECT 135.400 131.450 135.660 131.770 ;
        RECT 134.940 131.110 135.200 131.430 ;
        RECT 134.470 129.365 134.750 129.735 ;
        RECT 134.540 128.710 134.680 129.365 ;
        RECT 134.480 128.390 134.740 128.710 ;
        RECT 134.010 126.365 134.290 126.735 ;
        RECT 135.000 125.235 135.140 131.110 ;
        RECT 135.460 126.735 135.600 131.450 ;
        RECT 135.390 126.365 135.670 126.735 ;
        RECT 131.235 124.865 131.515 125.235 ;
        RECT 134.930 124.865 135.210 125.235 ;
        RECT 139.500 99.000 140.500 149.500 ;
        RECT 141.000 104.000 142.000 149.500 ;
        RECT 143.000 99.000 144.250 199.000 ;
        RECT 145.250 104.000 146.500 204.000 ;
      LAYER met3 ;
        RECT 5.000 223.500 89.000 224.500 ;
        RECT 0.000 200.000 4.000 204.000 ;
        RECT 5.000 195.000 9.000 199.000 ;
        RECT 123.750 191.250 132.750 192.250 ;
        RECT 144.500 190.250 160.500 190.500 ;
        RECT 29.250 188.500 29.750 189.500 ;
        RECT 38.750 188.500 39.250 189.500 ;
        RECT 48.250 188.500 49.250 189.500 ;
        RECT 94.000 189.250 160.500 190.250 ;
        RECT 144.500 189.000 160.500 189.250 ;
        RECT 144.500 188.250 145.500 188.500 ;
        RECT 22.250 186.500 22.750 187.000 ;
        RECT 23.750 186.500 24.250 187.000 ;
        RECT 21.250 185.500 23.500 186.000 ;
        RECT 25.590 185.100 29.750 187.500 ;
        RECT 31.750 186.500 32.250 187.000 ;
        RECT 33.250 186.500 33.750 187.000 ;
        RECT 30.750 185.500 33.000 186.000 ;
        RECT 35.090 185.100 39.250 187.500 ;
        RECT 41.250 186.500 41.750 187.000 ;
        RECT 42.750 186.500 43.250 187.000 ;
        RECT 40.250 185.500 42.500 186.000 ;
        RECT 44.590 185.100 48.750 187.500 ;
        RECT 88.000 187.250 147.500 188.250 ;
        RECT 144.500 187.000 145.500 187.250 ;
        RECT 22.250 182.750 22.750 183.250 ;
        RECT 23.750 182.750 24.250 183.250 ;
        RECT 21.250 181.750 23.500 182.250 ;
        RECT 25.590 181.350 29.750 183.750 ;
        RECT 31.750 182.750 32.250 183.250 ;
        RECT 33.250 182.750 33.750 183.250 ;
        RECT 30.750 181.750 33.000 182.250 ;
        RECT 35.090 181.350 39.250 183.750 ;
        RECT 41.250 182.750 41.750 183.250 ;
        RECT 42.750 182.750 43.250 183.250 ;
        RECT 40.250 181.750 42.500 182.250 ;
        RECT 44.590 181.350 48.750 183.750 ;
        RECT 22.250 179.000 22.750 179.500 ;
        RECT 23.750 179.000 24.250 179.500 ;
        RECT 21.250 178.000 23.500 178.500 ;
        RECT 25.590 177.600 29.750 180.000 ;
        RECT 31.750 179.000 32.250 179.500 ;
        RECT 33.250 179.000 33.750 179.500 ;
        RECT 30.750 178.000 33.000 178.500 ;
        RECT 35.090 177.600 39.250 180.000 ;
        RECT 41.250 179.000 41.750 179.500 ;
        RECT 42.750 179.000 43.250 179.500 ;
        RECT 40.250 178.000 42.500 178.500 ;
        RECT 44.590 177.600 48.750 180.000 ;
        RECT 22.250 175.250 22.750 175.750 ;
        RECT 23.750 175.250 24.250 175.750 ;
        RECT 21.250 174.250 23.500 174.750 ;
        RECT 25.590 173.850 29.750 176.250 ;
        RECT 31.750 175.250 32.250 175.750 ;
        RECT 33.250 175.250 33.750 175.750 ;
        RECT 30.750 174.250 33.000 174.750 ;
        RECT 35.090 173.850 39.250 176.250 ;
        RECT 41.250 175.250 41.750 175.750 ;
        RECT 42.750 175.250 43.250 175.750 ;
        RECT 40.250 174.250 42.500 174.750 ;
        RECT 44.590 173.850 48.750 176.250 ;
        RECT 100.500 175.500 101.500 176.500 ;
        RECT 113.500 175.500 114.500 176.500 ;
        RECT 119.000 175.750 120.250 176.250 ;
        RECT 122.250 173.600 127.500 178.000 ;
        RECT 128.000 175.750 128.500 176.250 ;
        RECT 22.250 171.500 22.750 172.000 ;
        RECT 23.750 171.500 24.250 172.000 ;
        RECT 21.250 170.500 23.500 171.000 ;
        RECT 25.590 170.100 29.750 172.500 ;
        RECT 31.750 171.500 32.250 172.000 ;
        RECT 33.250 171.500 33.750 172.000 ;
        RECT 30.750 170.500 33.000 171.000 ;
        RECT 35.090 170.100 39.250 172.500 ;
        RECT 41.250 171.500 41.750 172.000 ;
        RECT 42.750 171.500 43.250 172.000 ;
        RECT 40.250 170.500 42.500 171.000 ;
        RECT 44.590 170.100 48.750 172.500 ;
        RECT 22.250 167.750 22.750 168.250 ;
        RECT 23.750 167.750 24.250 168.250 ;
        RECT 21.250 166.750 23.500 167.250 ;
        RECT 25.590 166.350 29.750 168.750 ;
        RECT 31.750 167.750 32.250 168.250 ;
        RECT 33.250 167.750 33.750 168.250 ;
        RECT 30.750 166.750 33.000 167.250 ;
        RECT 35.090 166.350 39.250 168.750 ;
        RECT 41.250 167.750 41.750 168.250 ;
        RECT 42.750 167.750 43.250 168.250 ;
        RECT 40.250 166.750 42.500 167.250 ;
        RECT 44.590 166.350 48.750 168.750 ;
        RECT 93.000 168.500 94.000 169.500 ;
        RECT 106.000 168.500 107.000 169.500 ;
        RECT 115.750 166.600 121.000 171.000 ;
        RECT 122.250 166.600 127.500 171.000 ;
        RECT 128.000 168.750 128.500 169.250 ;
        RECT 22.250 164.000 22.750 164.500 ;
        RECT 23.750 164.000 24.250 164.500 ;
        RECT 21.250 163.000 23.500 163.500 ;
        RECT 25.590 162.600 29.750 165.000 ;
        RECT 31.750 164.000 32.250 164.500 ;
        RECT 33.250 164.000 33.750 164.500 ;
        RECT 30.750 163.000 33.000 163.500 ;
        RECT 35.090 162.600 39.250 165.000 ;
        RECT 41.250 164.000 41.750 164.500 ;
        RECT 42.750 164.000 43.250 164.500 ;
        RECT 40.250 163.000 42.500 163.500 ;
        RECT 44.590 162.600 48.750 165.000 ;
        RECT 100.500 162.000 154.500 163.000 ;
        RECT 22.250 160.250 22.750 160.750 ;
        RECT 23.750 160.250 24.250 160.750 ;
        RECT 21.250 159.250 23.500 159.750 ;
        RECT 25.590 158.850 29.750 161.250 ;
        RECT 31.750 160.250 32.250 160.750 ;
        RECT 33.250 160.250 33.750 160.750 ;
        RECT 30.750 159.250 33.000 159.750 ;
        RECT 35.090 158.850 39.250 161.250 ;
        RECT 41.250 160.250 41.750 160.750 ;
        RECT 42.750 160.250 43.250 160.750 ;
        RECT 40.250 159.250 42.500 159.750 ;
        RECT 44.590 158.850 48.750 161.250 ;
        RECT 113.500 160.500 153.000 161.500 ;
        RECT 106.000 159.000 151.500 160.000 ;
        RECT 93.000 157.500 150.000 158.500 ;
        RECT 20.750 156.500 25.250 157.500 ;
        RECT 30.250 156.500 31.250 157.500 ;
        RECT 36.250 156.500 40.750 157.500 ;
        RECT 48.250 156.500 49.250 157.500 ;
        RECT 12.250 155.250 56.000 156.000 ;
        RECT 36.750 154.250 50.750 154.750 ;
        RECT 30.750 153.250 47.250 153.750 ;
        RECT 24.750 152.250 43.750 152.750 ;
        RECT 24.750 150.750 38.250 151.250 ;
        RECT 9.500 150.250 12.750 150.750 ;
        RECT 9.500 149.250 13.250 150.250 ;
        RECT 13.750 149.500 18.250 150.000 ;
        RECT 19.250 149.500 24.750 150.000 ;
        RECT 25.750 149.500 30.750 150.000 ;
        RECT 31.750 149.500 36.750 150.000 ;
        RECT 9.500 148.750 12.750 149.250 ;
        RECT 42.500 149.000 75.500 150.500 ;
        RECT 130.750 150.000 132.750 152.000 ;
        RECT 24.750 148.250 38.250 148.750 ;
        RECT 57.000 147.700 112.750 148.000 ;
        RECT 137.205 147.700 137.535 147.715 ;
        RECT 57.000 147.400 137.535 147.700 ;
        RECT 24.750 146.750 43.750 147.250 ;
        RECT 57.000 147.000 112.750 147.400 ;
        RECT 137.205 147.385 137.535 147.400 ;
        RECT 30.750 145.750 47.250 146.250 ;
        RECT 58.000 146.200 112.750 146.500 ;
        RECT 132.145 146.200 132.475 146.215 ;
        RECT 58.000 145.900 132.475 146.200 ;
        RECT 58.000 145.500 112.750 145.900 ;
        RECT 132.145 145.885 132.475 145.900 ;
        RECT 36.750 144.750 50.750 145.250 ;
        RECT 59.000 144.600 112.750 145.000 ;
        RECT 131.225 144.600 131.555 144.615 ;
        RECT 59.000 144.300 131.555 144.600 ;
        RECT 12.250 143.500 56.000 144.250 ;
        RECT 59.000 144.000 112.750 144.300 ;
        RECT 131.225 144.285 131.555 144.300 ;
        RECT 60.000 143.200 112.750 143.500 ;
        RECT 136.285 143.200 136.615 143.215 ;
        RECT 20.750 142.000 25.250 143.000 ;
        RECT 30.250 142.000 31.250 143.000 ;
        RECT 36.250 142.000 40.750 143.000 ;
        RECT 60.000 142.900 136.615 143.200 ;
        RECT 60.000 142.500 112.750 142.900 ;
        RECT 136.285 142.885 136.615 142.900 ;
        RECT 61.000 141.700 112.750 142.000 ;
        RECT 133.985 141.700 134.315 141.715 ;
        RECT 61.000 141.400 134.315 141.700 ;
        RECT 61.000 141.000 112.750 141.400 ;
        RECT 133.985 141.385 134.315 141.400 ;
        RECT 21.250 139.750 23.500 140.250 ;
        RECT 22.250 138.750 22.750 139.250 ;
        RECT 23.750 138.750 24.250 139.250 ;
        RECT 25.590 138.250 29.750 140.650 ;
        RECT 30.750 139.750 33.000 140.250 ;
        RECT 31.750 138.750 32.250 139.250 ;
        RECT 33.250 138.750 33.750 139.250 ;
        RECT 35.090 138.250 39.250 140.650 ;
        RECT 40.250 139.750 42.500 140.250 ;
        RECT 41.250 138.750 41.750 139.250 ;
        RECT 42.750 138.750 43.250 139.250 ;
        RECT 44.590 138.250 48.750 140.650 ;
        RECT 62.000 140.200 112.750 140.500 ;
        RECT 135.825 140.200 136.155 140.215 ;
        RECT 62.000 139.900 136.155 140.200 ;
        RECT 62.000 139.500 112.750 139.900 ;
        RECT 135.825 139.885 136.155 139.900 ;
        RECT 63.000 138.700 112.750 139.000 ;
        RECT 118.805 138.700 119.135 138.715 ;
        RECT 63.000 138.400 119.135 138.700 ;
        RECT 63.000 138.000 112.750 138.400 ;
        RECT 118.805 138.385 119.135 138.400 ;
        RECT 64.000 137.200 112.750 137.500 ;
        RECT 114.665 137.200 114.995 137.215 ;
        RECT 64.000 136.900 114.995 137.200 ;
        RECT 21.250 136.000 23.500 136.500 ;
        RECT 22.250 135.000 22.750 135.500 ;
        RECT 23.750 135.000 24.250 135.500 ;
        RECT 25.590 134.500 29.750 136.900 ;
        RECT 30.750 136.000 33.000 136.500 ;
        RECT 31.750 135.000 32.250 135.500 ;
        RECT 33.250 135.000 33.750 135.500 ;
        RECT 35.090 134.500 39.250 136.900 ;
        RECT 40.250 136.000 42.500 136.500 ;
        RECT 41.250 135.000 41.750 135.500 ;
        RECT 42.750 135.000 43.250 135.500 ;
        RECT 44.590 134.500 48.750 136.900 ;
        RECT 64.000 136.500 112.750 136.900 ;
        RECT 114.665 136.885 114.995 136.900 ;
        RECT 65.000 135.700 112.750 136.000 ;
        RECT 118.345 135.700 118.675 135.715 ;
        RECT 65.000 135.400 118.675 135.700 ;
        RECT 65.000 135.000 112.750 135.400 ;
        RECT 118.345 135.385 118.675 135.400 ;
        RECT 66.000 134.200 112.750 134.500 ;
        RECT 116.965 134.200 117.295 134.215 ;
        RECT 66.000 133.900 117.295 134.200 ;
        RECT 66.000 133.500 112.750 133.900 ;
        RECT 116.965 133.885 117.295 133.900 ;
        RECT 21.250 132.250 23.500 132.750 ;
        RECT 22.250 131.250 22.750 131.750 ;
        RECT 23.750 131.250 24.250 131.750 ;
        RECT 25.590 130.750 29.750 133.150 ;
        RECT 30.750 132.250 33.000 132.750 ;
        RECT 31.750 131.250 32.250 131.750 ;
        RECT 33.250 131.250 33.750 131.750 ;
        RECT 35.090 130.750 39.250 133.150 ;
        RECT 40.250 132.250 42.500 132.750 ;
        RECT 41.250 131.250 41.750 131.750 ;
        RECT 42.750 131.250 43.250 131.750 ;
        RECT 44.590 130.750 48.750 133.150 ;
        RECT 67.000 132.700 112.750 133.000 ;
        RECT 117.425 132.700 117.755 132.715 ;
        RECT 67.000 132.400 117.755 132.700 ;
        RECT 67.000 132.000 112.750 132.400 ;
        RECT 117.425 132.385 117.755 132.400 ;
        RECT 68.000 131.200 112.750 131.500 ;
        RECT 117.885 131.200 118.215 131.215 ;
        RECT 68.000 130.900 118.215 131.200 ;
        RECT 68.000 130.500 112.750 130.900 ;
        RECT 117.885 130.885 118.215 130.900 ;
        RECT 69.000 129.700 112.750 130.000 ;
        RECT 130.260 129.700 130.590 129.715 ;
        RECT 69.000 129.400 130.590 129.700 ;
        RECT 21.250 128.500 23.500 129.000 ;
        RECT 22.250 127.500 22.750 128.000 ;
        RECT 23.750 127.500 24.250 128.000 ;
        RECT 25.590 127.000 29.750 129.400 ;
        RECT 30.750 128.500 33.000 129.000 ;
        RECT 31.750 127.500 32.250 128.000 ;
        RECT 33.250 127.500 33.750 128.000 ;
        RECT 35.090 127.000 39.250 129.400 ;
        RECT 40.250 128.500 42.500 129.000 ;
        RECT 41.250 127.500 41.750 128.000 ;
        RECT 42.750 127.500 43.250 128.000 ;
        RECT 44.590 127.000 48.750 129.400 ;
        RECT 69.000 129.000 112.750 129.400 ;
        RECT 130.260 129.385 130.590 129.400 ;
        RECT 134.445 129.700 134.775 129.715 ;
        RECT 142.500 129.700 147.500 130.000 ;
        RECT 134.445 129.400 147.500 129.700 ;
        RECT 134.445 129.385 134.775 129.400 ;
        RECT 142.500 129.000 147.500 129.400 ;
        RECT 70.000 128.200 112.750 128.500 ;
        RECT 130.735 128.200 131.065 128.215 ;
        RECT 70.000 127.900 131.065 128.200 ;
        RECT 70.000 127.500 112.750 127.900 ;
        RECT 130.735 127.885 131.065 127.900 ;
        RECT 131.685 128.200 132.015 128.215 ;
        RECT 142.500 128.200 147.500 128.500 ;
        RECT 131.685 127.900 147.500 128.200 ;
        RECT 131.685 127.885 132.015 127.900 ;
        RECT 118.570 127.195 120.150 127.525 ;
        RECT 142.500 127.500 147.500 127.900 ;
        RECT 71.000 126.700 112.750 127.000 ;
        RECT 133.985 126.700 134.315 126.715 ;
        RECT 71.000 126.400 134.315 126.700 ;
        RECT 71.000 126.000 112.750 126.400 ;
        RECT 133.985 126.385 134.315 126.400 ;
        RECT 135.365 126.700 135.695 126.715 ;
        RECT 142.500 126.700 147.500 127.000 ;
        RECT 135.365 126.400 147.500 126.700 ;
        RECT 135.365 126.385 135.695 126.400 ;
        RECT 142.500 126.000 147.500 126.400 ;
        RECT 21.250 124.750 23.500 125.250 ;
        RECT 22.250 123.750 22.750 124.250 ;
        RECT 23.750 123.750 24.250 124.250 ;
        RECT 25.590 123.250 29.750 125.650 ;
        RECT 30.750 124.750 33.000 125.250 ;
        RECT 31.750 123.750 32.250 124.250 ;
        RECT 33.250 123.750 33.750 124.250 ;
        RECT 35.090 123.250 39.250 125.650 ;
        RECT 40.250 124.750 42.500 125.250 ;
        RECT 41.250 123.750 41.750 124.250 ;
        RECT 42.750 123.750 43.250 124.250 ;
        RECT 44.590 123.250 48.750 125.650 ;
        RECT 72.000 125.200 112.750 125.500 ;
        RECT 131.210 125.200 131.540 125.215 ;
        RECT 72.000 124.900 131.540 125.200 ;
        RECT 72.000 124.500 112.750 124.900 ;
        RECT 131.210 124.885 131.540 124.900 ;
        RECT 134.905 125.200 135.235 125.215 ;
        RECT 142.500 125.200 148.500 125.500 ;
        RECT 134.905 124.900 148.500 125.200 ;
        RECT 134.905 124.885 135.235 124.900 ;
        RECT 142.500 124.500 148.500 124.900 ;
        RECT 21.250 121.000 23.500 121.500 ;
        RECT 22.250 120.000 22.750 120.500 ;
        RECT 23.750 120.000 24.250 120.500 ;
        RECT 25.590 119.500 29.750 121.900 ;
        RECT 30.750 121.000 33.000 121.500 ;
        RECT 31.750 120.000 32.250 120.500 ;
        RECT 33.250 120.000 33.750 120.500 ;
        RECT 35.090 119.500 39.250 121.900 ;
        RECT 40.250 121.000 42.500 121.500 ;
        RECT 41.250 120.000 41.750 120.500 ;
        RECT 42.750 120.000 43.250 120.500 ;
        RECT 44.590 119.500 48.750 121.900 ;
        RECT 21.250 117.250 23.500 117.750 ;
        RECT 22.250 116.250 22.750 116.750 ;
        RECT 23.750 116.250 24.250 116.750 ;
        RECT 25.590 115.750 29.750 118.150 ;
        RECT 30.750 117.250 33.000 117.750 ;
        RECT 31.750 116.250 32.250 116.750 ;
        RECT 33.250 116.250 33.750 116.750 ;
        RECT 35.090 115.750 39.250 118.150 ;
        RECT 40.250 117.250 42.500 117.750 ;
        RECT 41.250 116.250 41.750 116.750 ;
        RECT 42.750 116.250 43.250 116.750 ;
        RECT 44.590 115.750 48.750 118.150 ;
        RECT 73.500 115.750 77.500 117.750 ;
        RECT 78.500 115.750 80.500 117.750 ;
        RECT 81.500 115.750 98.250 117.750 ;
        RECT 106.500 117.500 147.500 117.750 ;
        RECT 106.500 116.000 157.500 117.500 ;
        RECT 106.500 115.750 147.500 116.000 ;
        RECT 21.250 113.500 23.500 114.000 ;
        RECT 22.250 112.500 22.750 113.000 ;
        RECT 23.750 112.500 24.250 113.000 ;
        RECT 25.590 112.000 29.750 114.400 ;
        RECT 30.750 113.500 33.000 114.000 ;
        RECT 31.750 112.500 32.250 113.000 ;
        RECT 33.250 112.500 33.750 113.000 ;
        RECT 35.090 112.000 39.250 114.400 ;
        RECT 40.250 113.500 42.500 114.000 ;
        RECT 41.250 112.500 41.750 113.000 ;
        RECT 42.750 112.500 43.250 113.000 ;
        RECT 44.590 112.000 48.750 114.400 ;
        RECT 29.250 110.000 29.750 111.000 ;
        RECT 38.750 110.000 39.250 111.000 ;
        RECT 48.250 110.000 49.250 111.000 ;
        RECT 0.000 104.000 4.000 108.000 ;
        RECT 5.000 99.000 9.000 103.000 ;
        RECT 73.500 100.000 151.500 102.000 ;
        RECT 7.840 76.600 30.000 97.000 ;
        RECT 31.340 76.600 53.500 97.000 ;
        RECT 54.840 76.600 77.000 97.000 ;
        RECT 78.340 76.600 100.500 97.000 ;
        RECT 101.840 76.600 124.000 97.000 ;
        RECT 125.340 76.600 147.500 97.000 ;
        RECT 7.840 54.600 30.000 75.000 ;
        RECT 31.340 54.600 53.500 75.000 ;
        RECT 54.840 54.600 77.000 75.000 ;
        RECT 78.340 54.600 100.500 75.000 ;
        RECT 101.840 54.600 124.000 75.000 ;
        RECT 125.340 54.600 147.500 75.000 ;
        RECT 31.340 32.600 53.500 53.000 ;
        RECT 54.840 32.600 77.000 53.000 ;
        RECT 78.340 32.600 100.500 53.000 ;
        RECT 101.840 32.600 124.000 53.000 ;
        RECT 125.340 32.600 147.500 53.000 ;
        RECT 31.340 10.600 53.500 31.000 ;
        RECT 54.840 10.600 77.000 31.000 ;
        RECT 78.340 10.600 100.500 31.000 ;
        RECT 101.840 10.600 124.000 31.000 ;
        RECT 125.340 10.600 147.500 31.000 ;
      LAYER met4 ;
        RECT 30.500 223.500 31.500 224.760 ;
        RECT 33.000 223.500 34.000 224.760 ;
        RECT 36.000 223.500 37.000 224.760 ;
        RECT 38.500 223.500 39.500 224.760 ;
        RECT 41.500 223.500 42.500 224.760 ;
        RECT 44.000 223.500 45.000 224.760 ;
        RECT 47.000 223.500 48.000 224.760 ;
        RECT 49.500 223.500 50.500 224.760 ;
        RECT 52.500 223.500 53.500 224.760 ;
        RECT 55.000 223.500 56.000 224.760 ;
        RECT 58.000 223.500 59.000 224.760 ;
        RECT 60.500 223.500 61.500 224.760 ;
        RECT 63.500 223.500 64.500 224.760 ;
        RECT 66.000 223.500 67.000 224.760 ;
        RECT 69.000 223.500 70.000 224.760 ;
        RECT 71.500 223.500 72.500 224.760 ;
        RECT 74.500 223.500 75.500 224.760 ;
        RECT 77.500 223.500 78.500 224.760 ;
        RECT 80.000 223.500 81.000 224.760 ;
        RECT 82.500 223.500 83.500 224.760 ;
        RECT 85.500 223.500 86.500 224.760 ;
        RECT 88.000 223.500 89.000 224.760 ;
        RECT 25.985 187.000 27.595 187.105 ;
        RECT 22.250 186.500 27.595 187.000 ;
        RECT 20.750 156.500 21.750 186.000 ;
        RECT 25.985 185.495 27.595 186.500 ;
        RECT 25.985 183.250 27.595 183.355 ;
        RECT 22.250 182.750 27.595 183.250 ;
        RECT 25.985 181.745 27.595 182.750 ;
        RECT 25.985 179.500 27.595 179.605 ;
        RECT 22.250 179.000 27.595 179.500 ;
        RECT 25.985 177.995 27.595 179.000 ;
        RECT 25.985 175.750 27.595 175.855 ;
        RECT 22.250 175.250 27.595 175.750 ;
        RECT 25.985 174.245 27.595 175.250 ;
        RECT 25.985 172.000 27.595 172.105 ;
        RECT 22.250 171.500 27.595 172.000 ;
        RECT 25.985 170.495 27.595 171.500 ;
        RECT 25.985 168.250 27.595 168.355 ;
        RECT 22.250 167.750 27.595 168.250 ;
        RECT 25.985 166.745 27.595 167.750 ;
        RECT 25.985 164.500 27.595 164.605 ;
        RECT 22.250 164.000 27.595 164.500 ;
        RECT 25.985 162.995 27.595 164.000 ;
        RECT 25.985 160.750 27.595 160.855 ;
        RECT 22.250 160.250 27.595 160.750 ;
        RECT 25.985 159.245 27.595 160.250 ;
        RECT 29.250 158.750 29.750 189.500 ;
        RECT 35.485 187.000 37.095 187.105 ;
        RECT 31.750 186.500 37.095 187.000 ;
        RECT 30.250 156.500 31.250 186.000 ;
        RECT 35.485 185.495 37.095 186.500 ;
        RECT 35.485 183.250 37.095 183.355 ;
        RECT 31.750 182.750 37.095 183.250 ;
        RECT 35.485 181.745 37.095 182.750 ;
        RECT 35.485 179.500 37.095 179.605 ;
        RECT 31.750 179.000 37.095 179.500 ;
        RECT 35.485 177.995 37.095 179.000 ;
        RECT 35.485 175.750 37.095 175.855 ;
        RECT 31.750 175.250 37.095 175.750 ;
        RECT 35.485 174.245 37.095 175.250 ;
        RECT 35.485 172.000 37.095 172.105 ;
        RECT 31.750 171.500 37.095 172.000 ;
        RECT 35.485 170.495 37.095 171.500 ;
        RECT 35.485 168.250 37.095 168.355 ;
        RECT 31.750 167.750 37.095 168.250 ;
        RECT 35.485 166.745 37.095 167.750 ;
        RECT 35.485 164.500 37.095 164.605 ;
        RECT 31.750 164.000 37.095 164.500 ;
        RECT 35.485 162.995 37.095 164.000 ;
        RECT 35.485 160.750 37.095 160.855 ;
        RECT 31.750 160.250 37.095 160.750 ;
        RECT 35.485 159.245 37.095 160.250 ;
        RECT 38.750 158.750 39.250 189.500 ;
        RECT 44.985 187.000 46.595 187.105 ;
        RECT 41.250 186.500 46.595 187.000 ;
        RECT 39.750 156.500 40.750 186.000 ;
        RECT 44.985 185.495 46.595 186.500 ;
        RECT 44.985 183.250 46.595 183.355 ;
        RECT 41.250 182.750 46.595 183.250 ;
        RECT 44.985 181.745 46.595 182.750 ;
        RECT 44.985 179.500 46.595 179.605 ;
        RECT 41.250 179.000 46.595 179.500 ;
        RECT 44.985 177.995 46.595 179.000 ;
        RECT 44.985 175.750 46.595 175.855 ;
        RECT 41.250 175.250 46.595 175.750 ;
        RECT 44.985 174.245 46.595 175.250 ;
        RECT 44.985 172.000 46.595 172.105 ;
        RECT 41.250 171.500 46.595 172.000 ;
        RECT 44.985 170.495 46.595 171.500 ;
        RECT 44.985 168.250 46.595 168.355 ;
        RECT 41.250 167.750 46.595 168.250 ;
        RECT 44.985 166.745 46.595 167.750 ;
        RECT 44.985 164.500 46.595 164.605 ;
        RECT 41.250 164.000 46.595 164.500 ;
        RECT 44.985 162.995 46.595 164.000 ;
        RECT 44.985 160.750 46.595 160.855 ;
        RECT 41.250 160.250 46.595 160.750 ;
        RECT 44.985 159.245 46.595 160.250 ;
        RECT 20.750 113.500 21.750 143.000 ;
        RECT 25.985 139.250 27.595 140.255 ;
        RECT 22.250 138.750 27.595 139.250 ;
        RECT 25.985 138.645 27.595 138.750 ;
        RECT 25.985 135.500 27.595 136.505 ;
        RECT 22.250 135.000 27.595 135.500 ;
        RECT 25.985 134.895 27.595 135.000 ;
        RECT 25.985 131.750 27.595 132.755 ;
        RECT 22.250 131.250 27.595 131.750 ;
        RECT 25.985 131.145 27.595 131.250 ;
        RECT 25.985 128.000 27.595 129.005 ;
        RECT 22.250 127.500 27.595 128.000 ;
        RECT 25.985 127.395 27.595 127.500 ;
        RECT 25.985 124.250 27.595 125.255 ;
        RECT 22.250 123.750 27.595 124.250 ;
        RECT 25.985 123.645 27.595 123.750 ;
        RECT 25.985 120.500 27.595 121.505 ;
        RECT 22.250 120.000 27.595 120.500 ;
        RECT 25.985 119.895 27.595 120.000 ;
        RECT 25.985 116.750 27.595 117.755 ;
        RECT 22.250 116.250 27.595 116.750 ;
        RECT 25.985 116.145 27.595 116.250 ;
        RECT 25.985 113.000 27.595 114.005 ;
        RECT 22.250 112.500 27.595 113.000 ;
        RECT 25.985 112.395 27.595 112.500 ;
        RECT 29.250 110.000 29.750 140.750 ;
        RECT 30.250 113.500 31.250 143.000 ;
        RECT 35.485 139.250 37.095 140.255 ;
        RECT 31.750 138.750 37.095 139.250 ;
        RECT 35.485 138.645 37.095 138.750 ;
        RECT 35.485 135.500 37.095 136.505 ;
        RECT 31.750 135.000 37.095 135.500 ;
        RECT 35.485 134.895 37.095 135.000 ;
        RECT 35.485 131.750 37.095 132.755 ;
        RECT 31.750 131.250 37.095 131.750 ;
        RECT 35.485 131.145 37.095 131.250 ;
        RECT 35.485 128.000 37.095 129.005 ;
        RECT 31.750 127.500 37.095 128.000 ;
        RECT 35.485 127.395 37.095 127.500 ;
        RECT 35.485 124.250 37.095 125.255 ;
        RECT 31.750 123.750 37.095 124.250 ;
        RECT 35.485 123.645 37.095 123.750 ;
        RECT 35.485 120.500 37.095 121.505 ;
        RECT 31.750 120.000 37.095 120.500 ;
        RECT 35.485 119.895 37.095 120.000 ;
        RECT 35.485 116.750 37.095 117.755 ;
        RECT 31.750 116.250 37.095 116.750 ;
        RECT 35.485 116.145 37.095 116.250 ;
        RECT 35.485 113.000 37.095 114.005 ;
        RECT 31.750 112.500 37.095 113.000 ;
        RECT 35.485 112.395 37.095 112.500 ;
        RECT 38.750 110.000 39.250 140.750 ;
        RECT 39.750 113.500 40.750 143.000 ;
        RECT 44.985 139.250 46.595 140.255 ;
        RECT 41.250 138.750 46.595 139.250 ;
        RECT 44.985 138.645 46.595 138.750 ;
        RECT 44.985 135.500 46.595 136.505 ;
        RECT 41.250 135.000 46.595 135.500 ;
        RECT 44.985 134.895 46.595 135.000 ;
        RECT 44.985 131.750 46.595 132.755 ;
        RECT 41.250 131.250 46.595 131.750 ;
        RECT 44.985 131.145 46.595 131.250 ;
        RECT 44.985 128.000 46.595 129.005 ;
        RECT 41.250 127.500 46.595 128.000 ;
        RECT 44.985 127.395 46.595 127.500 ;
        RECT 44.985 124.250 46.595 125.255 ;
        RECT 41.250 123.750 46.595 124.250 ;
        RECT 44.985 123.645 46.595 123.750 ;
        RECT 44.985 120.500 46.595 121.505 ;
        RECT 41.250 120.000 46.595 120.500 ;
        RECT 44.985 119.895 46.595 120.000 ;
        RECT 44.985 116.750 46.595 117.755 ;
        RECT 41.250 116.250 46.595 116.750 ;
        RECT 44.985 116.145 46.595 116.250 ;
        RECT 44.985 113.000 46.595 114.005 ;
        RECT 41.250 112.500 46.595 113.000 ;
        RECT 44.985 112.395 46.595 112.500 ;
        RECT 48.250 110.000 49.250 189.500 ;
        RECT 90.500 187.250 92.000 224.760 ;
        RECT 94.000 189.250 95.500 224.760 ;
        RECT 118.500 206.000 119.500 224.760 ;
        RECT 121.500 208.000 122.500 224.760 ;
        RECT 124.000 210.000 125.000 224.760 ;
        RECT 127.000 212.000 128.000 224.760 ;
        RECT 130.000 215.000 131.000 224.760 ;
        RECT 132.500 217.000 133.500 224.760 ;
        RECT 135.500 219.000 136.500 224.760 ;
        RECT 138.000 221.000 139.000 224.760 ;
        RECT 143.500 224.000 145.000 224.760 ;
        RECT 143.500 222.000 157.500 224.000 ;
        RECT 138.000 220.000 154.500 221.000 ;
        RECT 135.500 218.000 153.000 219.000 ;
        RECT 132.500 216.000 151.500 217.000 ;
        RECT 130.000 214.000 150.000 215.000 ;
        RECT 127.000 211.000 148.500 212.000 ;
        RECT 124.000 209.000 147.000 210.000 ;
        RECT 121.500 207.000 145.500 208.000 ;
        RECT 118.500 205.000 144.000 206.000 ;
        RECT 93.000 157.500 94.000 169.500 ;
        RECT 100.500 162.000 101.500 176.500 ;
        RECT 106.000 159.000 107.000 169.500 ;
        RECT 113.500 160.500 114.500 176.500 ;
        RECT 122.645 176.250 126.255 177.605 ;
        RECT 119.000 170.605 119.500 176.250 ;
        RECT 122.645 175.750 128.500 176.250 ;
        RECT 122.645 173.995 126.255 175.750 ;
        RECT 116.145 166.995 119.755 170.605 ;
        RECT 122.645 169.250 126.255 170.605 ;
        RECT 122.645 168.750 128.500 169.250 ;
        RECT 122.645 166.995 126.255 168.750 ;
        RECT 73.500 102.000 75.500 150.500 ;
        RECT 130.750 150.000 132.750 192.250 ;
        RECT 143.000 129.000 144.000 205.000 ;
        RECT 144.500 127.500 145.500 207.000 ;
        RECT 146.000 126.000 147.000 209.000 ;
        RECT 147.500 124.500 148.500 211.000 ;
        RECT 149.000 157.500 150.000 214.000 ;
        RECT 150.500 159.000 151.500 216.000 ;
        RECT 152.000 160.500 153.000 218.000 ;
        RECT 153.500 162.000 154.500 220.000 ;
        RECT 19.000 100.000 75.500 102.000 ;
        RECT 19.000 96.605 21.000 100.000 ;
        RECT 78.250 99.500 80.750 118.500 ;
        RECT 155.500 116.000 157.500 222.000 ;
        RECT 42.500 97.500 138.500 99.500 ;
        RECT 9.995 76.995 29.605 96.605 ;
        RECT 19.000 74.605 21.000 76.995 ;
        RECT 9.995 54.995 29.605 74.605 ;
        RECT 19.000 54.500 21.000 54.995 ;
        RECT 30.500 10.000 32.500 97.000 ;
        RECT 42.500 96.605 44.500 97.500 ;
        RECT 33.495 76.995 53.105 96.605 ;
        RECT 42.500 74.605 44.500 76.995 ;
        RECT 33.495 54.995 53.105 74.605 ;
        RECT 42.500 52.605 44.500 54.995 ;
        RECT 33.495 32.995 53.105 52.605 ;
        RECT 42.500 30.605 44.500 32.995 ;
        RECT 33.495 10.995 53.105 30.605 ;
        RECT 42.500 10.500 44.500 10.995 ;
        RECT 54.000 10.000 56.000 97.000 ;
        RECT 66.000 96.605 68.000 97.500 ;
        RECT 56.995 76.995 76.605 96.605 ;
        RECT 66.000 74.605 68.000 76.995 ;
        RECT 56.995 54.995 76.605 74.605 ;
        RECT 66.000 52.605 68.000 54.995 ;
        RECT 56.995 32.995 76.605 52.605 ;
        RECT 66.000 30.605 68.000 32.995 ;
        RECT 56.995 10.995 76.605 30.605 ;
        RECT 66.000 10.500 68.000 10.995 ;
        RECT 77.500 10.000 79.500 97.000 ;
        RECT 89.500 96.605 91.500 97.500 ;
        RECT 80.495 76.995 100.105 96.605 ;
        RECT 89.500 74.605 91.500 76.995 ;
        RECT 80.495 54.995 100.105 74.605 ;
        RECT 89.500 52.605 91.500 54.995 ;
        RECT 80.495 32.995 100.105 52.605 ;
        RECT 89.500 30.605 91.500 32.995 ;
        RECT 80.495 10.995 100.105 30.605 ;
        RECT 89.500 10.500 91.500 10.995 ;
        RECT 101.000 10.000 103.000 97.000 ;
        RECT 113.000 96.605 115.000 97.500 ;
        RECT 103.995 76.995 123.605 96.605 ;
        RECT 113.000 74.605 115.000 76.995 ;
        RECT 103.995 54.995 123.605 74.605 ;
        RECT 113.000 52.605 115.000 54.995 ;
        RECT 103.995 32.995 123.605 52.605 ;
        RECT 113.000 30.605 115.000 32.995 ;
        RECT 103.995 10.995 123.605 30.605 ;
        RECT 113.000 10.500 115.000 10.995 ;
        RECT 124.500 10.000 126.500 97.000 ;
        RECT 136.500 96.605 138.500 97.500 ;
        RECT 127.495 76.995 147.105 96.605 ;
        RECT 136.500 74.605 138.500 76.995 ;
        RECT 127.495 54.995 147.105 74.605 ;
        RECT 136.500 52.605 138.500 54.995 ;
        RECT 127.495 32.995 147.105 52.605 ;
        RECT 136.500 30.605 138.500 32.995 ;
        RECT 127.495 10.995 147.105 30.605 ;
        RECT 136.500 10.500 138.500 10.995 ;
        RECT 9.000 8.000 126.500 10.000 ;
        RECT 149.500 8.000 151.500 102.000 ;
        RECT 132.000 6.000 151.500 8.000 ;
        RECT 132.000 1.000 134.000 6.000 ;
        RECT 158.500 4.000 160.500 190.500 ;
        RECT 151.500 2.000 160.500 4.000 ;
        RECT 151.500 1.000 153.500 2.000 ;
  END
END tt_um_assaify_mssf_pll
END LIBRARY

