module tt_um_SNPU (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;

 sky130_fd_sc_hd__mux4_1 _219_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_170_));
 sky130_fd_sc_hd__mux4_1 _220_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(_171_),
    .A1(_170_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_172_));
 sky130_fd_sc_hd__and2b_1 _222_ (.A_N(net15),
    .B(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_173_));
 sky130_fd_sc_hd__mux4_1 _223_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_174_));
 sky130_fd_sc_hd__mux4_1 _224_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _225_ (.A0(_174_),
    .A1(_175_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_176_));
 sky130_fd_sc_hd__a21o_1 _226_ (.A1(net15),
    .A2(_176_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_177_));
 sky130_fd_sc_hd__o22a_4 _227_ (.A1(net7),
    .A2(_169_),
    .B1(_173_),
    .B2(_177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__nand2b_1 _228_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _229_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _230_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _231_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _232_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _233_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _234_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _235_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _236_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _237_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _238_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _239_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _240_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _241_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _242_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _243_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _244_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _245_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _246_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _247_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _248_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _249_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _250_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _251_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _252_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _253_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _254_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _255_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _256_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _257_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _258_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _259_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _260_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_178_));
 sky130_fd_sc_hd__mux4_1 _261_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_179_));
 sky130_fd_sc_hd__mux4_1 _262_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_180_));
 sky130_fd_sc_hd__mux4_1 _263_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_181_));
 sky130_fd_sc_hd__mux4_1 _264_ (.A0(_179_),
    .A1(_181_),
    .A2(_178_),
    .A3(_180_),
    .S0(net15),
    .S1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_182_));
 sky130_fd_sc_hd__mux4_1 _265_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_183_));
 sky130_fd_sc_hd__mux4_1 _266_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(_184_),
    .A1(_183_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_185_));
 sky130_fd_sc_hd__mux4_1 _268_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_186_));
 sky130_fd_sc_hd__mux4_1 _269_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_187_));
 sky130_fd_sc_hd__mux2_1 _270_ (.A0(_187_),
    .A1(_186_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_188_));
 sky130_fd_sc_hd__and2b_1 _271_ (.A_N(net15),
    .B(_188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_189_));
 sky130_fd_sc_hd__a21o_1 _272_ (.A1(net15),
    .A2(_185_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_190_));
 sky130_fd_sc_hd__o22a_4 _273_ (.A1(net7),
    .A2(_182_),
    .B1(_189_),
    .B2(_190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__nand2b_1 _274_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _275_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _276_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _277_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _278_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _279_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _280_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _281_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _282_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _283_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _284_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _285_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _286_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _287_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _288_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _289_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _290_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _291_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _292_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _293_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _294_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _295_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _296_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _297_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _298_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _299_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _300_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _301_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _302_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _303_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _304_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _305_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _306_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_191_));
 sky130_fd_sc_hd__mux4_1 _307_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_192_));
 sky130_fd_sc_hd__mux4_1 _308_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_193_));
 sky130_fd_sc_hd__mux4_1 _309_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_194_));
 sky130_fd_sc_hd__mux4_1 _310_ (.A0(_192_),
    .A1(_194_),
    .A2(_191_),
    .A3(_193_),
    .S0(net12),
    .S1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_195_));
 sky130_fd_sc_hd__mux4_1 _311_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_196_));
 sky130_fd_sc_hd__mux4_1 _312_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_197_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(_197_),
    .A1(_196_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_198_));
 sky130_fd_sc_hd__and2b_1 _314_ (.A_N(net12),
    .B(_198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_199_));
 sky130_fd_sc_hd__mux4_1 _315_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_200_));
 sky130_fd_sc_hd__mux4_1 _316_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(_200_),
    .A1(_201_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_202_));
 sky130_fd_sc_hd__a21o_1 _318_ (.A1(net12),
    .A2(_202_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_203_));
 sky130_fd_sc_hd__o22a_4 _319_ (.A1(net7),
    .A2(_195_),
    .B1(_199_),
    .B2(_203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__nand2b_1 _320_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _321_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _322_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _323_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _324_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _325_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _326_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _327_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _328_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _329_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _330_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _331_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _332_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _333_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _334_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _335_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _336_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _337_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _338_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _339_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _340_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _341_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _342_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _343_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _344_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _345_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _346_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _347_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _348_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _349_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _350_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _351_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _352_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_204_));
 sky130_fd_sc_hd__mux4_1 _353_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(_205_),
    .A1(_204_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_206_));
 sky130_fd_sc_hd__mux4_1 _355_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_207_));
 sky130_fd_sc_hd__mux4_1 _356_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_208_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(_208_),
    .A1(_207_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_209_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(_206_),
    .A1(_209_),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_210_));
 sky130_fd_sc_hd__mux4_1 _359_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_211_));
 sky130_fd_sc_hd__mux4_1 _360_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_212_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(_212_),
    .A1(_211_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_213_));
 sky130_fd_sc_hd__and2b_1 _362_ (.A_N(net14),
    .B(_213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_214_));
 sky130_fd_sc_hd__mux4_1 _363_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_215_));
 sky130_fd_sc_hd__mux4_1 _364_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_216_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(_215_),
    .A1(_216_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_217_));
 sky130_fd_sc_hd__a21o_1 _366_ (.A1(net14),
    .A2(_217_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_218_));
 sky130_fd_sc_hd__o22a_4 _367_ (.A1(net8),
    .A2(_210_),
    .B1(_214_),
    .B2(_218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 _368_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hd__nand2b_1 _369_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _370_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _371_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _372_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _373_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _374_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _375_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _376_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _377_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _378_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _379_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _380_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _381_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _382_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _383_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _384_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _385_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _386_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _387_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _388_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _389_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _390_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _391_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _392_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _393_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _394_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _395_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _396_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _397_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _398_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _399_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _400_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _401_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__mux4_1 _402_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(_001_),
    .A1(_002_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__mux4_1 _404_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net54),
    .S1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__mux4_1 _405_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net54),
    .S1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(_005_),
    .A1(_004_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(_006_),
    .A1(_003_),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__mux4_1 _408_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__mux4_1 _409_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(_009_),
    .A1(_008_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__and2b_1 _411_ (.A_N(net11),
    .B(_010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__mux4_1 _412_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__mux4_1 _413_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(_012_),
    .A1(_013_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__a21o_1 _415_ (.A1(net14),
    .A2(_014_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__o22a_4 _416_ (.A1(net7),
    .A2(_007_),
    .B1(_011_),
    .B2(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__nand2b_1 _417_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _418_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _419_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _420_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _421_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _422_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _423_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _424_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _425_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _426_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _427_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _428_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _429_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _430_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _431_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _432_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _433_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _434_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _435_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _436_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _437_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _438_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _439_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _440_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _441_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _442_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _443_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _444_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _445_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _446_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _447_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _448_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _449_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__mux4_1 _450_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(_016_),
    .A1(_017_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__mux4_1 _452_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__mux4_1 _453_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(_020_),
    .A1(_019_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(_021_),
    .A1(_018_),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_022_));
 sky130_fd_sc_hd__mux4_1 _456_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__mux4_1 _457_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(_024_),
    .A1(_023_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__and2b_1 _459_ (.A_N(net14),
    .B(_025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__mux4_1 _460_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__mux4_1 _461_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net51),
    .S1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(_027_),
    .A1(_028_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__a21o_1 _463_ (.A1(net14),
    .A2(_029_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__o22a_4 _464_ (.A1(net8),
    .A2(_022_),
    .B1(_026_),
    .B2(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__nand2b_1 _465_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _466_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _467_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _468_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _469_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _470_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _471_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _472_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _473_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _474_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _475_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _476_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _477_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _478_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _479_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _480_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _481_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _482_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _483_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _484_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _485_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _486_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _487_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _488_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _489_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _490_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _491_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _492_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _493_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _494_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _495_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _496_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _497_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__mux4_1 _498_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(_032_),
    .A1(_031_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__mux4_1 _500_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__mux4_1 _501_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(_035_),
    .A1(_034_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(_033_),
    .A1(_036_),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__mux4_1 _504_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__mux4_1 _505_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(_039_),
    .A1(_038_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__mux4_1 _507_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__mux4_1 _508_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net44),
    .S1(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _509_ (.A0(_042_),
    .A1(_041_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__and2b_1 _510_ (.A_N(net13),
    .B(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__a21o_1 _511_ (.A1(net13),
    .A2(_040_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__o22a_4 _512_ (.A1(net7),
    .A2(_037_),
    .B1(_044_),
    .B2(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__nand2b_1 _513_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _514_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _515_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _516_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _517_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _518_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _519_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _520_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _521_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _522_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _523_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _524_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _525_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _526_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _527_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _528_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _529_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _530_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _531_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _532_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _533_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _534_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _535_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _536_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _537_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _538_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _539_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _540_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _541_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _542_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _543_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _544_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _545_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__mux4_1 _546_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__mux4_1 _547_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__mux4_1 _548_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net47),
    .S1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__mux4_1 _549_ (.A0(_047_),
    .A1(_049_),
    .A2(_046_),
    .A3(_048_),
    .S0(net12),
    .S1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__mux4_1 _550_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__mux4_1 _551_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _552_ (.A0(_052_),
    .A1(_051_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__mux4_1 _553_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__mux4_1 _554_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net49),
    .S1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(_055_),
    .A1(_054_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__and2b_1 _556_ (.A_N(net12),
    .B(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__a21o_1 _557_ (.A1(net12),
    .A2(_053_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__o22a_4 _558_ (.A1(net7),
    .A2(_050_),
    .B1(_057_),
    .B2(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__nand2b_1 _559_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _560_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _561_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _562_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _563_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _564_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _565_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _566_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _567_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _568_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _569_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _570_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _571_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _572_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _573_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _574_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _575_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _576_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _577_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _578_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _579_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _580_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _581_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _582_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _583_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _584_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _585_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _586_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _587_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _588_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _589_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _590_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _591_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__mux4_1 _592_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_060_));
 sky130_fd_sc_hd__mux4_1 _593_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__mux4_1 _594_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_062_));
 sky130_fd_sc_hd__mux4_1 _595_ (.A0(_060_),
    .A1(_062_),
    .A2(_059_),
    .A3(_061_),
    .S0(net12),
    .S1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__mux4_1 _596_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_064_));
 sky130_fd_sc_hd__mux4_1 _597_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net48),
    .S1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _598_ (.A0(_065_),
    .A1(_064_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__mux4_1 _599_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__mux4_1 _600_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _601_ (.A0(_068_),
    .A1(_067_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__and2b_1 _602_ (.A_N(net12),
    .B(_069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__a21o_1 _603_ (.A1(net13),
    .A2(_066_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_071_));
 sky130_fd_sc_hd__o22a_4 _604_ (.A1(net7),
    .A2(_063_),
    .B1(_070_),
    .B2(_071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__nand2b_1 _605_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _606_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _607_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _608_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _609_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _610_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _611_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _612_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _613_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _614_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _615_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _616_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _617_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _618_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _619_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _620_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _621_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _622_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _623_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _624_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _625_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _626_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _627_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _628_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _629_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _630_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _631_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _632_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _633_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _634_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _635_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _636_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _637_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_072_));
 sky130_fd_sc_hd__mux4_1 _638_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_073_));
 sky130_fd_sc_hd__mux4_1 _639_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_074_));
 sky130_fd_sc_hd__mux4_1 _640_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_075_));
 sky130_fd_sc_hd__mux4_1 _641_ (.A0(_073_),
    .A1(_075_),
    .A2(_072_),
    .A3(_074_),
    .S0(net12),
    .S1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_076_));
 sky130_fd_sc_hd__mux4_1 _642_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_077_));
 sky130_fd_sc_hd__mux4_1 _643_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net46),
    .S1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _644_ (.A0(_078_),
    .A1(_077_),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_079_));
 sky130_fd_sc_hd__and2b_1 _645_ (.A_N(net12),
    .B(_079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_080_));
 sky130_fd_sc_hd__mux4_1 _646_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__mux4_1 _647_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _648_ (.A0(_081_),
    .A1(_082_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_083_));
 sky130_fd_sc_hd__a21o_1 _649_ (.A1(net11),
    .A2(_083_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_084_));
 sky130_fd_sc_hd__o22a_4 _650_ (.A1(net7),
    .A2(_076_),
    .B1(_080_),
    .B2(_084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__nand2b_1 _651_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _652_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _653_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _654_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _655_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _656_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _657_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _658_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _659_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _660_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _661_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _662_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _663_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _664_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _665_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _666_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _667_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _668_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _669_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _670_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _671_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _672_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _673_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _674_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _675_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _676_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _677_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _678_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _679_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _680_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _681_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _682_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _683_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_085_));
 sky130_fd_sc_hd__mux4_1 _684_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_086_));
 sky130_fd_sc_hd__mux4_1 _685_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_087_));
 sky130_fd_sc_hd__mux4_1 _686_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_088_));
 sky130_fd_sc_hd__mux4_1 _687_ (.A0(_086_),
    .A1(_088_),
    .A2(_085_),
    .A3(_087_),
    .S0(net11),
    .S1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_089_));
 sky130_fd_sc_hd__mux4_1 _688_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_090_));
 sky130_fd_sc_hd__mux4_1 _689_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net43),
    .S1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _690_ (.A0(_091_),
    .A1(_090_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_092_));
 sky130_fd_sc_hd__and2b_1 _691_ (.A_N(net11),
    .B(_092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_093_));
 sky130_fd_sc_hd__mux4_1 _692_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_094_));
 sky130_fd_sc_hd__mux4_1 _693_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net45),
    .S1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _694_ (.A0(_094_),
    .A1(_095_),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_096_));
 sky130_fd_sc_hd__a21o_1 _695_ (.A1(net11),
    .A2(_096_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_097_));
 sky130_fd_sc_hd__o22a_4 _696_ (.A1(net7),
    .A2(_089_),
    .B1(_093_),
    .B2(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__nand2b_1 _697_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _698_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _699_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _700_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _701_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _702_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _703_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _704_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _705_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _706_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _707_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _708_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _709_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _710_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _711_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _712_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _713_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _714_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _715_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _716_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _717_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _718_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _719_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _720_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _721_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _722_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _723_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _724_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _725_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _726_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _727_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _728_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _729_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_098_));
 sky130_fd_sc_hd__mux4_1 _730_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_099_));
 sky130_fd_sc_hd__mux4_1 _731_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_100_));
 sky130_fd_sc_hd__mux4_1 _732_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_101_));
 sky130_fd_sc_hd__mux4_1 _733_ (.A0(_099_),
    .A1(_101_),
    .A2(_098_),
    .A3(_100_),
    .S0(net11),
    .S1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_102_));
 sky130_fd_sc_hd__mux4_1 _734_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_103_));
 sky130_fd_sc_hd__mux4_1 _735_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _736_ (.A0(_104_),
    .A1(_103_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_105_));
 sky130_fd_sc_hd__mux4_1 _737_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_106_));
 sky130_fd_sc_hd__mux4_1 _738_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net42),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _739_ (.A0(_107_),
    .A1(_106_),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__and2b_1 _740_ (.A_N(net11),
    .B(_108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_109_));
 sky130_fd_sc_hd__a21o_1 _741_ (.A1(net11),
    .A2(_105_),
    .B1(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_110_));
 sky130_fd_sc_hd__o22a_4 _742_ (.A1(net7),
    .A2(_102_),
    .B1(_109_),
    .B2(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__nand2b_1 _743_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _744_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _745_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _746_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _747_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _748_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _749_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _750_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _751_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _752_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _753_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _754_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _755_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _756_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _757_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _758_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _759_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _760_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _761_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _762_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _763_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _764_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _765_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _766_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _767_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _768_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _769_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _770_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _771_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _772_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _773_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _774_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _775_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net54),
    .S1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_111_));
 sky130_fd_sc_hd__mux4_1 _776_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_112_));
 sky130_fd_sc_hd__mux4_1 _777_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net54),
    .S1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__mux4_1 _778_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_114_));
 sky130_fd_sc_hd__mux4_1 _779_ (.A0(_112_),
    .A1(_114_),
    .A2(_111_),
    .A3(_113_),
    .S0(net14),
    .S1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__mux4_1 _780_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__mux4_1 _781_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _782_ (.A0(_117_),
    .A1(_116_),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_118_));
 sky130_fd_sc_hd__and2b_1 _783_ (.A_N(net14),
    .B(_118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_119_));
 sky130_fd_sc_hd__mux4_1 _784_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_120_));
 sky130_fd_sc_hd__mux4_1 _785_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net53),
    .S1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _786_ (.A0(_120_),
    .A1(_121_),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__a21o_1 _787_ (.A1(net14),
    .A2(_122_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_123_));
 sky130_fd_sc_hd__o22a_4 _788_ (.A1(net8),
    .A2(_115_),
    .B1(_119_),
    .B2(_123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__nand2b_1 _789_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _790_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _791_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _792_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _793_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _794_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _795_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _796_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _797_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _798_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _799_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _800_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _801_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _802_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _803_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _804_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _805_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _806_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _807_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _808_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _809_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _810_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _811_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _812_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _813_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _814_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _815_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _816_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _817_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _818_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _819_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _820_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _821_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_124_));
 sky130_fd_sc_hd__mux4_1 _822_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__mux4_1 _823_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net55),
    .S1(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__mux4_1 _824_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_127_));
 sky130_fd_sc_hd__mux4_1 _825_ (.A0(_125_),
    .A1(_127_),
    .A2(_124_),
    .A3(_126_),
    .S0(net15),
    .S1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_128_));
 sky130_fd_sc_hd__mux4_1 _826_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__mux4_1 _827_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _828_ (.A0(_130_),
    .A1(_129_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_131_));
 sky130_fd_sc_hd__and2b_1 _829_ (.A_N(net15),
    .B(_131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_132_));
 sky130_fd_sc_hd__mux4_1 _830_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__mux4_1 _831_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _832_ (.A0(_133_),
    .A1(_134_),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_135_));
 sky130_fd_sc_hd__a21o_1 _833_ (.A1(net15),
    .A2(_135_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__o22a_4 _834_ (.A1(net8),
    .A2(_128_),
    .B1(_132_),
    .B2(_136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__nand2b_1 _835_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _836_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _837_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _838_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _839_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _840_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _841_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _842_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _843_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _844_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _845_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _846_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _847_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _848_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _849_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _850_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _851_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _852_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _853_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _854_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _855_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _856_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _857_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _858_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _859_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _860_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _861_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _862_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _863_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _864_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _865_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _866_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _867_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_137_));
 sky130_fd_sc_hd__mux4_1 _868_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _869_ (.A0(_138_),
    .A1(_137_),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_139_));
 sky130_fd_sc_hd__mux4_1 _870_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_140_));
 sky130_fd_sc_hd__mux4_1 _871_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _872_ (.A0(_141_),
    .A1(_140_),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _873_ (.A0(_139_),
    .A1(_142_),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_143_));
 sky130_fd_sc_hd__mux4_1 _874_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_144_));
 sky130_fd_sc_hd__mux4_1 _875_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _876_ (.A0(_145_),
    .A1(_144_),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_146_));
 sky130_fd_sc_hd__mux4_1 _877_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_147_));
 sky130_fd_sc_hd__mux4_1 _878_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net52),
    .S1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _879_ (.A0(_148_),
    .A1(_147_),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_149_));
 sky130_fd_sc_hd__and2b_1 _880_ (.A_N(net16),
    .B(_149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_150_));
 sky130_fd_sc_hd__a21o_1 _881_ (.A1(net16),
    .A2(_146_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_151_));
 sky130_fd_sc_hd__o22a_4 _882_ (.A1(net8),
    .A2(_143_),
    .B1(_150_),
    .B2(_151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__nand2b_1 _883_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _884_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _885_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _886_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _887_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _888_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _889_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _890_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _891_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _892_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _893_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _894_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _895_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _896_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _897_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _898_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _899_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _900_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _901_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _902_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _903_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _904_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _905_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _906_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _907_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _908_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _909_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _910_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _911_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _912_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _913_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _914_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _915_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_152_));
 sky130_fd_sc_hd__mux4_1 _916_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_153_));
 sky130_fd_sc_hd__mux4_1 _917_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net57),
    .S1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_154_));
 sky130_fd_sc_hd__mux4_1 _918_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net58),
    .S1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_155_));
 sky130_fd_sc_hd__mux4_1 _919_ (.A0(_153_),
    .A1(_155_),
    .A2(_152_),
    .A3(_154_),
    .S0(net15),
    .S1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_156_));
 sky130_fd_sc_hd__mux4_1 _920_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net58),
    .S1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_157_));
 sky130_fd_sc_hd__mux4_1 _921_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net58),
    .S1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _922_ (.A0(_158_),
    .A1(_157_),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_159_));
 sky130_fd_sc_hd__and2b_1 _923_ (.A_N(net16),
    .B(_159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_160_));
 sky130_fd_sc_hd__mux4_1 _924_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net58),
    .S1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_161_));
 sky130_fd_sc_hd__mux4_1 _925_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net58),
    .S1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _926_ (.A0(_161_),
    .A1(_162_),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_163_));
 sky130_fd_sc_hd__a21o_1 _927_ (.A1(net16),
    .A2(_163_),
    .B1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_164_));
 sky130_fd_sc_hd__o22a_4 _928_ (.A1(net8),
    .A2(_156_),
    .B1(_160_),
    .B2(_164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__nand2b_1 _929_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _930_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _931_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _932_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _933_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _934_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _935_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _936_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _937_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _938_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _939_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _940_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _941_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _942_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _943_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _944_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _945_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _946_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _947_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _948_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _949_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _950_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _951_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _952_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _953_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _954_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _955_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _956_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _957_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _958_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _959_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _960_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__mux4_1 _961_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_165_));
 sky130_fd_sc_hd__mux4_1 _962_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_166_));
 sky130_fd_sc_hd__mux4_1 _963_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_167_));
 sky130_fd_sc_hd__mux4_1 _964_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net56),
    .S1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_168_));
 sky130_fd_sc_hd__mux4_1 _965_ (.A0(_166_),
    .A1(_168_),
    .A2(_165_),
    .A3(_167_),
    .S0(net15),
    .S1(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_169_));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net131));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net132));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net133));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net134));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net135));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net136));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net137));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 fanout7 (.A(_000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(_000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 fanout27 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout40 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout41 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout59 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout61 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout63 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__buf_1 fanout67 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout70 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__buf_2 fanout71 (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_1 fanout73 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout75 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_1 fanout77 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_1 fanout80 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__buf_1 fanout82 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_1 fanout86 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout88 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout94 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout95 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout97 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout100 (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__buf_2 fanout103 (.A(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 fanout104 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout122 (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__buf_1 fanout123 (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__buf_2 fanout124 (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__buf_2 fanout129 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net130));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_98 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_3_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_68 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_162 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_6_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_7_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_218 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_230 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_275 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_196 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_9_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_267 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_168 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_274 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_318 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_130 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_13_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_229 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_128 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_14_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_272 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_246 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_46 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_167 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_16_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_83 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_17_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_17_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_244 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_17_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_50 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_18_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_19_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_248 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_168 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_304 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_22_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_111 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_168 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_207 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_219 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_22_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_174 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_186 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_198 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_210 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_23_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_23_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_268 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_24_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_25_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_56 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_227 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_26_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_134 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_27_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_247 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_27_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_28_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_28_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_29_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_191 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_29_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_162 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_30_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_30_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_30_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_31_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_32_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_31 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_62 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_134 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_196 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_256 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_34_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_68 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_34_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_106 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_34_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_160 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_172 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_34_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_211 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_117 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_35_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_33 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_77 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_16 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_38_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net130;
 assign uio_oe[1] = net131;
 assign uio_oe[2] = net132;
 assign uio_oe[3] = net133;
 assign uio_oe[4] = net134;
 assign uio_oe[5] = net135;
 assign uio_oe[6] = net136;
 assign uio_oe[7] = net137;
endmodule
