module tt_um_SNPU (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[32].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[33].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ;
 wire \rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;

 sky130_fd_sc_hd__inv_2 _0342_ (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0343_ (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0344_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2b_1 _0345_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0346_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0347_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0348_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0349_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0350_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0351_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0352_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0353_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0354_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0355_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0356_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0357_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0358_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0359_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0360_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0361_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0362_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0363_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0364_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0365_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0366_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0367_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0368_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0369_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0370_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0371_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0372_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0373_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0374_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0375_ (.A_N(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0376_ (.A_N(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0377_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0378_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0379_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0380_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0381_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0382_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0383_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0384_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0385_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0386_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0387_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0388_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0389_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0390_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0391_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0392_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0393_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0394_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0395_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0396_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0397_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0398_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0399_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0400_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0401_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0402_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0403_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0404_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0405_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0406_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0407_ (.A_N(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0408_ (.A_N(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0409_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0410_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0411_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0412_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0413_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0414_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0415_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0416_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0417_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0418_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0419_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0420_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0421_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0422_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0423_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0424_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0425_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0426_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0427_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0428_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0429_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0430_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0431_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0432_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0433_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0434_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0435_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0436_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0437_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0438_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0439_ (.A_N(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0440_ (.A_N(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0441_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0442_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0443_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0444_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0445_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0446_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0447_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0448_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0449_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0450_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0451_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0452_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0453_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0454_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0455_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0456_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0457_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0458_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0459_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0460_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0461_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0462_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0463_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0464_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0465_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0466_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0467_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0468_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0469_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0470_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0471_ (.A_N(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0472_ (.A_N(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0473_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0474_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0475_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0476_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0477_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0478_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0479_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0480_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0481_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0482_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0483_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0484_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0485_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0486_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0487_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0488_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0489_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0490_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0491_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0492_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0493_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0494_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0495_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0496_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0497_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0498_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0499_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0500_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0501_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0502_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0503_ (.A_N(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0504_ (.A_N(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0505_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0506_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0507_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0508_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0509_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0510_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0511_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0512_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0513_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0514_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0515_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0516_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0517_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0518_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0519_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0520_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0521_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0522_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0523_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0524_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0525_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0526_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0527_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0528_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0529_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0530_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0531_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0532_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0533_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0534_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0535_ (.A_N(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0536_ (.A_N(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0537_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0538_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0539_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0540_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0541_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0542_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0543_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0544_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0545_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0546_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0547_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0548_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0549_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0550_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0551_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0552_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0553_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0554_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0555_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0556_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0557_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0558_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0559_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0560_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0561_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0562_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0563_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0564_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0565_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0566_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0567_ (.A_N(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0568_ (.A_N(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0569_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0570_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0571_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0572_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0573_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0574_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0575_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0576_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0577_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0578_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0579_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0580_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0581_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0582_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0583_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0584_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0585_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0586_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0587_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0588_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0589_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0590_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0591_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0592_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0593_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0594_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0595_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0596_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0597_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0598_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0599_ (.A_N(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0600_ (.A_N(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0601_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0602_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0603_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0604_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0605_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0606_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0607_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0608_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0609_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0610_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0611_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0612_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0613_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0614_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0615_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0616_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0617_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0618_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0619_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0620_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0621_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0622_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0623_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0624_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0625_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0626_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0627_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0628_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0629_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0630_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0631_ (.A_N(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0632_ (.A_N(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0633_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0634_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0635_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0636_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0637_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0638_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0639_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0640_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0641_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0642_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0643_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0644_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0645_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0646_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0647_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0648_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0649_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0650_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0651_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0652_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0653_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0654_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0655_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0656_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0657_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0658_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0659_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0660_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0661_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0662_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0663_ (.A_N(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0664_ (.A_N(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0665_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0666_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0667_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0668_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0669_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0670_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0671_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0672_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0673_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0674_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0675_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0676_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0677_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0678_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0679_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0680_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0681_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0682_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0683_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0684_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0685_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0686_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0687_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0688_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0689_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0690_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0691_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0692_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0693_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0694_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0695_ (.A_N(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0696_ (.A_N(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0697_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0698_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0699_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0700_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0701_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0702_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0703_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0704_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0705_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0706_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0707_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0708_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0709_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0710_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0711_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0712_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0713_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0714_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0715_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0716_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0717_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0718_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0719_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0720_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0721_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0722_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0723_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0724_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0725_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0726_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0727_ (.A_N(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0728_ (.A_N(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0729_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0730_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0731_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0732_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0733_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0734_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0735_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0736_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0737_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0738_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0739_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0740_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0741_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0742_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0743_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0744_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0745_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0746_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0747_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0748_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0749_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0750_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0751_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0752_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0753_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0754_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0755_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0756_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0757_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0758_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0759_ (.A_N(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0760_ (.A_N(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0761_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0762_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0763_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0764_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0765_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0766_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0767_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0768_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0769_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0770_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0771_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0772_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0773_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0774_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0775_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0776_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0777_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0778_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0779_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0780_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0781_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0782_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0783_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0784_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0785_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0786_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0787_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0788_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0789_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0790_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0791_ (.A_N(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0792_ (.A_N(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0793_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0794_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0795_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0796_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0797_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0798_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0799_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0800_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0801_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0802_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0803_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0804_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0805_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0806_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0807_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0808_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0809_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0810_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0811_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0812_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0813_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0814_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0815_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0816_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0817_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0818_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0819_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0820_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0821_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0822_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0823_ (.A_N(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0824_ (.A_N(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0825_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0826_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0827_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0828_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0829_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0830_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0831_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0832_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0833_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0834_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0835_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0836_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0837_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0838_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0839_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0840_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0841_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0842_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0843_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0844_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0845_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0846_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0847_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0848_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0849_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0850_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0851_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0852_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0853_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0854_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0855_ (.A_N(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0856_ (.A_N(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0857_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0858_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[0].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0859_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0860_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[1].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0861_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0862_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[2].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0863_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0864_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[3].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0865_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0866_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[4].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0867_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0868_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[5].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0869_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0870_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[6].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0871_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0872_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[7].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0873_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0874_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .B(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[8].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0875_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0876_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .B(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[9].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0877_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0878_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[10].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0879_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0880_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[11].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0881_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0882_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[12].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0883_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0884_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[13].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0885_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0886_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[14].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0887_ (.A_N(\rnd_blocks[32].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[32].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nand2b_1 _0888_ (.A_N(\rnd_blocks[33].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\rnd_blocks[33].rnd_bank.rnd_gen[15].rnd_inst.R ));
 sky130_fd_sc_hd__nor3_2 _0889_ (.A(net49),
    .B(net39),
    .C(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0003_));
 sky130_fd_sc_hd__and3_1 _0890_ (.A(net30),
    .B(net7),
    .C(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0891_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__mux4_1 _0892_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(net25),
    .B(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _0894_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__o211a_1 _0895_ (.A1(net37),
    .A2(_0008_),
    .B1(_0007_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__nor3b_1 _0897_ (.A(net39),
    .B(net35),
    .C_N(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0011_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__a221o_1 _0899_ (.A1(net19),
    .A2(_0010_),
    .B1(net14),
    .B2(_0012_),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__nor2_2 _0900_ (.A(net27),
    .B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0014_));
 sky130_fd_sc_hd__mux4_1 _0901_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__a211o_1 _0902_ (.A1(net8),
    .A2(_0015_),
    .B1(_0009_),
    .C1(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_1 _0903_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _0904_ (.A(net37),
    .B(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_1 _0905_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__o211a_1 _0906_ (.A1(net25),
    .A2(_0019_),
    .B1(_0018_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _0907_ (.A1(\rnd_blocks[17].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(net19),
    .B1(net14),
    .B2(\rnd_blocks[19].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(\rnd_blocks[16].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(net19),
    .B1(net14),
    .B2(\rnd_blocks[18].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0909_ (.A0(_0022_),
    .A1(_0021_),
    .S(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _0910_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[0].rnd_inst.R ),
    .S0(net58),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__a21o_1 _0911_ (.A1(net8),
    .A2(_0024_),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__or3_1 _0912_ (.A(_0020_),
    .B(_0023_),
    .C(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__a32o_4 _0913_ (.A1(net23),
    .A2(_0016_),
    .A3(_0026_),
    .B1(net12),
    .B2(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__mux4_1 _0915_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net57),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__or2_1 _0916_ (.A(net37),
    .B(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_1 _0917_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net57),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _0918_ (.A(net25),
    .B(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__mux4_1 _0919_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net66),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0921_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__a221o_1 _0922_ (.A1(net16),
    .A2(_0033_),
    .B1(_0034_),
    .B2(net20),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__a21o_1 _0923_ (.A1(net10),
    .A2(_0032_),
    .B1(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__a31o_1 _0924_ (.A1(net33),
    .A2(_0029_),
    .A3(_0031_),
    .B1(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__mux4_1 _0925_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net57),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _0926_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net57),
    .S1(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _0927_ (.A(net37),
    .B(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__o211a_1 _0928_ (.A1(net25),
    .A2(_0038_),
    .B1(_0040_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _0929_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S0(net59),
    .S1(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _0930_ (.A(net8),
    .B(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[1].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__a221o_1 _0933_ (.A1(net19),
    .A2(_0044_),
    .B1(_0045_),
    .B2(net14),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__or3_1 _0934_ (.A(_0041_),
    .B(_0043_),
    .C(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__a32o_4 _0935_ (.A1(net23),
    .A2(_0037_),
    .A3(_0047_),
    .B1(net12),
    .B2(_0027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _0937_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net62),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__or2_1 _0938_ (.A(net37),
    .B(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__mux4_1 _0939_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net62),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__o211a_1 _0940_ (.A1(net26),
    .A2(_0051_),
    .B1(_0050_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _0941_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net62),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _0942_ (.A(net9),
    .B(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__a221o_1 _0945_ (.A1(net20),
    .A2(_0055_),
    .B1(_0056_),
    .B2(net15),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__or3_1 _0946_ (.A(_0052_),
    .B(_0054_),
    .C(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _0947_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net63),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__or2_1 _0948_ (.A(net26),
    .B(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _0949_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net63),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _0950_ (.A(net38),
    .B(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _0951_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S0(net63),
    .S1(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[2].rnd_inst.R ),
    .S(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__a221o_1 _0954_ (.A1(net15),
    .A2(_0064_),
    .B1(_0065_),
    .B2(net20),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__a21o_1 _0955_ (.A1(net9),
    .A2(_0063_),
    .B1(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__a31o_1 _0956_ (.A1(net34),
    .A2(_0060_),
    .A3(_0062_),
    .B1(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__a32o_4 _0957_ (.A1(net23),
    .A2(_0058_),
    .A3(_0068_),
    .B1(net12),
    .B2(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__mux4_1 _0959_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net56),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0070_));
 sky130_fd_sc_hd__mux4_1 _0960_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net56),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _0961_ (.A(net37),
    .B(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__o211a_1 _0962_ (.A1(net25),
    .A2(_0070_),
    .B1(_0072_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__a221o_1 _0965_ (.A1(net19),
    .A2(_0074_),
    .B1(_0075_),
    .B2(net14),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__mux4_1 _0966_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net56),
    .S1(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__a211o_1 _0967_ (.A1(net8),
    .A2(_0077_),
    .B1(_0076_),
    .C1(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__mux4_1 _0968_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(net26),
    .B(_0079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__mux4_1 _0970_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__o211a_1 _0971_ (.A1(net38),
    .A2(_0081_),
    .B1(_0080_),
    .C1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__mux4_1 _0972_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _0973_ (.A(net9),
    .B(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[3].rnd_inst.R ),
    .S(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__a221o_1 _0976_ (.A1(net20),
    .A2(_0085_),
    .B1(_0086_),
    .B2(net15),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__or3_1 _0977_ (.A(_0082_),
    .B(_0084_),
    .C(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__a32o_4 _0978_ (.A1(net23),
    .A2(_0078_),
    .A3(_0088_),
    .B1(net12),
    .B2(_0069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__mux4_1 _0980_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net56),
    .S1(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0981_ (.A(net37),
    .B(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__mux4_1 _0982_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net56),
    .S1(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0983_ (.A(net25),
    .B(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _0984_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net57),
    .S1(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0987_ (.A1(net14),
    .A2(_0095_),
    .B1(_0096_),
    .B2(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__a211o_1 _0988_ (.A1(net8),
    .A2(_0094_),
    .B1(_0097_),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__a31o_1 _0989_ (.A1(net33),
    .A2(_0091_),
    .A3(_0093_),
    .B1(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__mux4_1 _0990_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net59),
    .S1(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__mux4_1 _0991_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net55),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__or2_1 _0992_ (.A(net37),
    .B(_0101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__o211a_1 _0993_ (.A1(net25),
    .A2(_0100_),
    .B1(_0102_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__mux4_1 _0994_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S0(net59),
    .S1(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__and2_1 _0995_ (.A(net8),
    .B(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[4].rnd_inst.R ),
    .S(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__a221o_1 _0998_ (.A1(net19),
    .A2(_0106_),
    .B1(_0107_),
    .B2(net14),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__or3_1 _0999_ (.A(_0103_),
    .B(_0105_),
    .C(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__a32o_4 _1000_ (.A1(net23),
    .A2(_0099_),
    .A3(_0109_),
    .B1(net12),
    .B2(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__mux4_1 _1002_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net60),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(net38),
    .B(_0111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_1 _1004_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net60),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__o211a_1 _1005_ (.A1(net26),
    .A2(_0113_),
    .B1(_0112_),
    .C1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _1006_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net60),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _1007_ (.A(net9),
    .B(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0118_));
 sky130_fd_sc_hd__a221o_1 _1010_ (.A1(net20),
    .A2(_0117_),
    .B1(_0118_),
    .B2(net15),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0119_));
 sky130_fd_sc_hd__or3_1 _1011_ (.A(_0114_),
    .B(_0116_),
    .C(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0120_));
 sky130_fd_sc_hd__mux4_1 _1012_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__mux4_1 _1013_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__or2_1 _1014_ (.A(net38),
    .B(_0122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0123_));
 sky130_fd_sc_hd__o211a_1 _1015_ (.A1(net25),
    .A2(_0121_),
    .B1(_0123_),
    .C1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__mux4_1 _1016_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S0(net62),
    .S1(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _1017_ (.A(net9),
    .B(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[5].rnd_inst.R ),
    .S(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__a221o_1 _1020_ (.A1(net20),
    .A2(_0127_),
    .B1(_0128_),
    .B2(net15),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__or3_1 _1021_ (.A(_0124_),
    .B(_0126_),
    .C(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__a32o_4 _1022_ (.A1(net23),
    .A2(_0120_),
    .A3(_0130_),
    .B1(net12),
    .B2(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__mux4_1 _1024_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_1 _1025_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net61),
    .S1(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _1026_ (.A(net38),
    .B(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__o211a_1 _1027_ (.A1(net26),
    .A2(_0132_),
    .B1(_0134_),
    .C1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__mux4_1 _1028_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net60),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _1029_ (.A(net9),
    .B(_0136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__a221o_1 _1032_ (.A1(net20),
    .A2(_0138_),
    .B1(_0139_),
    .B2(net15),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__or3_1 _1033_ (.A(_0135_),
    .B(_0137_),
    .C(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__mux4_1 _1034_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net60),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__mux4_1 _1035_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net60),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _1036_ (.A(net38),
    .B(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__o211a_1 _1037_ (.A1(net26),
    .A2(_0142_),
    .B1(_0144_),
    .C1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1038_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__mux4_1 _1040_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[6].rnd_inst.R ),
    .S0(net64),
    .S1(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _1041_ (.A(net9),
    .B(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__a221o_1 _1042_ (.A1(net15),
    .A2(_0146_),
    .B1(_0147_),
    .B2(net20),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__or3_1 _1043_ (.A(_0145_),
    .B(_0149_),
    .C(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__a32o_4 _1044_ (.A1(net23),
    .A2(_0141_),
    .A3(_0151_),
    .B1(net12),
    .B2(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__mux2_1 _1045_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__mux4_1 _1046_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net55),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__mux4_1 _1047_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net55),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _1048_ (.A(net37),
    .B(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__o211a_1 _1049_ (.A1(net25),
    .A2(_0153_),
    .B1(_0155_),
    .C1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1051_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__a221o_1 _1052_ (.A1(net19),
    .A2(_0157_),
    .B1(_0158_),
    .B2(net14),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__mux4_1 _1053_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net55),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__a211o_1 _1054_ (.A1(net8),
    .A2(_0160_),
    .B1(_0159_),
    .C1(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _1055_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__and2b_1 _1056_ (.A_N(net41),
    .B(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1057_ (.A0(\rnd_blocks[30].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[31].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__a211o_1 _1058_ (.A1(net41),
    .A2(_0164_),
    .B1(_0163_),
    .C1(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__mux4_1 _1059_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net55),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__or2_1 _1060_ (.A(net37),
    .B(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__mux4_1 _1061_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S0(net56),
    .S1(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _1063_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[7].rnd_inst.R ),
    .S(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__a221o_1 _1064_ (.A1(net19),
    .A2(_0169_),
    .B1(_0170_),
    .B2(net14),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__a21o_1 _1065_ (.A1(net8),
    .A2(_0168_),
    .B1(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__a31o_1 _1066_ (.A1(net33),
    .A2(_0165_),
    .A3(_0167_),
    .B1(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__a32o_4 _1067_ (.A1(net23),
    .A2(_0161_),
    .A3(_0173_),
    .B1(net12),
    .B2(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__mux2_1 _1068_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__mux4_1 _1069_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _1070_ (.A(net28),
    .B(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__mux4_1 _1071_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__or2_1 _1072_ (.A(net40),
    .B(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__mux4_1 _1073_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1074_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _1075_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__a221o_1 _1076_ (.A1(net21),
    .A2(_0180_),
    .B1(_0181_),
    .B2(net16),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__a21o_1 _1077_ (.A1(net10),
    .A2(_0179_),
    .B1(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__a31o_1 _1078_ (.A1(net36),
    .A2(_0176_),
    .A3(_0178_),
    .B1(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__mux4_1 _1079_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__mux4_1 _1080_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _1081_ (.A(net40),
    .B(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__o211a_1 _1082_ (.A1(net28),
    .A2(_0185_),
    .B1(_0187_),
    .C1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _1083_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S0(net74),
    .S1(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _1084_ (.A(net10),
    .B(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _1085_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[8].rnd_inst.R ),
    .S(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__a221o_1 _1087_ (.A1(net22),
    .A2(_0191_),
    .B1(_0192_),
    .B2(net17),
    .C1(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__or3_1 _1088_ (.A(_0188_),
    .B(_0190_),
    .C(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__a32o_4 _1089_ (.A1(net23),
    .A2(_0184_),
    .A3(_0194_),
    .B1(net12),
    .B2(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__mux4_1 _1091_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net72),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _1092_ (.A(net28),
    .B(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__mux4_1 _1093_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net72),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(net40),
    .B(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__mux4_1 _1095_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net72),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _1097_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__a221o_1 _1098_ (.A1(net21),
    .A2(_0201_),
    .B1(_0202_),
    .B2(net17),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__a21o_1 _1099_ (.A1(net11),
    .A2(_0200_),
    .B1(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__a31o_1 _1100_ (.A1(net36),
    .A2(_0197_),
    .A3(_0199_),
    .B1(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__mux4_1 _1101_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net63),
    .S1(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(net28),
    .B(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__mux4_1 _1103_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net72),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__o211a_1 _1104_ (.A1(net40),
    .A2(_0208_),
    .B1(_0207_),
    .C1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__mux4_1 _1105_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S0(net76),
    .S1(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__and2_1 _1106_ (.A(net8),
    .B(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1107_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[9].rnd_inst.R ),
    .S(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__a221o_1 _1109_ (.A1(net20),
    .A2(_0212_),
    .B1(_0213_),
    .B2(net15),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__or3_1 _1110_ (.A(_0209_),
    .B(_0211_),
    .C(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__a32o_4 _1111_ (.A1(net24),
    .A2(_0205_),
    .A3(_0215_),
    .B1(net13),
    .B2(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__mux4_1 _1113_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__or2_1 _1114_ (.A(net39),
    .B(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__mux4_1 _1115_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__or2_1 _1116_ (.A(net27),
    .B(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__mux4_1 _1117_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__a221o_1 _1120_ (.A1(net21),
    .A2(_0222_),
    .B1(_0223_),
    .B2(net16),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__a32o_1 _1121_ (.A1(net35),
    .A2(_0218_),
    .A3(_0220_),
    .B1(_0221_),
    .B2(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__or2_1 _1122_ (.A(_0224_),
    .B(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__and2b_1 _1124_ (.A_N(net50),
    .B(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1125_ (.A0(\rnd_blocks[30].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[31].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_1 _1126_ (.A1(net50),
    .A2(_0229_),
    .B1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__mux4_1 _1127_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net68),
    .S1(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__o221a_1 _1128_ (.A1(_0228_),
    .A2(_0230_),
    .B1(_0231_),
    .B2(net39),
    .C1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__mux4_1 _1129_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S0(net68),
    .S1(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1130_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[10].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__a221o_1 _1132_ (.A1(net16),
    .A2(_0234_),
    .B1(_0235_),
    .B2(net21),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__a211o_1 _1133_ (.A1(net10),
    .A2(_0233_),
    .B1(_0236_),
    .C1(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__a32o_4 _1134_ (.A1(net24),
    .A2(_0226_),
    .A3(_0237_),
    .B1(net13),
    .B2(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__mux4_1 _1136_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net73),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(net28),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__mux4_1 _1138_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net74),
    .S1(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(net40),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__mux4_1 _1140_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net75),
    .S1(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _1141_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1142_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__a221o_1 _1143_ (.A1(net22),
    .A2(_0244_),
    .B1(_0245_),
    .B2(net17),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__a21o_1 _1144_ (.A1(net11),
    .A2(_0243_),
    .B1(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__a31o_1 _1145_ (.A1(net36),
    .A2(_0240_),
    .A3(_0242_),
    .B1(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__mux4_1 _1146_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net73),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__mux4_1 _1147_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net73),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _1148_ (.A(net40),
    .B(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__o211a_1 _1149_ (.A1(net28),
    .A2(_0249_),
    .B1(_0251_),
    .C1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__mux4_1 _1150_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S0(net73),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__and2_1 _1151_ (.A(net11),
    .B(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[11].rnd_inst.R ),
    .S(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__a221o_1 _1154_ (.A1(net22),
    .A2(_0255_),
    .B1(_0256_),
    .B2(net17),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__or3_1 _1155_ (.A(_0252_),
    .B(_0254_),
    .C(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__a32o_4 _1156_ (.A1(net24),
    .A2(_0248_),
    .A3(_0258_),
    .B1(net13),
    .B2(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__mux4_1 _1158_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _1159_ (.A(net27),
    .B(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__mux4_1 _1160_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _1161_ (.A(net40),
    .B(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__mux4_1 _1162_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _1165_ (.A1(net17),
    .A2(_0265_),
    .B1(_0266_),
    .B2(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__a211o_1 _1166_ (.A1(net11),
    .A2(_0264_),
    .B1(_0267_),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__a31o_1 _1167_ (.A1(net36),
    .A2(_0261_),
    .A3(_0263_),
    .B1(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__mux4_1 _1168_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__mux4_1 _1169_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _1170_ (.A(net40),
    .B(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__o211a_1 _1171_ (.A1(net28),
    .A2(_0270_),
    .B1(_0272_),
    .C1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__mux4_1 _1172_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S0(net71),
    .S1(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__and2_1 _1173_ (.A(net11),
    .B(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[12].rnd_inst.R ),
    .S(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__a221o_1 _1176_ (.A1(net22),
    .A2(_0276_),
    .B1(_0277_),
    .B2(net16),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _1177_ (.A(_0273_),
    .B(_0275_),
    .C(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__a32o_4 _1178_ (.A1(net24),
    .A2(_0269_),
    .A3(_0279_),
    .B1(net13),
    .B2(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__mux2_1 _1179_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__mux4_1 _1180_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net75),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_1 _1181_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net68),
    .S1(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _1182_ (.A(net39),
    .B(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__o211a_1 _1183_ (.A1(net27),
    .A2(_0281_),
    .B1(_0283_),
    .C1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__a221o_1 _1186_ (.A1(net21),
    .A2(_0285_),
    .B1(_0286_),
    .B2(net16),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__mux4_1 _1187_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net73),
    .S1(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__a211o_1 _1188_ (.A1(net10),
    .A2(_0288_),
    .B1(_0287_),
    .C1(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__mux4_1 _1189_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net66),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _1190_ (.A(net27),
    .B(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__mux4_1 _1191_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net70),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1192_ (.A(net39),
    .B(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _1193_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__mux4_1 _1194_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S0(net70),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[13].rnd_inst.R ),
    .S(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(net16),
    .A2(_0294_),
    .B1(_0296_),
    .B2(net21),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__a32o_1 _1197_ (.A1(net35),
    .A2(_0291_),
    .A3(_0293_),
    .B1(_0295_),
    .B2(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _1198_ (.A(_0297_),
    .B(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__a32o_4 _1199_ (.A1(net24),
    .A2(_0289_),
    .A3(_0299_),
    .B1(net13),
    .B2(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__mux4_1 _1201_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _1202_ (.A(net27),
    .B(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__mux4_1 _1203_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__or2_1 _1204_ (.A(net39),
    .B(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__mux4_1 _1205_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net69),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1206_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1207_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__a221o_1 _1208_ (.A1(net21),
    .A2(_0306_),
    .B1(_0307_),
    .B2(net16),
    .C1(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__a21o_1 _1209_ (.A1(net10),
    .A2(_0305_),
    .B1(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__a31o_1 _1210_ (.A1(net35),
    .A2(_0302_),
    .A3(_0304_),
    .B1(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__mux4_1 _1211_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__mux4_1 _1212_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net67),
    .S1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__or2_1 _1213_ (.A(net40),
    .B(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__o211a_1 _1214_ (.A1(net27),
    .A2(_0311_),
    .B1(_0313_),
    .C1(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1215_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__mux4_1 _1216_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S0(net70),
    .S1(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1217_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[14].rnd_inst.R ),
    .S(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _1218_ (.A1(net16),
    .A2(_0315_),
    .B1(_0317_),
    .B2(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__a21o_1 _1219_ (.A1(net10),
    .A2(_0316_),
    .B1(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _1220_ (.A(net32),
    .B(_0314_),
    .C(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__a32o_4 _1221_ (.A1(net24),
    .A2(_0310_),
    .A3(_0320_),
    .B1(net13),
    .B2(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(\rnd_blocks[32].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[33].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__mux4_1 _1223_ (.A0(\rnd_blocks[24].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[25].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[26].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[27].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net65),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _1224_ (.A(net39),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__mux4_1 _1225_ (.A0(\rnd_blocks[28].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[29].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[30].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[31].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net65),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _1226_ (.A(net27),
    .B(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(\rnd_blocks[16].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[17].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _1228_ (.A0(\rnd_blocks[18].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[19].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__a221o_1 _1229_ (.A1(net19),
    .A2(_0326_),
    .B1(_0327_),
    .B2(net14),
    .C1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__mux4_1 _1230_ (.A0(\rnd_blocks[20].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[21].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[22].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[23].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net65),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__a32o_1 _1231_ (.A1(net35),
    .A2(_0323_),
    .A3(_0325_),
    .B1(_0329_),
    .B2(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _1232_ (.A(_0328_),
    .B(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__mux4_1 _1233_ (.A0(\rnd_blocks[12].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[13].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[14].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[15].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net65),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _1234_ (.A(net27),
    .B(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__mux4_1 _1235_ (.A0(\rnd_blocks[8].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[9].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[10].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[11].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net65),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _1236_ (.A(net39),
    .B(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__mux4_1 _1237_ (.A0(\rnd_blocks[4].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[5].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A2(\rnd_blocks[6].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A3(\rnd_blocks[7].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S0(net66),
    .S1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1238_ (.A0(\rnd_blocks[0].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[1].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(\rnd_blocks[2].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .A1(\rnd_blocks[3].rnd_bank.rnd_gen[15].rnd_inst.R ),
    .S(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__a221o_1 _1240_ (.A1(net21),
    .A2(_0337_),
    .B1(_0338_),
    .B2(net16),
    .C1(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__a32o_1 _1241_ (.A1(net35),
    .A2(_0333_),
    .A3(_0335_),
    .B1(_0336_),
    .B2(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _1242_ (.A(_0339_),
    .B(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__a32o_4 _1243_ (.A1(net23),
    .A2(_0331_),
    .A3(_0341_),
    .B1(net12),
    .B2(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net151));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net152));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net153));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net154));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net155));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net156));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net157));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout11 (.A(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_8 fanout12 (.A(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 max_cap18 (.A(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout38 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout42 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout44 (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 fanout80 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_1 fanout90 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout92 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout93 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__buf_2 fanout97 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout98 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__buf_2 fanout100 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__buf_1 fanout109 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout112 (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__buf_1 fanout115 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__buf_1 fanout126 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout128 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__buf_1 fanout133 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__buf_1 fanout136 (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__buf_1 fanout138 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout140 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 fanout142 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout147 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__buf_1 fanout148 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__conb_1 tt_um_SNPU_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net150));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_230 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_314 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_2_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_178 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_226 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_274 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_2_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_80 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_3_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_247 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_259 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_227 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_5_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_80 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_62 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_6_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_91 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_6_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_214 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_275 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_6_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_25 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_128 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_152 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_7_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_8_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_9_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_123 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_10_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_88 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_192 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_117 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_12_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_13_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_247 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_15_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_254 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_101 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_16_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_16_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_202 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_16_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_16_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_17_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_17_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_211 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_92 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_104 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_145 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_180 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_21_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_98 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_21_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_228 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_23_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_145 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_23_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_92 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_104 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_116 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_24_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_25_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_25_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_268 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_26_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_26_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_27_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_76 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_27_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_112 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_214 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_226 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_28_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_230 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_108 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_30_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_30_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_199 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_31_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_32_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_32_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_32_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_83 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_196 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_245 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_34_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_102 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_228 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_284 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_34_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_35_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_35_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_142 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_144 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_38_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_38_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_38_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_38_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net150;
 assign uio_oe[1] = net151;
 assign uio_oe[2] = net152;
 assign uio_oe[3] = net153;
 assign uio_oe[4] = net154;
 assign uio_oe[5] = net155;
 assign uio_oe[6] = net156;
 assign uio_oe[7] = net157;
endmodule
