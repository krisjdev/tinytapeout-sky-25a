VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_asic_1
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_asic_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 77.574997 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 180.000000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 50.000000 ;
    ANTENNADIFFAREA 0.290000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.000000 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.000000 ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.000000 ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 947.392456 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 315.000 5.000 317.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER pwell ;
        RECT 15.745 153.590 31.075 214.700 ;
      LAYER nwell ;
        RECT 32.750 154.785 56.960 158.755 ;
      LAYER pwell ;
        RECT 63.685 135.215 93.795 141.140 ;
        RECT 63.435 134.660 93.795 135.215 ;
        RECT 63.685 122.850 93.795 134.660 ;
        RECT 94.690 140.420 114.830 141.185 ;
        RECT 94.690 135.250 95.455 140.420 ;
        RECT 100.625 135.250 102.175 140.420 ;
        RECT 107.345 135.250 108.895 140.420 ;
        RECT 114.065 135.250 114.830 140.420 ;
        RECT 94.690 133.700 114.830 135.250 ;
        RECT 94.690 128.530 95.455 133.700 ;
        RECT 100.625 128.530 102.175 133.700 ;
        RECT 107.345 128.530 108.895 133.700 ;
        RECT 114.065 128.530 114.830 133.700 ;
        RECT 94.690 126.980 114.830 128.530 ;
        RECT 94.690 121.810 95.455 126.980 ;
        RECT 100.625 121.810 102.175 126.980 ;
        RECT 107.345 121.810 108.895 126.980 ;
        RECT 114.065 121.810 114.830 126.980 ;
        RECT 80.650 121.165 81.120 121.480 ;
        RECT 56.055 98.885 81.120 121.165 ;
        RECT 94.690 121.045 114.830 121.810 ;
        RECT 104.660 117.130 126.940 119.130 ;
        RECT 82.380 111.550 126.940 117.130 ;
        RECT 82.415 105.190 126.940 110.770 ;
        RECT 82.415 103.190 104.695 105.190 ;
        RECT 80.650 98.340 81.120 98.885 ;
      LAYER nwell ;
        RECT 57.315 83.515 79.895 96.485 ;
        RECT 67.365 71.495 79.895 75.465 ;
        RECT 82.755 71.495 126.965 96.485 ;
        RECT 129.595 72.065 135.585 94.645 ;
      LAYER pwell ;
        RECT 240.550 84.250 244.130 90.640 ;
        RECT 259.745 89.030 272.565 93.540 ;
        RECT 264.710 87.085 272.530 89.030 ;
        RECT 246.175 85.010 271.995 87.020 ;
      LAYER nwell ;
        RECT 72.245 59.755 77.425 59.905 ;
        RECT 48.670 54.625 61.300 58.440 ;
        RECT 72.190 56.440 77.585 59.755 ;
        RECT 72.245 56.365 77.425 56.440 ;
        RECT 38.670 54.470 61.300 54.625 ;
        RECT 38.670 49.785 61.250 54.470 ;
      LAYER pwell ;
        RECT 69.185 50.290 80.305 53.870 ;
      LAYER nwell ;
        RECT 165.740 51.355 189.545 56.450 ;
        RECT 193.920 51.355 223.950 68.110 ;
        RECT 229.890 62.035 234.860 78.010 ;
        RECT 165.740 51.200 223.950 51.355 ;
        RECT 164.450 51.185 223.950 51.200 ;
        RECT 38.670 49.655 63.200 49.785 ;
        RECT 39.230 39.015 48.890 49.655 ;
        RECT 53.560 38.890 63.200 49.655 ;
      LAYER pwell ;
        RECT 35.780 24.305 52.340 38.625 ;
        RECT 53.710 35.045 58.190 38.625 ;
        RECT 58.570 35.050 63.050 38.630 ;
        RECT 91.745 30.570 104.325 49.940 ;
        RECT 109.450 41.175 129.270 47.625 ;
        RECT 104.680 30.550 116.960 39.990 ;
        RECT 116.990 30.550 129.270 39.990 ;
        RECT 87.160 18.090 129.270 30.460 ;
        RECT 146.080 28.240 158.660 50.720 ;
      LAYER nwell ;
        RECT 161.370 44.715 223.950 51.185 ;
        RECT 161.355 43.605 223.950 44.715 ;
        RECT 161.350 43.480 223.950 43.605 ;
        RECT 161.350 42.640 178.345 43.480 ;
        RECT 189.415 43.385 223.950 43.480 ;
        RECT 165.735 32.095 178.345 42.640 ;
        RECT 181.185 34.370 186.055 41.340 ;
        RECT 193.920 40.280 223.950 43.385 ;
        RECT 229.885 61.650 234.860 62.035 ;
      LAYER pwell ;
        RECT 240.550 77.775 253.130 84.250 ;
        RECT 240.550 65.080 244.130 77.775 ;
      LAYER nwell ;
        RECT 193.920 39.465 224.225 40.280 ;
        RECT 189.690 35.495 224.225 39.465 ;
      LAYER pwell ;
        RECT 145.760 18.525 160.650 26.105 ;
        RECT 161.500 18.950 174.080 30.230 ;
      LAYER nwell ;
        RECT 193.920 19.385 224.225 35.495 ;
        RECT 229.885 20.120 234.855 61.650 ;
      LAYER pwell ;
        RECT 240.550 26.655 246.130 65.080 ;
        RECT 240.550 23.550 244.130 26.655 ;
        RECT 240.550 23.460 244.145 23.550 ;
        RECT 240.565 20.270 244.145 23.460 ;
        RECT 256.620 20.030 261.590 81.040 ;
      LAYER nwell ;
        RECT 209.035 19.310 224.225 19.385 ;
      LAYER li1 ;
        RECT 14.670 215.780 31.615 215.790 ;
        RECT 14.670 214.235 31.850 215.780 ;
        RECT 14.670 184.230 16.225 214.235 ;
        RECT 16.575 211.710 16.925 213.870 ;
        RECT 16.575 184.710 16.925 186.870 ;
        RECT 17.405 184.230 17.575 214.235 ;
        RECT 18.055 211.710 18.405 213.870 ;
        RECT 18.055 184.710 18.405 186.870 ;
        RECT 18.885 184.230 19.055 214.235 ;
        RECT 19.535 211.710 19.885 213.870 ;
        RECT 19.535 184.710 19.885 186.870 ;
        RECT 20.365 184.230 20.535 214.235 ;
        RECT 21.015 211.710 21.365 213.870 ;
        RECT 21.015 184.710 21.365 186.870 ;
        RECT 21.845 184.230 22.015 214.235 ;
        RECT 22.495 211.710 22.845 213.870 ;
        RECT 22.495 184.710 22.845 186.870 ;
        RECT 23.325 184.230 23.495 214.235 ;
        RECT 23.975 211.710 24.325 213.870 ;
        RECT 23.975 184.710 24.325 186.870 ;
        RECT 24.805 184.230 24.975 214.235 ;
        RECT 25.455 211.710 25.805 213.870 ;
        RECT 25.455 184.710 25.805 186.870 ;
        RECT 26.285 184.230 26.455 214.235 ;
        RECT 26.935 211.710 27.285 213.870 ;
        RECT 26.935 184.710 27.285 186.870 ;
        RECT 27.765 184.230 27.935 214.235 ;
        RECT 28.415 211.710 28.765 213.870 ;
        RECT 28.415 184.710 28.765 186.870 ;
        RECT 29.245 184.230 29.415 214.235 ;
        RECT 29.895 211.710 30.245 213.870 ;
        RECT 29.895 184.710 30.245 186.870 ;
        RECT 30.595 184.230 31.850 214.235 ;
        RECT 14.670 184.060 31.850 184.230 ;
        RECT 14.670 154.150 16.225 184.060 ;
        RECT 16.575 181.420 16.925 183.580 ;
        RECT 16.575 154.420 16.925 156.580 ;
        RECT 17.405 154.150 17.575 184.060 ;
        RECT 18.055 181.420 18.405 183.580 ;
        RECT 18.055 154.420 18.405 156.580 ;
        RECT 18.885 154.150 19.055 184.060 ;
        RECT 19.535 181.420 19.885 183.580 ;
        RECT 19.535 154.420 19.885 156.580 ;
        RECT 20.365 154.150 20.535 184.060 ;
        RECT 21.015 181.420 21.365 183.580 ;
        RECT 21.015 154.420 21.365 156.580 ;
        RECT 21.845 154.150 22.015 184.060 ;
        RECT 22.495 181.420 22.845 183.580 ;
        RECT 22.495 154.420 22.845 156.580 ;
        RECT 23.325 154.150 23.495 184.060 ;
        RECT 23.975 181.420 24.325 183.580 ;
        RECT 23.975 154.420 24.325 156.580 ;
        RECT 24.805 154.150 24.975 184.060 ;
        RECT 25.455 181.420 25.805 183.580 ;
        RECT 25.455 154.420 25.805 156.580 ;
        RECT 26.285 154.150 26.455 184.060 ;
        RECT 26.935 181.420 27.285 183.580 ;
        RECT 26.935 154.420 27.285 156.580 ;
        RECT 27.765 154.150 27.935 184.060 ;
        RECT 28.415 181.420 28.765 183.580 ;
        RECT 28.415 154.420 28.765 156.580 ;
        RECT 29.245 154.150 29.415 184.060 ;
        RECT 29.895 181.420 30.245 183.580 ;
        RECT 29.895 154.420 30.245 156.580 ;
        RECT 30.595 154.150 31.850 184.060 ;
        RECT 32.805 159.100 57.060 159.195 ;
        RECT 32.755 158.170 57.165 159.100 ;
        RECT 32.755 155.415 33.445 158.170 ;
        RECT 34.040 157.505 44.040 157.675 ;
        RECT 33.810 156.250 33.980 157.290 ;
        RECT 44.100 156.250 44.270 157.290 ;
        RECT 34.040 155.865 44.040 156.035 ;
        RECT 44.770 155.415 44.940 158.170 ;
        RECT 45.670 157.505 55.670 157.675 ;
        RECT 45.440 156.250 45.610 157.290 ;
        RECT 55.730 156.250 55.900 157.290 ;
        RECT 45.670 155.865 55.670 156.035 ;
        RECT 56.385 155.415 57.165 158.170 ;
        RECT 32.755 154.355 57.165 155.415 ;
        RECT 14.670 152.820 31.850 154.150 ;
        RECT 63.260 140.660 114.750 141.530 ;
        RECT 63.260 139.615 64.060 140.660 ;
        RECT 64.515 139.960 66.675 140.310 ;
        RECT 76.015 139.960 78.175 140.310 ;
        RECT 78.470 139.615 78.960 140.660 ;
        RECT 79.305 139.960 81.465 140.310 ;
        RECT 90.805 139.960 92.965 140.310 ;
        RECT 93.435 139.880 114.750 140.660 ;
        RECT 93.435 139.615 95.995 139.880 ;
        RECT 63.260 139.060 95.995 139.615 ;
        RECT 63.260 138.150 64.060 139.060 ;
        RECT 64.515 138.480 66.675 138.830 ;
        RECT 76.015 138.480 78.175 138.830 ;
        RECT 78.470 138.150 78.960 139.060 ;
        RECT 79.305 138.480 81.465 138.830 ;
        RECT 90.805 138.480 92.965 138.830 ;
        RECT 93.435 138.150 95.995 139.060 ;
        RECT 63.260 137.595 95.995 138.150 ;
        RECT 63.260 136.680 64.060 137.595 ;
        RECT 64.515 137.000 66.675 137.350 ;
        RECT 76.015 137.000 78.175 137.350 ;
        RECT 78.470 136.680 78.960 137.595 ;
        RECT 79.305 137.000 81.465 137.350 ;
        RECT 90.805 137.000 92.965 137.350 ;
        RECT 93.435 136.680 95.995 137.595 ;
        RECT 63.260 136.125 95.995 136.680 ;
        RECT 63.260 135.215 64.060 136.125 ;
        RECT 64.515 135.520 66.675 135.870 ;
        RECT 76.015 135.520 78.175 135.870 ;
        RECT 78.470 135.215 78.960 136.125 ;
        RECT 79.305 135.520 81.465 135.870 ;
        RECT 90.805 135.520 92.965 135.870 ;
        RECT 93.435 135.790 95.995 136.125 ;
        RECT 96.305 136.100 99.775 139.570 ;
        RECT 100.085 135.790 102.715 139.880 ;
        RECT 103.025 136.100 106.495 139.570 ;
        RECT 106.805 135.790 109.435 139.880 ;
        RECT 109.745 136.100 113.215 139.570 ;
        RECT 113.525 135.790 114.750 139.880 ;
        RECT 93.435 135.215 114.750 135.790 ;
        RECT 63.260 134.660 114.750 135.215 ;
        RECT 63.260 133.750 64.060 134.660 ;
        RECT 64.515 134.040 66.675 134.390 ;
        RECT 76.015 134.040 78.175 134.390 ;
        RECT 78.470 133.750 78.960 134.660 ;
        RECT 79.305 134.040 81.465 134.390 ;
        RECT 90.805 134.040 92.965 134.390 ;
        RECT 93.435 133.840 114.750 134.660 ;
        RECT 93.435 133.750 95.855 133.840 ;
        RECT 63.260 133.520 95.855 133.750 ;
        RECT 100.170 133.520 102.585 133.840 ;
        RECT 106.950 133.520 109.250 133.840 ;
        RECT 113.665 133.520 114.750 133.840 ;
        RECT 63.260 133.195 114.750 133.520 ;
        RECT 63.260 132.285 64.060 133.195 ;
        RECT 64.515 132.560 66.675 132.910 ;
        RECT 76.015 132.560 78.175 132.910 ;
        RECT 78.470 132.285 78.960 133.195 ;
        RECT 93.435 133.160 114.750 133.195 ;
        RECT 79.305 132.560 81.465 132.910 ;
        RECT 90.805 132.560 92.965 132.910 ;
        RECT 93.435 132.285 95.995 133.160 ;
        RECT 63.260 131.730 95.995 132.285 ;
        RECT 63.260 130.785 64.060 131.730 ;
        RECT 64.515 131.080 66.675 131.430 ;
        RECT 76.015 131.080 78.175 131.430 ;
        RECT 78.470 130.785 78.960 131.730 ;
        RECT 79.305 131.080 81.465 131.430 ;
        RECT 90.805 131.080 92.965 131.430 ;
        RECT 93.435 130.785 95.995 131.730 ;
        RECT 63.260 130.230 95.995 130.785 ;
        RECT 63.260 129.250 64.060 130.230 ;
        RECT 64.515 129.600 66.675 129.950 ;
        RECT 76.015 129.600 78.175 129.950 ;
        RECT 78.470 129.250 78.960 130.230 ;
        RECT 79.305 129.600 81.465 129.950 ;
        RECT 90.805 129.600 92.965 129.950 ;
        RECT 93.435 129.250 95.995 130.230 ;
        RECT 96.305 129.380 99.775 132.850 ;
        RECT 63.260 129.070 95.995 129.250 ;
        RECT 100.085 129.070 102.715 133.160 ;
        RECT 103.025 129.380 106.495 132.850 ;
        RECT 106.805 129.070 109.435 133.160 ;
        RECT 109.745 129.380 113.215 132.850 ;
        RECT 113.525 129.070 114.750 133.160 ;
        RECT 63.260 128.695 114.750 129.070 ;
        RECT 63.260 127.820 64.060 128.695 ;
        RECT 64.515 128.120 66.675 128.470 ;
        RECT 76.015 128.120 78.175 128.470 ;
        RECT 78.470 127.820 78.960 128.695 ;
        RECT 79.305 128.120 81.465 128.470 ;
        RECT 90.805 128.120 92.965 128.470 ;
        RECT 93.435 127.820 114.750 128.695 ;
        RECT 63.260 127.265 114.750 127.820 ;
        RECT 63.260 126.355 64.060 127.265 ;
        RECT 64.515 126.640 66.675 126.990 ;
        RECT 76.015 126.640 78.175 126.990 ;
        RECT 78.470 126.355 78.960 127.265 ;
        RECT 79.305 126.640 81.465 126.990 ;
        RECT 90.805 126.640 92.965 126.990 ;
        RECT 93.435 126.440 114.750 127.265 ;
        RECT 93.435 126.355 95.995 126.440 ;
        RECT 63.260 125.800 95.995 126.355 ;
        RECT 63.260 124.820 64.060 125.800 ;
        RECT 64.515 125.160 66.675 125.510 ;
        RECT 76.015 125.160 78.175 125.510 ;
        RECT 78.470 124.820 78.960 125.800 ;
        RECT 79.305 125.160 81.465 125.510 ;
        RECT 90.805 125.160 92.965 125.510 ;
        RECT 93.435 124.820 95.995 125.800 ;
        RECT 63.260 124.265 95.995 124.820 ;
        RECT 63.260 123.250 64.060 124.265 ;
        RECT 64.515 123.680 66.675 124.030 ;
        RECT 76.015 123.680 78.175 124.030 ;
        RECT 78.470 123.250 78.960 124.265 ;
        RECT 79.305 123.680 81.465 124.030 ;
        RECT 90.805 123.680 92.965 124.030 ;
        RECT 93.435 123.250 95.995 124.265 ;
        RECT 63.260 123.195 95.995 123.250 ;
        RECT 55.295 122.350 95.995 123.195 ;
        RECT 96.305 122.660 99.775 126.130 ;
        RECT 100.085 122.350 102.715 126.440 ;
        RECT 103.025 122.660 106.495 126.130 ;
        RECT 106.805 122.350 109.435 126.440 ;
        RECT 109.745 122.660 113.215 126.130 ;
        RECT 113.525 122.350 114.750 126.440 ;
        RECT 55.295 120.585 114.750 122.350 ;
        RECT 55.295 99.515 56.490 120.585 ;
        RECT 57.325 120.085 57.865 120.255 ;
        RECT 56.985 100.025 57.155 120.025 ;
        RECT 58.035 100.025 58.205 120.025 ;
        RECT 57.325 99.795 57.865 99.965 ;
        RECT 58.725 99.515 58.895 120.585 ;
        RECT 59.755 120.085 60.295 120.255 ;
        RECT 59.415 100.025 59.585 120.025 ;
        RECT 60.465 100.025 60.635 120.025 ;
        RECT 59.755 99.795 60.295 99.965 ;
        RECT 61.155 99.515 61.325 120.585 ;
        RECT 62.185 120.085 62.725 120.255 ;
        RECT 61.845 100.025 62.015 120.025 ;
        RECT 62.895 100.025 63.065 120.025 ;
        RECT 62.185 99.795 62.725 99.965 ;
        RECT 63.585 99.515 63.755 120.585 ;
        RECT 64.615 120.085 65.155 120.255 ;
        RECT 64.275 100.025 64.445 120.025 ;
        RECT 65.325 100.025 65.495 120.025 ;
        RECT 64.615 99.795 65.155 99.965 ;
        RECT 66.015 99.515 66.185 120.585 ;
        RECT 67.045 120.085 67.585 120.255 ;
        RECT 66.705 100.025 66.875 120.025 ;
        RECT 67.755 100.025 67.925 120.025 ;
        RECT 67.045 99.795 67.585 99.965 ;
        RECT 68.445 99.515 68.615 120.585 ;
        RECT 69.475 120.085 70.015 120.255 ;
        RECT 69.135 100.025 69.305 120.025 ;
        RECT 70.185 100.025 70.355 120.025 ;
        RECT 69.475 99.795 70.015 99.965 ;
        RECT 70.875 99.515 71.045 120.585 ;
        RECT 71.905 120.085 72.445 120.255 ;
        RECT 71.565 100.025 71.735 120.025 ;
        RECT 72.615 100.025 72.785 120.025 ;
        RECT 71.905 99.795 72.445 99.965 ;
        RECT 73.305 99.515 73.475 120.585 ;
        RECT 74.335 120.085 74.875 120.255 ;
        RECT 73.995 100.025 74.165 120.025 ;
        RECT 75.045 100.025 75.215 120.025 ;
        RECT 74.335 99.795 74.875 99.965 ;
        RECT 75.735 99.515 75.905 120.585 ;
        RECT 76.765 120.085 77.305 120.255 ;
        RECT 76.425 100.025 76.595 120.025 ;
        RECT 77.475 100.025 77.645 120.025 ;
        RECT 76.765 99.795 77.305 99.965 ;
        RECT 78.165 99.515 78.335 120.585 ;
        RECT 79.195 120.085 79.735 120.255 ;
        RECT 80.400 120.085 114.750 120.585 ;
        RECT 78.855 100.025 79.025 120.025 ;
        RECT 79.905 100.025 80.075 120.025 ;
        RECT 80.400 118.625 127.360 120.085 ;
        RECT 80.400 116.565 105.165 118.625 ;
        RECT 105.800 118.030 125.800 118.200 ;
        RECT 80.400 112.030 82.845 116.565 ;
        RECT 83.520 116.030 103.520 116.200 ;
        RECT 83.290 112.820 83.460 115.860 ;
        RECT 103.580 112.820 103.750 115.860 ;
        RECT 83.520 112.480 103.520 112.650 ;
        RECT 104.215 112.030 105.165 116.565 ;
        RECT 105.570 112.820 105.740 117.860 ;
        RECT 125.860 112.820 126.030 117.860 ;
        RECT 105.800 112.480 125.800 112.650 ;
        RECT 126.410 112.030 127.360 118.625 ;
        RECT 80.400 110.225 127.360 112.030 ;
        RECT 80.400 103.665 82.890 110.225 ;
        RECT 83.555 109.670 103.555 109.840 ;
        RECT 83.325 104.460 83.495 109.500 ;
        RECT 103.615 104.460 103.785 109.500 ;
        RECT 104.150 105.690 105.135 110.225 ;
        RECT 105.800 109.670 125.800 109.840 ;
        RECT 105.570 106.460 105.740 109.500 ;
        RECT 125.860 106.460 126.030 109.500 ;
        RECT 105.800 106.120 125.800 106.290 ;
        RECT 126.410 105.690 127.360 110.225 ;
        RECT 104.150 105.150 127.360 105.690 ;
        RECT 83.555 104.120 103.555 104.290 ;
        RECT 80.400 103.660 82.900 103.665 ;
        RECT 104.245 103.660 104.585 105.150 ;
        RECT 80.400 103.225 104.600 103.660 ;
        RECT 79.195 99.795 79.735 99.965 ;
        RECT 80.400 99.515 81.055 103.225 ;
        RECT 55.295 98.400 81.055 99.515 ;
        RECT 82.655 96.575 127.125 96.580 ;
        RECT 57.265 95.725 127.125 96.575 ;
        RECT 57.265 95.700 83.405 95.725 ;
        RECT 57.265 89.950 57.930 95.700 ;
        RECT 58.605 95.235 78.605 95.405 ;
        RECT 58.375 93.480 58.545 95.020 ;
        RECT 78.665 93.480 78.835 95.020 ;
        RECT 58.605 93.095 78.605 93.265 ;
        RECT 58.605 92.555 78.605 92.725 ;
        RECT 58.375 90.800 58.545 92.340 ;
        RECT 78.665 90.800 78.835 92.340 ;
        RECT 58.605 90.415 78.605 90.585 ;
        RECT 79.170 89.950 83.405 95.700 ;
        RECT 84.045 95.235 104.045 95.405 ;
        RECT 57.265 88.765 83.405 89.950 ;
        RECT 57.265 84.180 57.930 88.765 ;
        RECT 58.605 88.235 78.605 88.405 ;
        RECT 58.375 84.980 58.545 88.020 ;
        RECT 78.665 84.980 78.835 88.020 ;
        RECT 58.605 84.595 78.605 84.765 ;
        RECT 57.265 84.145 69.330 84.180 ;
        RECT 57.265 84.140 78.520 84.145 ;
        RECT 79.170 84.140 83.405 88.765 ;
        RECT 83.815 84.980 83.985 95.020 ;
        RECT 104.105 84.980 104.275 95.020 ;
        RECT 84.045 84.595 104.045 84.765 ;
        RECT 57.265 84.075 83.405 84.140 ;
        RECT 104.775 84.075 104.945 95.725 ;
        RECT 105.675 95.235 125.675 95.405 ;
        RECT 105.445 84.980 105.615 95.020 ;
        RECT 125.735 84.980 125.905 95.020 ;
        RECT 126.345 94.705 127.095 95.725 ;
        RECT 126.345 93.985 135.740 94.705 ;
        RECT 105.675 84.595 125.675 84.765 ;
        RECT 126.345 84.075 130.270 93.985 ;
        RECT 131.060 93.415 131.600 93.585 ;
        RECT 57.265 83.905 130.270 84.075 ;
        RECT 57.265 83.450 83.405 83.905 ;
        RECT 57.350 83.430 83.405 83.450 ;
        RECT 66.865 74.855 83.405 83.430 ;
        RECT 84.045 83.215 104.045 83.385 ;
        RECT 66.840 74.785 83.405 74.855 ;
        RECT 66.840 72.155 67.930 74.785 ;
        RECT 68.655 74.215 78.605 74.385 ;
        RECT 68.425 72.960 68.595 74.000 ;
        RECT 78.665 72.960 78.835 74.000 ;
        RECT 68.655 72.575 78.605 72.745 ;
        RECT 79.270 72.155 83.405 74.785 ;
        RECT 83.815 72.960 83.985 83.000 ;
        RECT 104.105 72.960 104.275 83.000 ;
        RECT 84.045 72.575 104.045 72.745 ;
        RECT 104.775 72.155 104.945 83.905 ;
        RECT 105.675 83.215 125.675 83.385 ;
        RECT 105.445 72.960 105.615 83.000 ;
        RECT 125.735 72.960 125.905 83.000 ;
        RECT 105.675 72.575 125.675 72.745 ;
        RECT 126.345 72.670 130.270 83.905 ;
        RECT 130.675 73.355 130.845 93.355 ;
        RECT 131.815 73.355 131.985 93.355 ;
        RECT 131.060 73.125 131.600 73.295 ;
        RECT 132.505 72.670 132.675 93.985 ;
        RECT 133.580 93.415 134.120 93.585 ;
        RECT 133.195 73.355 133.365 93.355 ;
        RECT 134.335 73.355 134.505 93.355 ;
        RECT 133.580 73.125 134.120 73.295 ;
        RECT 134.915 72.670 135.740 93.985 ;
        RECT 259.700 92.980 272.575 93.680 ;
        RECT 240.550 90.730 246.630 90.770 ;
        RECT 240.520 90.520 246.630 90.730 ;
        RECT 240.510 90.175 246.630 90.520 ;
        RECT 240.510 87.770 241.085 90.175 ;
        RECT 243.640 90.000 246.630 90.175 ;
        RECT 241.820 89.560 242.860 89.730 ;
        RECT 243.640 89.505 246.635 90.000 ;
        RECT 241.480 88.500 241.650 89.500 ;
        RECT 243.030 88.500 243.200 89.500 ;
        RECT 243.640 88.505 246.630 89.505 ;
        RECT 259.700 89.485 260.150 92.980 ;
        RECT 260.575 89.860 262.735 92.710 ;
        RECT 269.575 89.860 271.735 92.710 ;
        RECT 271.925 89.485 272.575 92.980 ;
        RECT 259.700 88.705 272.575 89.485 ;
        RECT 241.820 88.270 242.860 88.440 ;
        RECT 243.640 88.010 246.635 88.505 ;
        RECT 243.640 87.770 246.630 88.010 ;
        RECT 240.510 87.055 246.630 87.770 ;
        RECT 259.700 87.450 265.140 88.705 ;
        RECT 265.540 87.915 267.700 88.265 ;
        RECT 269.540 87.915 271.700 88.265 ;
        RECT 271.925 87.450 272.575 88.705 ;
        RECT 240.510 87.035 246.635 87.055 ;
        RECT 240.510 84.595 241.085 87.035 ;
        RECT 243.640 86.990 246.635 87.035 ;
        RECT 259.700 86.990 272.575 87.450 ;
        RECT 243.640 86.560 272.575 86.990 ;
        RECT 241.820 86.365 242.860 86.535 ;
        RECT 241.480 85.305 241.650 86.305 ;
        RECT 243.030 85.305 243.200 86.305 ;
        RECT 243.640 85.445 246.630 86.560 ;
        RECT 247.005 85.840 249.165 86.190 ;
        RECT 269.005 85.840 271.165 86.190 ;
        RECT 271.610 85.475 272.575 86.560 ;
        RECT 252.585 85.445 272.575 85.475 ;
        RECT 241.820 85.075 242.860 85.245 ;
        RECT 243.640 84.595 272.575 85.445 ;
        RECT 240.510 83.840 272.575 84.595 ;
        RECT 240.510 81.380 241.085 83.840 ;
        RECT 241.820 83.170 251.860 83.340 ;
        RECT 241.480 82.110 241.650 83.110 ;
        RECT 252.030 82.110 252.200 83.110 ;
        RECT 241.820 81.880 251.860 82.050 ;
        RECT 252.540 81.380 272.575 83.840 ;
        RECT 240.510 80.710 272.575 81.380 ;
        RECT 240.510 80.690 261.780 80.710 ;
        RECT 240.510 80.645 257.145 80.690 ;
        RECT 240.510 78.185 241.085 80.645 ;
        RECT 241.820 79.975 251.860 80.145 ;
        RECT 241.480 78.915 241.650 79.915 ;
        RECT 252.030 78.915 252.200 79.915 ;
        RECT 241.820 78.685 251.860 78.855 ;
        RECT 252.540 78.185 257.145 80.645 ;
        RECT 229.620 78.050 234.745 78.090 ;
        RECT 126.340 72.155 135.740 72.670 ;
        RECT 66.840 70.450 135.740 72.155 ;
        RECT 66.865 69.750 135.740 70.450 ;
        RECT 229.555 77.400 234.860 78.050 ;
        RECT 229.555 74.990 230.505 77.400 ;
        RECT 231.355 76.780 233.395 76.950 ;
        RECT 230.970 75.720 231.140 76.720 ;
        RECT 233.610 75.720 233.780 76.720 ;
        RECT 231.355 75.490 233.395 75.660 ;
        RECT 234.150 74.990 234.860 77.400 ;
        RECT 229.555 74.255 234.860 74.990 ;
        RECT 229.555 71.795 230.505 74.255 ;
        RECT 231.355 73.585 233.395 73.755 ;
        RECT 230.970 72.525 231.140 73.525 ;
        RECT 233.610 72.525 233.780 73.525 ;
        RECT 231.355 72.295 233.395 72.465 ;
        RECT 234.150 71.795 234.860 74.255 ;
        RECT 229.555 71.055 234.860 71.795 ;
        RECT 192.975 68.715 224.570 68.870 ;
        RECT 191.640 67.545 224.570 68.715 ;
        RECT 229.555 68.600 230.505 71.055 ;
        RECT 231.355 70.390 233.395 70.560 ;
        RECT 230.970 69.330 231.140 70.330 ;
        RECT 233.610 69.330 233.780 70.330 ;
        RECT 231.355 69.100 233.395 69.270 ;
        RECT 234.150 68.600 234.860 71.055 ;
        RECT 229.555 67.865 234.860 68.600 ;
        RECT 48.365 59.425 63.255 59.460 ;
        RECT 48.365 59.385 63.320 59.425 ;
        RECT 48.300 57.850 63.320 59.385 ;
        RECT 48.300 55.265 49.495 57.850 ;
        RECT 49.960 57.190 60.010 57.360 ;
        RECT 49.730 55.935 49.900 56.975 ;
        RECT 60.070 55.935 60.240 56.975 ;
        RECT 49.960 55.550 60.010 55.720 ;
        RECT 60.620 55.265 63.320 57.850 ;
        RECT 72.205 59.285 77.600 59.970 ;
        RECT 72.205 56.885 72.980 59.285 ;
        RECT 73.405 58.890 73.905 59.060 ;
        RECT 74.195 58.890 74.695 59.060 ;
        RECT 74.985 58.890 75.485 59.060 ;
        RECT 75.775 58.890 76.275 59.060 ;
        RECT 73.175 57.635 73.345 58.675 ;
        RECT 73.965 57.635 74.135 58.675 ;
        RECT 74.755 57.635 74.925 58.675 ;
        RECT 75.545 57.635 75.715 58.675 ;
        RECT 76.335 57.635 76.505 58.675 ;
        RECT 73.405 57.250 73.905 57.420 ;
        RECT 74.195 57.250 74.695 57.420 ;
        RECT 74.985 57.250 75.485 57.420 ;
        RECT 75.775 57.250 76.275 57.420 ;
        RECT 76.825 56.885 77.600 59.285 ;
        RECT 191.640 57.135 194.575 67.545 ;
        RECT 195.210 66.860 196.210 67.030 ;
        RECT 196.500 66.860 197.500 67.030 ;
        RECT 197.790 66.860 198.790 67.030 ;
        RECT 199.080 66.860 200.080 67.030 ;
        RECT 200.370 66.860 201.370 67.030 ;
        RECT 201.660 66.860 202.660 67.030 ;
        RECT 202.950 66.860 203.950 67.030 ;
        RECT 204.240 66.860 205.240 67.030 ;
        RECT 205.530 66.860 206.530 67.030 ;
        RECT 206.820 66.860 207.820 67.030 ;
        RECT 165.430 56.905 194.575 57.135 ;
        RECT 72.190 56.090 77.600 56.885 ;
        RECT 165.420 55.820 194.575 56.905 ;
        RECT 38.485 53.955 63.320 55.265 ;
        RECT 38.485 50.360 39.345 53.955 ;
        RECT 39.960 53.375 59.960 53.545 ;
        RECT 39.730 51.120 39.900 53.160 ;
        RECT 60.020 51.120 60.190 53.160 ;
        RECT 39.960 50.735 59.960 50.905 ;
        RECT 60.620 50.360 63.320 53.955 ;
        RECT 38.485 49.125 63.320 50.360 ;
        RECT 69.150 53.460 80.340 53.905 ;
        RECT 69.150 50.835 69.655 53.460 ;
        RECT 70.325 52.770 70.825 52.940 ;
        RECT 70.095 51.560 70.265 52.600 ;
        RECT 70.885 51.560 71.055 52.600 ;
        RECT 70.325 51.220 70.825 51.390 ;
        RECT 71.555 50.835 72.375 53.460 ;
        RECT 73.105 52.770 73.605 52.940 ;
        RECT 72.875 51.560 73.045 52.600 ;
        RECT 73.665 51.560 73.835 52.600 ;
        RECT 73.105 51.220 73.605 51.390 ;
        RECT 74.335 50.835 75.155 53.460 ;
        RECT 75.885 52.770 76.385 52.940 ;
        RECT 75.655 51.560 75.825 52.600 ;
        RECT 76.445 51.560 76.615 52.600 ;
        RECT 75.885 51.220 76.385 51.390 ;
        RECT 77.110 50.835 77.935 53.460 ;
        RECT 78.665 52.770 79.165 52.940 ;
        RECT 78.435 51.560 78.605 52.600 ;
        RECT 79.225 51.560 79.395 52.600 ;
        RECT 78.665 51.220 79.165 51.390 ;
        RECT 79.885 50.835 80.340 53.460 ;
        RECT 161.315 51.555 161.975 51.585 ;
        RECT 165.430 51.555 166.430 55.820 ;
        RECT 167.030 55.200 168.030 55.370 ;
        RECT 168.320 55.200 169.320 55.370 ;
        RECT 169.610 55.200 170.610 55.370 ;
        RECT 170.900 55.200 171.900 55.370 ;
        RECT 172.190 55.200 173.190 55.370 ;
        RECT 173.480 55.200 174.480 55.370 ;
        RECT 174.770 55.200 175.770 55.370 ;
        RECT 176.060 55.200 177.060 55.370 ;
        RECT 177.350 55.200 178.350 55.370 ;
        RECT 178.640 55.200 179.640 55.370 ;
        RECT 69.150 50.035 80.340 50.835 ;
        RECT 145.475 51.290 146.555 51.320 ;
        RECT 145.475 51.275 159.245 51.290 ;
        RECT 38.485 44.785 39.910 49.125 ;
        RECT 40.520 48.445 42.920 48.615 ;
        RECT 40.290 45.690 40.460 48.230 ;
        RECT 42.980 45.690 43.150 48.230 ;
        RECT 40.520 45.305 42.920 45.475 ;
        RECT 43.580 44.785 44.590 49.125 ;
        RECT 45.200 48.445 47.600 48.615 ;
        RECT 44.970 45.690 45.140 48.230 ;
        RECT 47.660 45.690 47.830 48.230 ;
        RECT 45.200 45.305 47.600 45.475 ;
        RECT 48.185 45.020 54.255 49.125 ;
        RECT 54.850 48.535 57.250 48.705 ;
        RECT 54.620 45.780 54.790 48.320 ;
        RECT 57.310 45.780 57.480 48.320 ;
        RECT 54.850 45.395 57.250 45.565 ;
        RECT 57.970 45.020 58.890 49.125 ;
        RECT 59.510 48.535 61.910 48.705 ;
        RECT 59.280 45.780 59.450 48.320 ;
        RECT 61.970 45.780 62.140 48.320 ;
        RECT 59.510 45.395 61.910 45.565 ;
        RECT 62.530 45.020 63.320 49.125 ;
        RECT 48.185 44.785 63.320 45.020 ;
        RECT 38.485 44.615 63.320 44.785 ;
        RECT 38.485 44.095 39.910 44.615 ;
        RECT 43.580 44.095 44.590 44.615 ;
        RECT 48.185 44.095 63.320 44.615 ;
        RECT 38.485 43.925 63.320 44.095 ;
        RECT 38.485 39.760 39.910 43.925 ;
        RECT 40.520 43.235 42.920 43.405 ;
        RECT 40.290 40.480 40.460 43.020 ;
        RECT 42.980 40.480 43.150 43.020 ;
        RECT 40.520 40.095 42.920 40.265 ;
        RECT 43.580 39.760 44.590 43.925 ;
        RECT 48.185 43.760 63.320 43.925 ;
        RECT 45.200 43.235 47.600 43.405 ;
        RECT 44.970 40.480 45.140 43.020 ;
        RECT 47.660 40.480 47.830 43.020 ;
        RECT 45.200 40.095 47.600 40.265 ;
        RECT 48.185 39.760 54.255 43.760 ;
        RECT 54.850 43.110 57.250 43.280 ;
        RECT 54.620 40.355 54.790 42.895 ;
        RECT 57.310 40.355 57.480 42.895 ;
        RECT 54.850 39.970 57.250 40.140 ;
        RECT 38.485 39.725 54.440 39.760 ;
        RECT 57.970 39.725 58.890 43.760 ;
        RECT 59.510 43.110 61.910 43.280 ;
        RECT 59.280 40.355 59.450 42.895 ;
        RECT 61.970 40.355 62.140 42.895 ;
        RECT 59.510 39.970 61.910 40.140 ;
        RECT 62.530 39.725 63.320 43.760 ;
        RECT 38.485 39.085 63.320 39.725 ;
        RECT 38.485 39.050 39.910 39.085 ;
        RECT 53.425 39.050 63.320 39.085 ;
        RECT 86.095 49.420 130.420 50.660 ;
        RECT 53.425 39.045 63.245 39.050 ;
        RECT 53.470 39.025 63.245 39.045 ;
        RECT 62.640 38.980 63.245 39.025 ;
        RECT 43.505 38.595 44.665 38.615 ;
        RECT 53.985 38.595 63.475 38.615 ;
        RECT 35.775 38.055 63.475 38.595 ;
        RECT 35.775 35.565 36.315 38.055 ;
        RECT 36.920 37.525 42.920 37.695 ;
        RECT 36.690 36.315 36.860 37.355 ;
        RECT 42.980 36.315 43.150 37.355 ;
        RECT 36.920 35.975 42.920 36.145 ;
        RECT 43.505 35.565 44.665 38.055 ;
        RECT 51.840 38.035 63.475 38.055 ;
        RECT 45.200 37.525 51.200 37.695 ;
        RECT 44.970 36.315 45.140 37.355 ;
        RECT 51.260 36.315 51.430 37.355 ;
        RECT 45.200 35.975 51.200 36.145 ;
        RECT 51.840 35.630 54.200 38.035 ;
        RECT 54.850 37.525 57.050 37.695 ;
        RECT 54.620 36.315 54.790 37.355 ;
        RECT 57.110 36.315 57.280 37.355 ;
        RECT 54.850 35.975 57.050 36.145 ;
        RECT 57.635 35.630 59.140 38.035 ;
        RECT 59.710 37.530 61.910 37.700 ;
        RECT 59.480 36.320 59.650 37.360 ;
        RECT 61.970 36.320 62.140 37.360 ;
        RECT 59.710 35.980 61.910 36.150 ;
        RECT 62.550 35.630 63.475 38.035 ;
        RECT 51.840 35.565 63.495 35.630 ;
        RECT 35.775 34.795 63.495 35.565 ;
        RECT 35.775 34.520 52.525 34.795 ;
        RECT 62.550 34.770 63.475 34.795 ;
        RECT 35.775 32.010 36.315 34.520 ;
        RECT 36.920 33.945 42.920 34.115 ;
        RECT 36.690 32.735 36.860 33.775 ;
        RECT 42.980 32.735 43.150 33.775 ;
        RECT 36.920 32.395 42.920 32.565 ;
        RECT 43.505 32.010 44.665 34.520 ;
        RECT 45.200 33.945 51.200 34.115 ;
        RECT 44.970 32.735 45.140 33.775 ;
        RECT 51.260 32.735 51.430 33.775 ;
        RECT 45.200 32.395 51.200 32.565 ;
        RECT 51.840 32.010 52.525 34.520 ;
        RECT 35.775 30.965 52.525 32.010 ;
        RECT 35.775 28.390 36.315 30.965 ;
        RECT 36.920 30.365 42.920 30.535 ;
        RECT 36.690 29.155 36.860 30.195 ;
        RECT 42.980 29.155 43.150 30.195 ;
        RECT 36.920 28.815 42.920 28.985 ;
        RECT 43.505 28.390 44.665 30.965 ;
        RECT 45.200 30.365 51.200 30.535 ;
        RECT 44.970 29.155 45.140 30.195 ;
        RECT 51.260 29.155 51.430 30.195 ;
        RECT 45.200 28.815 51.200 28.985 ;
        RECT 51.840 28.390 52.525 30.965 ;
        RECT 35.775 27.345 52.525 28.390 ;
        RECT 35.775 24.895 36.315 27.345 ;
        RECT 36.920 26.785 42.920 26.955 ;
        RECT 36.690 25.575 36.860 26.615 ;
        RECT 42.980 25.575 43.150 26.615 ;
        RECT 36.920 25.235 42.920 25.405 ;
        RECT 43.505 24.895 44.665 27.345 ;
        RECT 45.200 26.785 51.200 26.955 ;
        RECT 44.970 25.575 45.140 26.615 ;
        RECT 51.260 25.575 51.430 26.615 ;
        RECT 45.200 25.235 51.200 25.405 ;
        RECT 51.840 24.895 52.525 27.345 ;
        RECT 35.775 23.885 52.525 24.895 ;
        RECT 51.840 23.865 52.525 23.885 ;
        RECT 86.095 31.155 92.325 49.420 ;
        RECT 93.015 48.860 103.055 49.030 ;
        RECT 92.675 48.300 92.845 48.800 ;
        RECT 103.225 48.300 103.395 48.800 ;
        RECT 93.015 48.070 103.055 48.240 ;
        RECT 92.675 47.510 92.845 48.010 ;
        RECT 103.225 47.510 103.395 48.010 ;
        RECT 93.015 47.280 103.055 47.450 ;
        RECT 103.810 47.275 130.420 49.420 ;
        RECT 92.675 46.720 92.845 47.220 ;
        RECT 103.225 46.720 103.395 47.220 ;
        RECT 93.015 46.490 103.055 46.660 ;
        RECT 92.675 45.930 92.845 46.430 ;
        RECT 103.225 45.930 103.395 46.430 ;
        RECT 103.810 45.965 109.825 47.275 ;
        RECT 110.280 46.445 112.440 46.795 ;
        RECT 126.280 46.445 128.440 46.795 ;
        RECT 128.775 45.965 130.420 47.275 ;
        RECT 93.015 45.700 103.055 45.870 ;
        RECT 103.810 45.795 130.420 45.965 ;
        RECT 92.675 45.140 92.845 45.640 ;
        RECT 103.225 45.140 103.395 45.640 ;
        RECT 93.015 44.910 103.055 45.080 ;
        RECT 92.675 44.350 92.845 44.850 ;
        RECT 103.225 44.350 103.395 44.850 ;
        RECT 103.810 44.485 109.825 45.795 ;
        RECT 110.280 44.965 112.440 45.315 ;
        RECT 126.280 44.965 128.440 45.315 ;
        RECT 128.775 44.485 130.420 45.795 ;
        RECT 103.810 44.315 130.420 44.485 ;
        RECT 93.015 44.120 103.055 44.290 ;
        RECT 92.675 43.560 92.845 44.060 ;
        RECT 103.225 43.560 103.395 44.060 ;
        RECT 93.015 43.330 103.055 43.500 ;
        RECT 92.675 42.770 92.845 43.270 ;
        RECT 103.225 42.770 103.395 43.270 ;
        RECT 103.810 43.005 109.825 44.315 ;
        RECT 110.280 43.485 112.440 43.835 ;
        RECT 126.280 43.485 128.440 43.835 ;
        RECT 128.775 43.005 130.420 44.315 ;
        RECT 103.810 42.835 130.420 43.005 ;
        RECT 93.015 42.540 103.055 42.710 ;
        RECT 92.675 41.980 92.845 42.480 ;
        RECT 103.225 41.980 103.395 42.480 ;
        RECT 93.015 41.750 103.055 41.920 ;
        RECT 92.675 41.190 92.845 41.690 ;
        RECT 103.225 41.190 103.395 41.690 ;
        RECT 103.810 41.540 109.825 42.835 ;
        RECT 110.280 42.005 112.440 42.355 ;
        RECT 126.280 42.005 128.440 42.355 ;
        RECT 128.775 41.540 130.420 42.835 ;
        RECT 93.015 40.960 103.055 41.130 ;
        RECT 92.675 40.400 92.845 40.900 ;
        RECT 103.225 40.400 103.395 40.900 ;
        RECT 93.015 40.170 103.055 40.340 ;
        RECT 92.675 39.610 92.845 40.110 ;
        RECT 103.225 39.610 103.395 40.110 ;
        RECT 103.810 39.615 130.420 41.540 ;
        RECT 103.810 39.580 116.720 39.615 ;
        RECT 93.015 39.380 103.055 39.550 ;
        RECT 92.675 38.820 92.845 39.320 ;
        RECT 103.225 38.820 103.395 39.320 ;
        RECT 93.015 38.590 103.055 38.760 ;
        RECT 92.675 38.030 92.845 38.530 ;
        RECT 103.225 38.030 103.395 38.530 ;
        RECT 93.015 37.800 103.055 37.970 ;
        RECT 92.675 37.240 92.845 37.740 ;
        RECT 103.225 37.240 103.395 37.740 ;
        RECT 93.015 37.010 103.055 37.180 ;
        RECT 92.675 36.450 92.845 36.950 ;
        RECT 103.225 36.450 103.395 36.950 ;
        RECT 103.810 36.820 105.155 39.580 ;
        RECT 105.820 38.890 115.820 39.060 ;
        RECT 105.590 37.680 105.760 38.720 ;
        RECT 115.880 37.680 116.050 38.720 ;
        RECT 105.820 37.340 115.820 37.510 ;
        RECT 116.550 36.820 116.720 39.580 ;
        RECT 103.810 36.650 116.720 36.820 ;
        RECT 93.015 36.220 103.055 36.390 ;
        RECT 92.675 35.660 92.845 36.160 ;
        RECT 103.225 35.660 103.395 36.160 ;
        RECT 93.015 35.430 103.055 35.600 ;
        RECT 92.675 34.870 92.845 35.370 ;
        RECT 103.225 34.870 103.395 35.370 ;
        RECT 93.015 34.640 103.055 34.810 ;
        RECT 92.675 34.080 92.845 34.580 ;
        RECT 103.225 34.080 103.395 34.580 ;
        RECT 93.015 33.850 103.055 34.020 ;
        RECT 103.810 33.890 105.155 36.650 ;
        RECT 105.820 35.960 115.820 36.130 ;
        RECT 105.590 34.750 105.760 35.790 ;
        RECT 115.880 34.750 116.050 35.790 ;
        RECT 105.820 34.410 115.820 34.580 ;
        RECT 116.550 33.890 116.720 36.650 ;
        RECT 92.675 33.290 92.845 33.790 ;
        RECT 103.225 33.290 103.395 33.790 ;
        RECT 103.810 33.720 116.720 33.890 ;
        RECT 93.015 33.060 103.055 33.230 ;
        RECT 92.675 32.500 92.845 33.000 ;
        RECT 103.225 32.500 103.395 33.000 ;
        RECT 93.015 32.270 103.055 32.440 ;
        RECT 92.675 31.710 92.845 32.210 ;
        RECT 103.225 31.710 103.395 32.210 ;
        RECT 93.015 31.480 103.055 31.650 ;
        RECT 103.810 31.155 105.155 33.720 ;
        RECT 105.820 33.030 115.820 33.200 ;
        RECT 105.590 31.820 105.760 32.860 ;
        RECT 115.880 31.820 116.050 32.860 ;
        RECT 105.820 31.480 115.820 31.650 ;
        RECT 116.550 31.155 116.720 33.720 ;
        RECT 117.230 39.580 130.420 39.615 ;
        RECT 117.230 36.820 117.400 39.580 ;
        RECT 118.130 38.890 128.130 39.060 ;
        RECT 117.900 37.680 118.070 38.720 ;
        RECT 128.190 37.680 128.360 38.720 ;
        RECT 118.130 37.340 128.130 37.510 ;
        RECT 128.775 36.820 130.420 39.580 ;
        RECT 117.230 36.650 130.420 36.820 ;
        RECT 117.230 33.890 117.400 36.650 ;
        RECT 118.130 35.960 128.130 36.130 ;
        RECT 117.900 34.750 118.070 35.790 ;
        RECT 128.190 34.750 128.360 35.790 ;
        RECT 118.130 34.410 128.130 34.580 ;
        RECT 128.775 33.890 130.420 36.650 ;
        RECT 117.230 33.720 130.420 33.890 ;
        RECT 117.230 31.155 117.400 33.720 ;
        RECT 118.130 33.030 128.130 33.200 ;
        RECT 117.900 31.820 118.070 32.860 ;
        RECT 128.190 31.820 128.360 32.860 ;
        RECT 118.130 31.480 128.130 31.650 ;
        RECT 128.775 31.155 130.420 33.720 ;
        RECT 86.095 30.085 130.420 31.155 ;
        RECT 86.095 28.800 87.530 30.085 ;
        RECT 92.110 30.025 130.420 30.085 ;
        RECT 87.990 29.280 90.150 29.630 ;
        RECT 105.490 29.280 107.650 29.630 ;
        RECT 108.130 28.800 108.300 30.025 ;
        RECT 108.780 29.280 110.940 29.630 ;
        RECT 126.280 29.280 128.440 29.630 ;
        RECT 128.775 28.800 130.420 30.025 ;
        RECT 86.095 28.630 130.420 28.800 ;
        RECT 86.095 27.320 87.530 28.630 ;
        RECT 87.990 27.800 90.150 28.150 ;
        RECT 105.490 27.800 107.650 28.150 ;
        RECT 108.130 27.320 108.300 28.630 ;
        RECT 108.780 27.800 110.940 28.150 ;
        RECT 126.280 27.800 128.440 28.150 ;
        RECT 128.775 27.320 130.420 28.630 ;
        RECT 145.475 50.215 159.255 51.275 ;
        RECT 161.310 51.205 166.430 51.555 ;
        RECT 161.310 50.575 166.380 51.205 ;
        RECT 145.475 39.850 146.600 50.215 ;
        RECT 147.350 49.640 157.390 49.810 ;
        RECT 147.010 40.580 147.180 49.580 ;
        RECT 157.560 40.580 157.730 49.580 ;
        RECT 147.350 40.350 157.390 40.520 ;
        RECT 158.170 39.850 159.255 50.215 ;
        RECT 161.315 44.905 162.060 50.575 ;
        RECT 162.660 49.935 163.660 50.105 ;
        RECT 162.430 45.680 162.600 49.720 ;
        RECT 163.720 45.680 163.890 49.720 ;
        RECT 162.660 45.295 163.660 45.465 ;
        RECT 164.355 44.905 166.380 50.575 ;
        RECT 166.800 44.945 166.970 54.985 ;
        RECT 168.090 44.945 168.260 54.985 ;
        RECT 169.380 44.945 169.550 54.985 ;
        RECT 170.670 44.945 170.840 54.985 ;
        RECT 171.960 44.945 172.130 54.985 ;
        RECT 173.250 44.945 173.420 54.985 ;
        RECT 174.540 44.945 174.710 54.985 ;
        RECT 175.830 44.945 176.000 54.985 ;
        RECT 177.120 44.945 177.290 54.985 ;
        RECT 178.410 44.945 178.580 54.985 ;
        RECT 179.700 44.945 179.870 54.985 ;
        RECT 161.315 44.245 166.380 44.905 ;
        RECT 167.030 44.560 168.030 44.730 ;
        RECT 168.320 44.560 169.320 44.730 ;
        RECT 169.610 44.560 170.610 44.730 ;
        RECT 170.900 44.560 171.900 44.730 ;
        RECT 172.190 44.560 173.190 44.730 ;
        RECT 173.480 44.560 174.480 44.730 ;
        RECT 174.770 44.560 175.770 44.730 ;
        RECT 176.060 44.560 177.060 44.730 ;
        RECT 177.350 44.560 178.350 44.730 ;
        RECT 178.640 44.560 179.640 44.730 ;
        RECT 161.355 44.085 166.380 44.245 ;
        RECT 180.320 44.085 181.440 55.820 ;
        RECT 182.095 55.200 183.095 55.370 ;
        RECT 183.385 55.200 184.385 55.370 ;
        RECT 184.675 55.200 185.675 55.370 ;
        RECT 185.965 55.200 186.965 55.370 ;
        RECT 187.255 55.200 188.255 55.370 ;
        RECT 181.865 44.945 182.035 54.985 ;
        RECT 183.155 44.945 183.325 54.985 ;
        RECT 184.445 44.945 184.615 54.985 ;
        RECT 185.735 44.945 185.905 54.985 ;
        RECT 187.025 44.945 187.195 54.985 ;
        RECT 188.315 44.945 188.485 54.985 ;
        RECT 188.875 50.735 194.575 55.820 ;
        RECT 182.095 44.560 183.095 44.730 ;
        RECT 183.385 44.560 184.385 44.730 ;
        RECT 184.675 44.560 185.675 44.730 ;
        RECT 185.965 44.560 186.965 44.730 ;
        RECT 187.255 44.560 188.255 44.730 ;
        RECT 188.875 44.085 190.025 50.735 ;
        RECT 190.705 50.105 191.705 50.275 ;
        RECT 191.995 50.105 192.995 50.275 ;
        RECT 190.475 44.850 190.645 49.890 ;
        RECT 191.765 44.850 191.935 49.890 ;
        RECT 193.055 44.850 193.225 49.890 ;
        RECT 190.705 44.465 191.705 44.635 ;
        RECT 191.995 44.465 192.995 44.635 ;
        RECT 161.355 44.025 190.025 44.085 ;
        RECT 193.670 44.025 194.575 50.735 ;
        RECT 161.355 43.640 194.695 44.025 ;
        RECT 161.360 42.860 194.695 43.640 ;
        RECT 145.475 39.680 159.255 39.850 ;
        RECT 145.475 39.280 146.600 39.680 ;
        RECT 158.170 39.280 159.255 39.680 ;
        RECT 145.475 39.110 159.255 39.280 ;
        RECT 145.475 28.775 146.600 39.110 ;
        RECT 147.350 38.440 157.390 38.610 ;
        RECT 147.010 29.380 147.180 38.380 ;
        RECT 157.560 29.380 157.730 38.380 ;
        RECT 158.170 31.010 159.255 39.110 ;
        RECT 165.445 32.845 166.315 42.860 ;
        RECT 167.025 42.315 168.025 42.485 ;
        RECT 168.315 42.315 169.315 42.485 ;
        RECT 169.605 42.315 170.605 42.485 ;
        RECT 170.895 42.315 171.895 42.485 ;
        RECT 172.185 42.315 173.185 42.485 ;
        RECT 173.475 42.315 174.475 42.485 ;
        RECT 174.765 42.315 175.765 42.485 ;
        RECT 176.055 42.315 177.055 42.485 ;
        RECT 166.795 33.560 166.965 42.100 ;
        RECT 168.085 33.560 168.255 42.100 ;
        RECT 169.375 33.560 169.545 42.100 ;
        RECT 170.665 33.560 170.835 42.100 ;
        RECT 171.955 33.560 172.125 42.100 ;
        RECT 173.245 33.560 173.415 42.100 ;
        RECT 174.535 33.560 174.705 42.100 ;
        RECT 175.825 33.560 175.995 42.100 ;
        RECT 177.115 33.560 177.285 42.100 ;
        RECT 177.770 40.840 194.695 42.860 ;
        RECT 194.980 41.605 195.150 66.645 ;
        RECT 196.270 41.605 196.440 66.645 ;
        RECT 197.560 41.605 197.730 66.645 ;
        RECT 198.850 41.605 199.020 66.645 ;
        RECT 200.140 41.605 200.310 66.645 ;
        RECT 201.430 41.605 201.600 66.645 ;
        RECT 202.720 41.605 202.890 66.645 ;
        RECT 204.010 41.605 204.180 66.645 ;
        RECT 205.300 41.605 205.470 66.645 ;
        RECT 206.590 41.605 206.760 66.645 ;
        RECT 207.880 41.605 208.050 66.645 ;
        RECT 195.210 41.220 196.210 41.390 ;
        RECT 196.500 41.220 197.500 41.390 ;
        RECT 197.790 41.220 198.790 41.390 ;
        RECT 199.080 41.220 200.080 41.390 ;
        RECT 200.370 41.220 201.370 41.390 ;
        RECT 201.660 41.220 202.660 41.390 ;
        RECT 202.950 41.220 203.950 41.390 ;
        RECT 204.240 41.220 205.240 41.390 ;
        RECT 205.530 41.220 206.530 41.390 ;
        RECT 206.820 41.220 207.820 41.390 ;
        RECT 208.395 40.840 209.475 67.545 ;
        RECT 210.050 66.860 211.050 67.030 ;
        RECT 211.340 66.860 212.340 67.030 ;
        RECT 212.630 66.860 213.630 67.030 ;
        RECT 213.920 66.860 214.920 67.030 ;
        RECT 215.210 66.860 216.210 67.030 ;
        RECT 216.500 66.860 217.500 67.030 ;
        RECT 217.790 66.860 218.790 67.030 ;
        RECT 219.080 66.860 220.080 67.030 ;
        RECT 220.370 66.860 221.370 67.030 ;
        RECT 221.660 66.860 222.660 67.030 ;
        RECT 209.820 41.605 209.990 66.645 ;
        RECT 211.110 41.605 211.280 66.645 ;
        RECT 212.400 41.605 212.570 66.645 ;
        RECT 213.690 41.605 213.860 66.645 ;
        RECT 214.980 41.605 215.150 66.645 ;
        RECT 216.270 41.605 216.440 66.645 ;
        RECT 217.560 41.605 217.730 66.645 ;
        RECT 218.850 41.605 219.020 66.645 ;
        RECT 220.140 41.605 220.310 66.645 ;
        RECT 221.430 41.605 221.600 66.645 ;
        RECT 222.720 41.605 222.890 66.645 ;
        RECT 210.050 41.220 211.050 41.390 ;
        RECT 211.340 41.220 212.340 41.390 ;
        RECT 212.630 41.220 213.630 41.390 ;
        RECT 213.920 41.220 214.920 41.390 ;
        RECT 215.210 41.220 216.210 41.390 ;
        RECT 216.500 41.220 217.500 41.390 ;
        RECT 217.790 41.220 218.790 41.390 ;
        RECT 219.080 41.220 220.080 41.390 ;
        RECT 220.370 41.220 221.370 41.390 ;
        RECT 221.660 41.220 222.660 41.390 ;
        RECT 223.260 40.840 224.510 67.545 ;
        RECT 177.770 40.760 224.510 40.840 ;
        RECT 177.770 35.005 181.975 40.760 ;
        RECT 182.475 40.090 183.475 40.260 ;
        RECT 183.765 40.090 184.765 40.260 ;
        RECT 182.245 35.835 182.415 39.875 ;
        RECT 183.535 35.835 183.705 39.875 ;
        RECT 184.825 35.835 184.995 39.875 ;
        RECT 185.400 39.705 224.510 40.760 ;
        RECT 185.400 38.815 194.695 39.705 ;
        RECT 195.210 39.105 196.210 39.275 ;
        RECT 196.500 39.105 197.500 39.275 ;
        RECT 197.790 39.105 198.790 39.275 ;
        RECT 199.080 39.105 200.080 39.275 ;
        RECT 200.370 39.105 201.370 39.275 ;
        RECT 201.660 39.105 202.660 39.275 ;
        RECT 202.950 39.105 203.950 39.275 ;
        RECT 204.240 39.105 205.240 39.275 ;
        RECT 205.530 39.105 206.530 39.275 ;
        RECT 206.820 39.105 207.820 39.275 ;
        RECT 185.400 36.055 190.380 38.815 ;
        RECT 190.980 38.215 192.980 38.385 ;
        RECT 190.750 36.960 190.920 38.000 ;
        RECT 193.040 36.960 193.210 38.000 ;
        RECT 190.980 36.575 192.980 36.745 ;
        RECT 193.685 36.055 194.695 38.815 ;
        RECT 182.475 35.450 183.475 35.620 ;
        RECT 183.765 35.450 184.765 35.620 ;
        RECT 185.400 35.005 194.695 36.055 ;
        RECT 177.770 34.380 194.695 35.005 ;
        RECT 167.025 33.175 168.025 33.345 ;
        RECT 168.315 33.175 169.315 33.345 ;
        RECT 169.605 33.175 170.605 33.345 ;
        RECT 170.895 33.175 171.895 33.345 ;
        RECT 172.185 33.175 173.185 33.345 ;
        RECT 173.475 33.175 174.475 33.345 ;
        RECT 174.765 33.175 175.765 33.345 ;
        RECT 176.055 33.175 177.055 33.345 ;
        RECT 177.770 32.845 194.655 34.380 ;
        RECT 165.445 31.970 194.655 32.845 ;
        RECT 165.720 31.955 194.655 31.970 ;
        RECT 177.775 31.930 194.655 31.955 ;
        RECT 180.770 31.890 194.655 31.930 ;
        RECT 158.170 29.670 174.475 31.010 ;
        RECT 147.350 29.150 157.390 29.320 ;
        RECT 158.170 28.775 161.925 29.670 ;
        RECT 162.770 29.150 172.810 29.320 ;
        RECT 145.475 28.510 161.970 28.775 ;
        RECT 86.095 27.150 130.420 27.320 ;
        RECT 86.095 25.840 87.530 27.150 ;
        RECT 87.990 26.320 90.150 26.670 ;
        RECT 105.490 26.320 107.650 26.670 ;
        RECT 108.130 25.840 108.300 27.150 ;
        RECT 108.780 26.320 110.940 26.670 ;
        RECT 126.280 26.320 128.440 26.670 ;
        RECT 128.775 25.840 130.420 27.150 ;
        RECT 145.480 26.165 161.970 28.510 ;
        RECT 145.480 26.020 161.975 26.165 ;
        RECT 86.095 25.670 130.420 25.840 ;
        RECT 86.095 24.360 87.530 25.670 ;
        RECT 87.990 24.840 90.150 25.190 ;
        RECT 105.490 24.840 107.650 25.190 ;
        RECT 108.130 24.360 108.300 25.670 ;
        RECT 108.780 24.840 110.940 25.190 ;
        RECT 126.280 24.840 128.440 25.190 ;
        RECT 128.775 24.360 130.420 25.670 ;
        RECT 86.095 24.190 130.420 24.360 ;
        RECT 86.095 22.880 87.530 24.190 ;
        RECT 87.990 23.360 90.150 23.710 ;
        RECT 105.490 23.360 107.650 23.710 ;
        RECT 108.130 22.880 108.300 24.190 ;
        RECT 108.780 23.360 110.940 23.710 ;
        RECT 126.280 23.360 128.440 23.710 ;
        RECT 128.775 22.880 130.420 24.190 ;
        RECT 86.095 22.710 130.420 22.880 ;
        RECT 86.095 21.400 87.530 22.710 ;
        RECT 87.990 21.880 90.150 22.230 ;
        RECT 105.490 21.880 107.650 22.230 ;
        RECT 108.130 21.400 108.300 22.710 ;
        RECT 108.780 21.880 110.940 22.230 ;
        RECT 126.280 21.880 128.440 22.230 ;
        RECT 128.775 21.400 130.420 22.710 ;
        RECT 86.095 21.230 130.420 21.400 ;
        RECT 86.095 19.920 87.530 21.230 ;
        RECT 87.990 20.400 90.150 20.750 ;
        RECT 105.490 20.400 107.650 20.750 ;
        RECT 108.130 19.920 108.300 21.230 ;
        RECT 108.780 20.400 110.940 20.750 ;
        RECT 126.280 20.400 128.440 20.750 ;
        RECT 128.775 19.920 130.420 21.230 ;
        RECT 86.095 19.750 130.420 19.920 ;
        RECT 86.095 18.480 87.530 19.750 ;
        RECT 87.990 18.920 90.150 19.270 ;
        RECT 105.490 18.920 107.650 19.270 ;
        RECT 108.130 18.480 108.300 19.750 ;
        RECT 108.780 18.920 110.940 19.270 ;
        RECT 126.280 18.920 128.440 19.270 ;
        RECT 128.775 18.480 130.420 19.750 ;
        RECT 145.485 25.605 161.975 26.020 ;
        RECT 145.485 19.240 146.290 25.605 ;
        RECT 146.900 25.005 147.900 25.175 ;
        RECT 148.190 25.005 149.190 25.175 ;
        RECT 149.480 25.005 150.480 25.175 ;
        RECT 150.770 25.005 151.770 25.175 ;
        RECT 152.060 25.005 153.060 25.175 ;
        RECT 153.350 25.005 154.350 25.175 ;
        RECT 154.640 25.005 155.640 25.175 ;
        RECT 155.930 25.005 156.930 25.175 ;
        RECT 157.220 25.005 158.220 25.175 ;
        RECT 158.510 25.005 159.510 25.175 ;
        RECT 146.670 19.795 146.840 24.835 ;
        RECT 147.960 19.795 148.130 24.835 ;
        RECT 149.250 19.795 149.420 24.835 ;
        RECT 150.540 19.795 150.710 24.835 ;
        RECT 151.830 19.795 152.000 24.835 ;
        RECT 153.120 19.795 153.290 24.835 ;
        RECT 154.410 19.795 154.580 24.835 ;
        RECT 155.700 19.795 155.870 24.835 ;
        RECT 156.990 19.795 157.160 24.835 ;
        RECT 158.280 19.795 158.450 24.835 ;
        RECT 159.570 19.795 159.740 24.835 ;
        RECT 146.900 19.455 147.900 19.625 ;
        RECT 148.190 19.455 149.190 19.625 ;
        RECT 149.480 19.455 150.480 19.625 ;
        RECT 150.770 19.455 151.770 19.625 ;
        RECT 152.060 19.455 153.060 19.625 ;
        RECT 153.350 19.455 154.350 19.625 ;
        RECT 154.640 19.455 155.640 19.625 ;
        RECT 155.930 19.455 156.930 19.625 ;
        RECT 157.220 19.455 158.220 19.625 ;
        RECT 158.510 19.455 159.510 19.625 ;
        RECT 160.190 19.605 161.975 25.605 ;
        RECT 162.430 20.090 162.600 29.090 ;
        RECT 172.980 20.090 173.150 29.090 ;
        RECT 162.770 19.860 172.810 20.030 ;
        RECT 173.585 19.605 174.475 29.670 ;
        RECT 160.190 19.240 174.475 19.605 ;
        RECT 193.680 20.045 194.655 31.890 ;
        RECT 194.980 20.850 195.150 38.890 ;
        RECT 196.270 20.850 196.440 38.890 ;
        RECT 197.560 20.850 197.730 38.890 ;
        RECT 198.850 20.850 199.020 38.890 ;
        RECT 200.140 20.850 200.310 38.890 ;
        RECT 201.430 20.850 201.600 38.890 ;
        RECT 202.720 20.850 202.890 38.890 ;
        RECT 204.010 20.850 204.180 38.890 ;
        RECT 205.300 20.850 205.470 38.890 ;
        RECT 206.590 20.850 206.760 38.890 ;
        RECT 207.880 20.850 208.050 38.890 ;
        RECT 195.210 20.465 196.210 20.635 ;
        RECT 196.500 20.465 197.500 20.635 ;
        RECT 197.790 20.465 198.790 20.635 ;
        RECT 199.080 20.465 200.080 20.635 ;
        RECT 200.370 20.465 201.370 20.635 ;
        RECT 201.660 20.465 202.660 20.635 ;
        RECT 202.950 20.465 203.950 20.635 ;
        RECT 204.240 20.465 205.240 20.635 ;
        RECT 205.530 20.465 206.530 20.635 ;
        RECT 206.820 20.465 207.820 20.635 ;
        RECT 208.505 20.045 209.670 39.705 ;
        RECT 210.325 39.030 211.325 39.200 ;
        RECT 211.615 39.030 212.615 39.200 ;
        RECT 212.905 39.030 213.905 39.200 ;
        RECT 214.195 39.030 215.195 39.200 ;
        RECT 215.485 39.030 216.485 39.200 ;
        RECT 216.775 39.030 217.775 39.200 ;
        RECT 218.065 39.030 219.065 39.200 ;
        RECT 219.355 39.030 220.355 39.200 ;
        RECT 220.645 39.030 221.645 39.200 ;
        RECT 221.935 39.030 222.935 39.200 ;
        RECT 210.095 20.775 210.265 38.815 ;
        RECT 211.385 20.775 211.555 38.815 ;
        RECT 212.675 20.775 212.845 38.815 ;
        RECT 213.965 20.775 214.135 38.815 ;
        RECT 215.255 20.775 215.425 38.815 ;
        RECT 216.545 20.775 216.715 38.815 ;
        RECT 217.835 20.775 218.005 38.815 ;
        RECT 219.125 20.775 219.295 38.815 ;
        RECT 220.415 20.775 220.585 38.815 ;
        RECT 221.705 20.775 221.875 38.815 ;
        RECT 222.995 20.775 223.165 38.815 ;
        RECT 210.325 20.390 211.325 20.560 ;
        RECT 211.615 20.390 212.615 20.560 ;
        RECT 212.905 20.390 213.905 20.560 ;
        RECT 214.195 20.390 215.195 20.560 ;
        RECT 215.485 20.390 216.485 20.560 ;
        RECT 216.775 20.390 217.775 20.560 ;
        RECT 218.065 20.390 219.065 20.560 ;
        RECT 219.355 20.390 220.355 20.560 ;
        RECT 220.645 20.390 221.645 20.560 ;
        RECT 221.935 20.390 222.935 20.560 ;
        RECT 223.520 20.045 224.510 39.705 ;
        RECT 86.095 16.895 130.420 18.480 ;
        RECT 145.480 18.435 174.490 19.240 ;
        RECT 193.680 18.940 224.510 20.045 ;
        RECT 229.555 65.405 230.505 67.865 ;
        RECT 231.355 67.195 233.395 67.365 ;
        RECT 230.970 66.135 231.140 67.135 ;
        RECT 233.610 66.135 233.780 67.135 ;
        RECT 231.355 65.905 233.395 66.075 ;
        RECT 234.150 65.405 234.860 67.865 ;
        RECT 229.555 64.670 234.860 65.405 ;
        RECT 229.555 62.210 230.505 64.670 ;
        RECT 231.355 64.000 233.395 64.170 ;
        RECT 230.970 62.940 231.140 63.940 ;
        RECT 233.610 62.940 233.780 63.940 ;
        RECT 231.355 62.710 233.395 62.880 ;
        RECT 234.150 62.210 234.860 64.670 ;
        RECT 229.555 61.475 234.860 62.210 ;
        RECT 229.555 59.015 230.505 61.475 ;
        RECT 231.350 60.805 233.390 60.975 ;
        RECT 230.965 59.745 231.135 60.745 ;
        RECT 233.605 59.745 233.775 60.745 ;
        RECT 231.350 59.515 233.390 59.685 ;
        RECT 234.150 59.015 234.860 61.475 ;
        RECT 229.555 58.280 234.860 59.015 ;
        RECT 229.555 55.820 230.505 58.280 ;
        RECT 231.350 57.610 233.390 57.780 ;
        RECT 230.965 56.550 231.135 57.550 ;
        RECT 233.605 56.550 233.775 57.550 ;
        RECT 231.350 56.320 233.390 56.490 ;
        RECT 234.150 55.820 234.860 58.280 ;
        RECT 229.555 55.085 234.860 55.820 ;
        RECT 229.555 52.625 230.505 55.085 ;
        RECT 231.350 54.415 233.390 54.585 ;
        RECT 230.965 53.355 231.135 54.355 ;
        RECT 233.605 53.355 233.775 54.355 ;
        RECT 231.350 53.125 233.390 53.295 ;
        RECT 234.150 52.625 234.860 55.085 ;
        RECT 229.555 51.890 234.860 52.625 ;
        RECT 229.555 49.430 230.505 51.890 ;
        RECT 231.350 51.220 233.390 51.390 ;
        RECT 230.965 50.160 231.135 51.160 ;
        RECT 233.605 50.160 233.775 51.160 ;
        RECT 231.350 49.930 233.390 50.100 ;
        RECT 234.150 49.430 234.860 51.890 ;
        RECT 229.555 48.690 234.860 49.430 ;
        RECT 229.555 46.235 230.505 48.690 ;
        RECT 231.350 48.025 233.390 48.195 ;
        RECT 230.965 46.965 231.135 47.965 ;
        RECT 233.605 46.965 233.775 47.965 ;
        RECT 231.350 46.735 233.390 46.905 ;
        RECT 234.150 46.235 234.860 48.690 ;
        RECT 229.555 45.500 234.860 46.235 ;
        RECT 229.555 43.040 230.505 45.500 ;
        RECT 231.350 44.830 233.390 45.000 ;
        RECT 230.965 43.770 231.135 44.770 ;
        RECT 233.605 43.770 233.775 44.770 ;
        RECT 231.350 43.540 233.390 43.710 ;
        RECT 234.150 43.040 234.860 45.500 ;
        RECT 229.555 42.305 234.860 43.040 ;
        RECT 229.555 39.845 230.505 42.305 ;
        RECT 231.350 41.635 233.390 41.805 ;
        RECT 230.965 40.575 231.135 41.575 ;
        RECT 233.605 40.575 233.775 41.575 ;
        RECT 231.350 40.345 233.390 40.515 ;
        RECT 234.150 39.845 234.860 42.305 ;
        RECT 229.555 39.110 234.860 39.845 ;
        RECT 229.555 36.650 230.505 39.110 ;
        RECT 231.350 38.440 233.390 38.610 ;
        RECT 230.965 37.380 231.135 38.380 ;
        RECT 233.605 37.380 233.775 38.380 ;
        RECT 231.350 37.150 233.390 37.320 ;
        RECT 234.150 36.650 234.860 39.110 ;
        RECT 229.555 35.915 234.860 36.650 ;
        RECT 229.555 33.455 230.505 35.915 ;
        RECT 231.350 35.245 233.390 35.415 ;
        RECT 230.965 34.185 231.135 35.185 ;
        RECT 233.605 34.185 233.775 35.185 ;
        RECT 231.350 33.955 233.390 34.125 ;
        RECT 234.150 33.455 234.860 35.915 ;
        RECT 229.555 32.720 234.860 33.455 ;
        RECT 229.555 30.260 230.505 32.720 ;
        RECT 231.350 32.050 233.390 32.220 ;
        RECT 230.965 30.990 231.135 31.990 ;
        RECT 233.605 30.990 233.775 31.990 ;
        RECT 231.350 30.760 233.390 30.930 ;
        RECT 234.150 30.260 234.860 32.720 ;
        RECT 229.555 29.525 234.860 30.260 ;
        RECT 229.555 27.065 230.505 29.525 ;
        RECT 231.350 28.855 233.390 29.025 ;
        RECT 230.965 27.795 231.135 28.795 ;
        RECT 233.605 27.795 233.775 28.795 ;
        RECT 231.350 27.565 233.390 27.735 ;
        RECT 234.150 27.065 234.860 29.525 ;
        RECT 229.555 26.330 234.860 27.065 ;
        RECT 229.555 23.875 230.505 26.330 ;
        RECT 231.350 25.660 233.390 25.830 ;
        RECT 230.965 24.600 231.135 25.600 ;
        RECT 233.605 24.600 233.775 25.600 ;
        RECT 231.350 24.370 233.390 24.540 ;
        RECT 234.150 23.875 234.860 26.330 ;
        RECT 229.555 23.140 234.860 23.875 ;
        RECT 229.555 20.680 230.505 23.140 ;
        RECT 231.350 22.470 233.390 22.640 ;
        RECT 230.965 21.410 231.135 22.410 ;
        RECT 233.605 21.410 233.775 22.410 ;
        RECT 231.350 21.180 233.390 21.350 ;
        RECT 234.150 20.680 234.860 23.140 ;
        RECT 229.555 19.875 234.860 20.680 ;
        RECT 240.510 77.450 257.145 78.185 ;
        RECT 257.450 78.050 257.800 80.210 ;
        RECT 240.510 74.990 241.085 77.450 ;
        RECT 241.820 76.780 242.860 76.950 ;
        RECT 243.690 76.770 257.145 77.450 ;
        RECT 241.480 75.720 241.650 76.720 ;
        RECT 243.030 75.720 243.200 76.720 ;
        RECT 241.820 75.490 242.860 75.660 ;
        RECT 243.720 74.990 257.145 76.770 ;
        RECT 240.510 74.255 257.145 74.990 ;
        RECT 240.510 71.795 241.085 74.255 ;
        RECT 241.820 73.585 242.860 73.755 ;
        RECT 241.480 72.525 241.650 73.525 ;
        RECT 243.030 72.525 243.200 73.525 ;
        RECT 241.820 72.295 242.860 72.465 ;
        RECT 243.720 71.795 257.145 74.255 ;
        RECT 240.510 71.060 257.145 71.795 ;
        RECT 240.510 68.600 241.085 71.060 ;
        RECT 241.820 70.390 242.860 70.560 ;
        RECT 241.480 69.330 241.650 70.330 ;
        RECT 243.030 69.330 243.200 70.330 ;
        RECT 241.820 69.100 242.860 69.270 ;
        RECT 243.720 68.600 257.145 71.060 ;
        RECT 240.510 67.865 257.145 68.600 ;
        RECT 240.510 65.405 241.085 67.865 ;
        RECT 241.820 67.195 242.860 67.365 ;
        RECT 241.480 66.135 241.650 67.135 ;
        RECT 243.030 66.135 243.200 67.135 ;
        RECT 241.820 65.905 242.860 66.075 ;
        RECT 243.720 65.405 257.145 67.865 ;
        RECT 240.510 64.670 257.145 65.405 ;
        RECT 240.510 62.210 241.085 64.670 ;
        RECT 241.820 64.000 244.860 64.170 ;
        RECT 241.480 62.940 241.650 63.940 ;
        RECT 245.030 62.940 245.200 63.940 ;
        RECT 241.820 62.710 244.860 62.880 ;
        RECT 245.535 62.210 257.145 64.670 ;
        RECT 240.510 61.475 257.145 62.210 ;
        RECT 240.510 59.015 241.085 61.475 ;
        RECT 241.820 60.805 244.860 60.975 ;
        RECT 241.480 59.745 241.650 60.745 ;
        RECT 245.030 59.745 245.200 60.745 ;
        RECT 241.820 59.515 244.860 59.685 ;
        RECT 245.535 59.015 257.145 61.475 ;
        RECT 240.510 58.280 257.145 59.015 ;
        RECT 240.510 55.820 241.085 58.280 ;
        RECT 241.820 57.610 244.860 57.780 ;
        RECT 241.480 56.550 241.650 57.550 ;
        RECT 245.030 56.550 245.200 57.550 ;
        RECT 241.820 56.320 244.860 56.490 ;
        RECT 245.535 55.820 257.145 58.280 ;
        RECT 240.510 55.085 257.145 55.820 ;
        RECT 240.510 52.625 241.085 55.085 ;
        RECT 241.820 54.415 244.860 54.585 ;
        RECT 241.480 53.355 241.650 54.355 ;
        RECT 245.030 53.355 245.200 54.355 ;
        RECT 241.820 53.125 244.860 53.295 ;
        RECT 245.535 52.625 257.145 55.085 ;
        RECT 240.510 51.890 257.145 52.625 ;
        RECT 240.510 49.430 241.085 51.890 ;
        RECT 241.820 51.220 244.860 51.390 ;
        RECT 241.480 50.160 241.650 51.160 ;
        RECT 245.030 50.160 245.200 51.160 ;
        RECT 245.535 50.620 257.145 51.890 ;
        RECT 257.450 51.100 257.800 53.260 ;
        RECT 258.075 50.620 258.585 80.690 ;
        RECT 258.930 78.050 259.280 80.210 ;
        RECT 258.930 51.100 259.280 53.260 ;
        RECT 259.560 50.620 260.070 80.690 ;
        RECT 260.410 78.050 260.760 80.210 ;
        RECT 260.410 51.100 260.760 53.260 ;
        RECT 261.230 50.620 261.780 80.690 ;
        RECT 245.535 50.450 261.780 50.620 ;
        RECT 241.820 49.930 244.860 50.100 ;
        RECT 245.535 49.430 257.145 50.450 ;
        RECT 240.510 48.695 257.145 49.430 ;
        RECT 240.510 46.235 241.085 48.695 ;
        RECT 241.820 48.025 244.860 48.195 ;
        RECT 241.480 46.965 241.650 47.965 ;
        RECT 245.030 46.965 245.200 47.965 ;
        RECT 241.820 46.735 244.860 46.905 ;
        RECT 245.535 46.235 257.145 48.695 ;
        RECT 257.450 47.810 257.800 49.970 ;
        RECT 240.510 45.500 257.145 46.235 ;
        RECT 240.510 43.040 241.085 45.500 ;
        RECT 241.820 44.830 244.860 45.000 ;
        RECT 241.480 43.770 241.650 44.770 ;
        RECT 245.030 43.770 245.200 44.770 ;
        RECT 241.820 43.540 244.860 43.710 ;
        RECT 245.535 43.040 257.145 45.500 ;
        RECT 240.510 42.305 257.145 43.040 ;
        RECT 240.510 39.845 241.085 42.305 ;
        RECT 241.820 41.635 244.860 41.805 ;
        RECT 241.480 40.575 241.650 41.575 ;
        RECT 245.030 40.575 245.200 41.575 ;
        RECT 241.820 40.345 244.860 40.515 ;
        RECT 245.535 39.845 257.145 42.305 ;
        RECT 240.510 39.110 257.145 39.845 ;
        RECT 240.510 36.650 241.085 39.110 ;
        RECT 241.820 38.440 244.860 38.610 ;
        RECT 241.480 37.380 241.650 38.380 ;
        RECT 245.030 37.380 245.200 38.380 ;
        RECT 241.820 37.150 244.860 37.320 ;
        RECT 245.535 36.650 257.145 39.110 ;
        RECT 240.510 35.915 257.145 36.650 ;
        RECT 240.510 33.455 241.085 35.915 ;
        RECT 241.820 35.245 244.860 35.415 ;
        RECT 241.480 34.185 241.650 35.185 ;
        RECT 245.030 34.185 245.200 35.185 ;
        RECT 241.820 33.955 244.860 34.125 ;
        RECT 245.535 33.455 257.145 35.915 ;
        RECT 240.510 32.720 257.145 33.455 ;
        RECT 240.510 30.260 241.085 32.720 ;
        RECT 241.820 32.050 244.860 32.220 ;
        RECT 241.480 30.990 241.650 31.990 ;
        RECT 245.030 30.990 245.200 31.990 ;
        RECT 241.820 30.760 244.860 30.930 ;
        RECT 245.535 30.260 257.145 32.720 ;
        RECT 240.510 29.525 257.145 30.260 ;
        RECT 240.510 27.065 241.085 29.525 ;
        RECT 241.820 28.855 244.860 29.025 ;
        RECT 241.480 27.795 241.650 28.795 ;
        RECT 245.030 27.795 245.200 28.795 ;
        RECT 241.820 27.565 244.860 27.735 ;
        RECT 245.535 27.065 257.145 29.525 ;
        RECT 240.510 26.330 257.145 27.065 ;
        RECT 240.510 23.870 241.085 26.330 ;
        RECT 241.820 25.660 242.860 25.830 ;
        RECT 241.480 24.600 241.650 25.600 ;
        RECT 243.030 24.600 243.200 25.600 ;
        RECT 241.820 24.370 242.860 24.540 ;
        RECT 243.640 23.870 257.145 26.330 ;
        RECT 240.510 23.140 257.145 23.870 ;
        RECT 240.510 20.765 241.085 23.140 ;
        RECT 241.835 22.470 242.875 22.640 ;
        RECT 241.495 21.410 241.665 22.410 ;
        RECT 243.045 21.410 243.215 22.410 ;
        RECT 241.835 21.180 242.875 21.350 ;
        RECT 243.640 20.765 257.145 23.140 ;
        RECT 257.450 20.860 257.800 23.020 ;
        RECT 240.510 20.445 257.145 20.765 ;
        RECT 258.075 20.445 258.585 50.450 ;
        RECT 258.930 47.810 259.280 49.970 ;
        RECT 258.930 20.860 259.280 23.020 ;
        RECT 259.560 20.445 260.070 50.450 ;
        RECT 260.410 47.810 260.760 49.970 ;
        RECT 260.410 20.860 260.760 23.020 ;
        RECT 261.230 20.445 261.780 50.450 ;
        RECT 240.510 19.435 261.780 20.445 ;
        RECT 240.565 19.385 261.780 19.435 ;
        RECT 257.085 19.375 261.780 19.385 ;
        RECT 193.680 18.870 224.415 18.940 ;
        RECT 193.745 18.860 224.415 18.870 ;
        RECT 193.745 18.830 224.400 18.860 ;
        RECT 145.575 18.410 174.475 18.435 ;
        RECT 145.760 18.395 174.415 18.410 ;
        RECT 86.095 16.890 87.530 16.895 ;
      LAYER met1 ;
        RECT 14.770 215.600 16.080 215.625 ;
        RECT 14.770 215.570 31.850 215.600 ;
        RECT 14.760 214.385 31.850 215.570 ;
        RECT 14.760 153.935 16.135 214.385 ;
        RECT 16.625 213.515 18.355 213.840 ;
        RECT 16.625 211.735 16.875 213.515 ;
        RECT 18.105 211.735 18.355 213.515 ;
        RECT 19.585 213.515 21.315 213.840 ;
        RECT 19.585 211.735 19.835 213.515 ;
        RECT 21.065 211.735 21.315 213.515 ;
        RECT 22.545 213.515 24.275 213.840 ;
        RECT 22.545 211.735 22.795 213.515 ;
        RECT 24.025 211.735 24.275 213.515 ;
        RECT 25.505 213.515 27.235 213.840 ;
        RECT 25.505 211.735 25.755 213.515 ;
        RECT 26.985 211.735 27.235 213.515 ;
        RECT 28.465 213.515 30.195 213.840 ;
        RECT 28.465 211.735 28.715 213.515 ;
        RECT 29.945 211.735 30.195 213.515 ;
        RECT 16.625 181.445 16.875 186.845 ;
        RECT 18.105 181.445 18.355 186.845 ;
        RECT 19.585 181.445 19.835 186.845 ;
        RECT 21.065 181.445 21.315 186.845 ;
        RECT 22.545 181.445 22.795 186.845 ;
        RECT 24.025 181.445 24.275 186.845 ;
        RECT 25.505 181.445 25.755 186.845 ;
        RECT 26.985 181.445 27.235 186.845 ;
        RECT 28.465 181.445 28.715 186.845 ;
        RECT 29.945 181.445 30.195 186.845 ;
        RECT 30.610 157.680 31.770 214.385 ;
        RECT 32.745 158.240 57.120 159.225 ;
        RECT 16.625 156.510 16.875 156.555 ;
        RECT 16.515 154.510 16.975 156.510 ;
        RECT 18.105 154.775 18.355 156.555 ;
        RECT 19.585 154.775 19.835 156.555 ;
        RECT 16.625 154.450 16.875 154.510 ;
        RECT 18.105 154.450 19.835 154.775 ;
        RECT 21.065 154.775 21.315 156.555 ;
        RECT 22.545 154.775 22.795 156.555 ;
        RECT 21.065 154.450 22.795 154.775 ;
        RECT 24.025 154.775 24.275 156.555 ;
        RECT 25.505 154.775 25.755 156.555 ;
        RECT 24.025 154.450 25.755 154.775 ;
        RECT 26.985 154.775 27.235 156.555 ;
        RECT 28.465 154.775 28.715 156.555 ;
        RECT 29.945 156.495 30.195 156.555 ;
        RECT 26.985 154.450 28.715 154.775 ;
        RECT 29.890 154.510 30.250 156.495 ;
        RECT 29.945 154.450 30.195 154.510 ;
        RECT 30.680 153.935 31.750 157.680 ;
        RECT 32.755 155.390 33.390 158.240 ;
        RECT 34.060 157.475 44.020 157.705 ;
        RECT 45.690 157.475 55.650 157.705 ;
        RECT 33.780 156.830 34.010 157.270 ;
        RECT 33.715 156.330 34.075 156.830 ;
        RECT 44.070 156.600 44.300 157.270 ;
        RECT 45.410 156.600 45.640 157.270 ;
        RECT 55.700 157.210 55.930 157.270 ;
        RECT 55.605 156.710 56.025 157.210 ;
        RECT 33.780 156.270 34.010 156.330 ;
        RECT 44.070 156.270 45.640 156.600 ;
        RECT 55.700 156.270 55.930 156.710 ;
        RECT 34.070 156.065 35.435 156.075 ;
        RECT 53.740 156.065 55.640 156.110 ;
        RECT 34.060 155.835 55.650 156.065 ;
        RECT 34.070 155.790 35.435 155.835 ;
        RECT 53.740 155.745 55.640 155.835 ;
        RECT 56.390 155.390 57.065 158.240 ;
        RECT 32.740 154.405 57.115 155.390 ;
        RECT 14.760 153.930 31.780 153.935 ;
        RECT 14.740 152.995 31.780 153.930 ;
        RECT 14.770 152.940 31.780 152.995 ;
        RECT 14.770 152.935 16.080 152.940 ;
        RECT 57.465 140.665 115.555 141.520 ;
        RECT 57.465 140.260 64.065 140.665 ;
        RECT 93.580 140.585 115.555 140.665 ;
        RECT 93.580 140.260 114.605 140.585 ;
        RECT 57.465 140.010 66.650 140.260 ;
        RECT 76.040 140.010 114.605 140.260 ;
        RECT 57.465 138.895 64.065 140.010 ;
        RECT 63.375 124.030 64.065 138.895 ;
        RECT 93.580 139.965 114.605 140.010 ;
        RECT 90.840 138.780 92.925 138.785 ;
        RECT 64.545 138.530 66.650 138.780 ;
        RECT 76.040 138.530 81.440 138.780 ;
        RECT 90.830 138.530 92.935 138.780 ;
        RECT 64.545 137.300 64.955 138.530 ;
        RECT 90.840 138.525 92.925 138.530 ;
        RECT 64.545 137.050 66.650 137.300 ;
        RECT 76.040 137.050 81.440 137.300 ;
        RECT 90.830 137.050 92.935 137.300 ;
        RECT 92.525 135.820 92.935 137.050 ;
        RECT 64.545 135.570 66.650 135.820 ;
        RECT 76.040 135.570 81.440 135.820 ;
        RECT 90.830 135.570 92.935 135.820 ;
        RECT 93.580 135.665 95.835 139.965 ;
        RECT 96.515 138.835 99.565 139.360 ;
        RECT 100.220 138.840 102.550 139.965 ;
        RECT 96.465 138.495 99.565 138.835 ;
        RECT 103.235 138.495 106.285 139.360 ;
        RECT 106.945 138.785 109.275 139.965 ;
        RECT 96.465 138.465 106.285 138.495 ;
        RECT 109.955 138.465 113.005 139.360 ;
        RECT 96.465 137.095 113.005 138.465 ;
        RECT 96.465 136.465 99.565 137.095 ;
        RECT 103.235 137.065 113.005 137.095 ;
        RECT 96.515 136.310 99.565 136.465 ;
        RECT 64.545 134.340 64.955 135.570 ;
        RECT 64.545 134.090 66.650 134.340 ;
        RECT 76.040 134.090 81.440 134.340 ;
        RECT 90.830 134.090 92.935 134.340 ;
        RECT 92.525 132.860 92.935 134.090 ;
        RECT 64.545 132.610 66.650 132.860 ;
        RECT 76.040 132.610 81.440 132.860 ;
        RECT 90.830 132.610 92.935 132.860 ;
        RECT 93.580 134.000 97.025 135.665 ;
        RECT 64.545 131.380 64.955 132.610 ;
        RECT 64.545 131.130 66.650 131.380 ;
        RECT 76.040 131.130 81.440 131.380 ;
        RECT 90.830 131.130 92.935 131.380 ;
        RECT 92.525 129.900 92.935 131.130 ;
        RECT 64.545 129.650 66.650 129.900 ;
        RECT 76.040 129.650 81.440 129.900 ;
        RECT 90.830 129.650 92.935 129.900 ;
        RECT 64.545 128.420 64.955 129.650 ;
        RECT 93.580 128.935 95.835 134.000 ;
        RECT 97.300 132.640 98.845 136.310 ;
        RECT 100.365 135.650 102.505 136.665 ;
        RECT 103.235 136.310 106.285 137.065 ;
        RECT 107.015 135.650 109.155 136.665 ;
        RECT 109.955 136.310 113.005 137.065 ;
        RECT 99.275 134.100 110.465 135.650 ;
        RECT 96.515 129.590 99.565 132.640 ;
        RECT 64.545 128.170 66.650 128.420 ;
        RECT 76.040 128.170 81.440 128.420 ;
        RECT 90.830 128.170 92.935 128.420 ;
        RECT 92.525 126.940 92.935 128.170 ;
        RECT 64.545 126.690 66.650 126.940 ;
        RECT 76.040 126.690 81.440 126.940 ;
        RECT 90.830 126.690 92.935 126.940 ;
        RECT 93.580 127.270 97.025 128.935 ;
        RECT 64.545 125.460 64.955 126.690 ;
        RECT 91.325 125.460 92.925 125.465 ;
        RECT 64.545 125.210 66.650 125.460 ;
        RECT 76.040 125.210 81.440 125.460 ;
        RECT 90.830 125.210 92.935 125.460 ;
        RECT 91.325 125.205 92.925 125.210 ;
        RECT 63.375 123.980 64.645 124.030 ;
        RECT 93.580 123.985 95.835 127.270 ;
        RECT 97.285 125.920 98.830 129.590 ;
        RECT 100.365 128.905 102.505 134.100 ;
        RECT 103.235 129.590 106.285 132.640 ;
        RECT 107.015 128.905 109.155 134.100 ;
        RECT 110.780 132.640 112.325 136.310 ;
        RECT 113.675 135.700 114.605 139.965 ;
        RECT 112.530 134.035 114.605 135.700 ;
        RECT 109.955 129.590 113.005 132.640 ;
        RECT 99.430 127.315 110.410 128.905 ;
        RECT 92.865 123.980 95.835 123.985 ;
        RECT 63.375 123.730 95.835 123.980 ;
        RECT 63.375 123.680 64.645 123.730 ;
        RECT 55.265 122.880 56.520 122.910 ;
        RECT 63.375 122.880 64.065 123.680 ;
        RECT 55.265 122.850 64.065 122.880 ;
        RECT 55.245 122.845 64.065 122.850 ;
        RECT 93.580 122.845 95.835 123.730 ;
        RECT 96.515 124.995 99.565 125.920 ;
        RECT 100.365 125.210 102.505 127.315 ;
        RECT 103.235 124.995 106.285 125.920 ;
        RECT 107.015 125.210 109.155 127.315 ;
        RECT 110.805 125.920 112.350 129.590 ;
        RECT 113.675 129.030 114.605 134.035 ;
        RECT 112.605 127.190 114.605 129.030 ;
        RECT 96.515 124.980 106.285 124.995 ;
        RECT 109.955 124.980 113.005 125.920 ;
        RECT 96.515 123.595 113.005 124.980 ;
        RECT 96.515 122.870 99.565 123.595 ;
        RECT 103.235 123.580 113.005 123.595 ;
        RECT 55.245 122.255 95.835 122.845 ;
        RECT 100.240 122.255 102.570 123.355 ;
        RECT 103.235 122.870 106.285 123.580 ;
        RECT 106.965 122.255 109.295 123.335 ;
        RECT 109.955 122.870 113.005 123.580 ;
        RECT 113.675 122.255 114.605 127.190 ;
        RECT 55.245 121.710 114.605 122.255 ;
        RECT 55.245 120.705 114.635 121.710 ;
        RECT 55.245 99.545 56.540 120.705 ;
        RECT 57.345 120.255 57.845 120.285 ;
        RECT 57.325 120.085 57.865 120.255 ;
        RECT 57.345 120.055 57.845 120.085 ;
        RECT 56.955 118.615 57.185 120.030 ;
        RECT 57.435 119.995 57.835 120.055 ;
        RECT 58.005 119.550 58.235 120.025 ;
        RECT 57.935 118.615 58.295 119.550 ;
        RECT 56.955 114.550 58.295 118.615 ;
        RECT 56.955 101.405 58.235 114.550 ;
        RECT 56.955 99.965 57.185 101.405 ;
        RECT 57.345 99.965 57.845 99.995 ;
        RECT 58.005 99.965 58.235 101.405 ;
        RECT 56.955 99.795 58.235 99.965 ;
        RECT 57.345 99.765 57.845 99.795 ;
        RECT 57.435 99.735 57.835 99.765 ;
        RECT 58.695 99.545 58.925 120.705 ;
        RECT 59.775 120.055 60.275 120.285 ;
        RECT 59.385 119.550 59.615 120.005 ;
        RECT 59.785 119.995 60.185 120.055 ;
        RECT 60.435 119.550 60.665 120.005 ;
        RECT 59.325 118.615 59.685 119.550 ;
        RECT 60.375 118.615 60.735 119.550 ;
        RECT 59.325 114.550 60.735 118.615 ;
        RECT 59.385 101.405 60.665 114.550 ;
        RECT 59.385 100.045 59.615 101.405 ;
        RECT 60.435 100.045 60.665 101.405 ;
        RECT 59.775 99.765 60.275 99.995 ;
        RECT 59.865 99.705 60.265 99.765 ;
        RECT 61.125 99.545 61.355 120.705 ;
        RECT 62.295 120.285 62.695 120.345 ;
        RECT 62.205 120.055 62.705 120.285 ;
        RECT 61.815 119.560 62.045 120.005 ;
        RECT 61.765 118.615 62.125 119.560 ;
        RECT 62.865 118.615 63.095 120.005 ;
        RECT 61.765 114.560 63.095 118.615 ;
        RECT 61.815 101.405 63.095 114.560 ;
        RECT 61.815 100.045 62.045 101.405 ;
        RECT 62.865 100.045 63.095 101.405 ;
        RECT 62.205 99.765 62.705 99.995 ;
        RECT 62.215 99.705 62.615 99.765 ;
        RECT 63.555 99.545 63.785 120.705 ;
        RECT 64.725 120.285 65.125 120.345 ;
        RECT 64.635 120.255 65.135 120.285 ;
        RECT 64.635 120.085 65.155 120.255 ;
        RECT 64.635 120.055 65.135 120.085 ;
        RECT 64.245 118.660 64.475 120.025 ;
        RECT 65.295 119.575 65.525 120.035 ;
        RECT 65.220 118.660 65.580 119.575 ;
        RECT 64.245 114.575 65.580 118.660 ;
        RECT 64.245 101.430 65.525 114.575 ;
        RECT 64.245 99.965 64.475 101.430 ;
        RECT 64.635 99.965 65.135 99.995 ;
        RECT 65.295 99.965 65.525 101.430 ;
        RECT 64.245 99.795 65.525 99.965 ;
        RECT 64.635 99.790 65.525 99.795 ;
        RECT 64.635 99.765 65.135 99.790 ;
        RECT 64.645 99.705 65.045 99.765 ;
        RECT 65.985 99.545 66.215 120.705 ;
        RECT 67.075 120.285 67.475 120.345 ;
        RECT 67.065 120.055 67.565 120.285 ;
        RECT 66.675 119.575 66.905 120.005 ;
        RECT 66.615 118.660 66.975 119.575 ;
        RECT 67.725 119.565 67.955 120.005 ;
        RECT 67.660 118.660 68.020 119.565 ;
        RECT 66.615 114.575 68.020 118.660 ;
        RECT 66.675 114.565 68.020 114.575 ;
        RECT 66.675 101.430 67.955 114.565 ;
        RECT 66.675 100.045 66.905 101.430 ;
        RECT 67.725 100.045 67.955 101.430 ;
        RECT 67.065 99.765 67.565 99.995 ;
        RECT 67.155 99.705 67.555 99.765 ;
        RECT 68.415 99.545 68.645 120.705 ;
        RECT 69.585 120.285 69.985 120.345 ;
        RECT 69.495 120.055 69.995 120.285 ;
        RECT 69.105 119.565 69.335 120.005 ;
        RECT 69.035 118.675 69.395 119.565 ;
        RECT 70.155 119.560 70.385 120.005 ;
        RECT 70.095 118.675 70.455 119.560 ;
        RECT 69.035 114.565 70.455 118.675 ;
        RECT 69.105 114.560 70.455 114.565 ;
        RECT 69.105 101.445 70.385 114.560 ;
        RECT 69.105 100.045 69.335 101.445 ;
        RECT 70.155 100.045 70.385 101.445 ;
        RECT 69.495 99.765 69.995 99.995 ;
        RECT 69.505 99.705 69.905 99.765 ;
        RECT 70.845 99.545 71.075 120.705 ;
        RECT 71.935 120.285 72.335 120.345 ;
        RECT 71.925 120.055 72.425 120.285 ;
        RECT 71.535 119.560 71.765 120.005 ;
        RECT 72.585 119.560 72.815 120.005 ;
        RECT 71.470 118.675 71.830 119.560 ;
        RECT 72.520 118.675 72.880 119.560 ;
        RECT 71.470 114.560 72.880 118.675 ;
        RECT 71.535 101.445 72.815 114.560 ;
        RECT 71.535 100.045 71.765 101.445 ;
        RECT 72.585 100.045 72.815 101.445 ;
        RECT 71.925 99.765 72.425 99.995 ;
        RECT 72.015 99.705 72.415 99.765 ;
        RECT 73.275 99.545 73.505 120.705 ;
        RECT 74.445 120.285 74.845 120.345 ;
        RECT 74.355 120.055 74.855 120.285 ;
        RECT 73.965 119.560 74.195 120.005 ;
        RECT 75.015 119.560 75.245 120.005 ;
        RECT 73.900 118.675 74.260 119.560 ;
        RECT 74.955 118.675 75.315 119.560 ;
        RECT 73.900 114.560 75.315 118.675 ;
        RECT 73.965 101.445 75.245 114.560 ;
        RECT 73.965 100.045 74.195 101.445 ;
        RECT 75.015 100.045 75.245 101.445 ;
        RECT 74.355 99.765 74.855 99.995 ;
        RECT 74.365 99.705 74.765 99.765 ;
        RECT 75.705 99.545 75.935 120.705 ;
        RECT 76.795 120.285 77.195 120.345 ;
        RECT 76.785 120.055 77.285 120.285 ;
        RECT 76.395 119.560 76.625 120.005 ;
        RECT 77.445 119.560 77.675 120.005 ;
        RECT 76.330 118.675 76.690 119.560 ;
        RECT 77.380 118.675 77.740 119.560 ;
        RECT 76.330 114.560 77.740 118.675 ;
        RECT 76.395 101.445 77.675 114.560 ;
        RECT 76.395 100.045 76.625 101.445 ;
        RECT 77.445 100.045 77.675 101.445 ;
        RECT 76.785 99.765 77.285 99.995 ;
        RECT 76.875 99.705 77.275 99.765 ;
        RECT 78.135 99.545 78.365 120.705 ;
        RECT 79.305 120.285 79.705 120.345 ;
        RECT 79.215 120.055 79.715 120.285 ;
        RECT 78.825 119.560 79.055 120.005 ;
        RECT 78.765 118.690 79.125 119.560 ;
        RECT 79.875 118.690 80.105 120.005 ;
        RECT 78.765 114.560 80.105 118.690 ;
        RECT 78.825 101.460 80.105 114.560 ;
        RECT 78.825 100.045 79.055 101.460 ;
        RECT 79.875 100.045 80.105 101.460 ;
        RECT 80.410 117.355 80.890 120.705 ;
        RECT 104.330 120.020 114.635 120.705 ;
        RECT 126.380 120.020 127.360 120.050 ;
        RECT 104.330 118.630 127.360 120.020 ;
        RECT 105.820 118.000 125.780 118.230 ;
        RECT 105.540 117.780 105.770 117.840 ;
        RECT 80.410 117.325 81.315 117.355 ;
        RECT 80.410 116.535 104.620 117.325 ;
        RECT 105.475 116.780 105.835 117.780 ;
        RECT 80.410 116.505 81.315 116.535 ;
        RECT 80.410 116.500 81.205 116.505 ;
        RECT 80.410 103.725 80.890 116.500 ;
        RECT 81.925 111.555 82.715 116.535 ;
        RECT 83.290 116.000 103.500 116.230 ;
        RECT 83.290 115.840 83.460 116.000 ;
        RECT 83.260 113.900 83.490 115.840 ;
        RECT 83.195 112.900 83.555 113.900 ;
        RECT 83.260 112.840 83.490 112.900 ;
        RECT 83.290 112.680 83.460 112.840 ;
        RECT 91.765 112.680 96.015 116.000 ;
        RECT 103.550 113.900 103.780 115.840 ;
        RECT 103.485 112.900 103.845 113.900 ;
        RECT 103.550 112.840 103.780 112.900 ;
        RECT 105.540 112.840 105.770 116.780 ;
        RECT 113.945 112.680 118.215 118.000 ;
        RECT 125.830 117.780 126.060 117.840 ;
        RECT 125.765 116.780 126.125 117.780 ;
        RECT 125.830 112.840 126.060 116.780 ;
        RECT 83.290 112.450 125.780 112.680 ;
        RECT 102.500 112.135 106.820 112.450 ;
        RECT 81.925 110.575 102.275 111.555 ;
        RECT 81.925 110.545 82.920 110.575 ;
        RECT 80.410 103.695 80.930 103.725 ;
        RECT 82.555 103.695 82.920 110.545 ;
        RECT 102.500 110.185 103.500 112.135 ;
        RECT 105.820 110.185 106.820 112.135 ;
        RECT 126.380 111.710 127.360 118.630 ;
        RECT 107.260 110.445 127.360 111.710 ;
        RECT 102.500 109.870 106.820 110.185 ;
        RECT 83.575 109.640 125.780 109.870 ;
        RECT 83.295 105.540 83.525 109.480 ;
        RECT 83.230 104.540 83.590 105.540 ;
        RECT 83.295 104.480 83.525 104.540 ;
        RECT 91.710 104.320 95.980 109.640 ;
        RECT 105.570 109.480 105.740 109.640 ;
        RECT 103.585 105.540 103.815 109.480 ;
        RECT 105.540 109.420 105.770 109.480 ;
        RECT 104.205 108.585 105.045 108.645 ;
        RECT 104.185 105.720 105.065 108.585 ;
        RECT 105.475 108.420 105.835 109.420 ;
        RECT 105.540 106.480 105.770 108.420 ;
        RECT 105.570 106.320 105.740 106.480 ;
        RECT 114.070 106.320 118.320 109.640 ;
        RECT 125.830 109.420 126.060 109.480 ;
        RECT 125.765 108.420 126.125 109.420 ;
        RECT 126.380 108.505 127.360 110.445 ;
        RECT 125.830 106.480 126.060 108.420 ;
        RECT 105.570 106.090 125.780 106.320 ;
        RECT 126.340 105.720 127.375 108.505 ;
        RECT 103.520 104.540 103.880 105.540 ;
        RECT 104.185 105.295 127.375 105.720 ;
        RECT 104.185 105.120 127.360 105.295 ;
        RECT 103.585 104.480 103.815 104.540 ;
        RECT 83.575 104.090 103.535 104.320 ;
        RECT 80.410 103.690 82.960 103.695 ;
        RECT 104.215 103.690 104.615 105.120 ;
        RECT 126.380 105.090 127.360 105.120 ;
        RECT 80.410 103.195 104.660 103.690 ;
        RECT 79.215 99.765 79.715 99.995 ;
        RECT 79.225 99.705 79.625 99.765 ;
        RECT 80.410 99.545 80.930 103.195 ;
        RECT 82.555 103.165 82.920 103.195 ;
        RECT 104.215 103.180 104.615 103.195 ;
        RECT 55.235 98.370 80.930 99.545 ;
        RECT 57.235 95.945 127.115 96.635 ;
        RECT 57.235 84.150 57.875 95.945 ;
        RECT 73.285 95.435 78.385 95.460 ;
        RECT 58.625 95.205 78.605 95.435 ;
        RECT 60.300 95.180 78.385 95.205 ;
        RECT 58.345 94.940 58.575 95.000 ;
        RECT 58.280 93.560 58.640 94.940 ;
        RECT 58.345 93.500 58.575 93.560 ;
        RECT 60.300 93.295 77.180 95.180 ;
        RECT 78.635 94.940 78.865 95.000 ;
        RECT 78.570 93.560 78.930 94.940 ;
        RECT 78.635 93.500 78.865 93.560 ;
        RECT 58.625 93.065 78.585 93.295 ;
        RECT 59.155 92.755 78.410 93.065 ;
        RECT 58.625 92.525 78.585 92.755 ;
        RECT 58.345 92.260 58.575 92.320 ;
        RECT 58.280 90.880 58.640 92.260 ;
        RECT 58.345 90.820 58.575 90.880 ;
        RECT 60.275 90.615 77.125 92.525 ;
        RECT 78.635 92.260 78.865 92.320 ;
        RECT 78.570 90.880 78.930 92.260 ;
        RECT 78.635 90.820 78.865 90.880 ;
        RECT 58.625 90.385 78.585 90.615 ;
        RECT 76.145 88.435 78.040 90.385 ;
        RECT 58.625 88.205 78.585 88.435 ;
        RECT 58.345 87.940 58.575 88.000 ;
        RECT 58.245 86.940 58.665 87.940 ;
        RECT 58.345 85.000 58.575 86.940 ;
        RECT 59.915 84.795 76.780 88.205 ;
        RECT 78.635 87.940 78.865 88.000 ;
        RECT 78.570 85.060 78.930 87.940 ;
        RECT 78.635 85.000 78.865 85.060 ;
        RECT 58.625 84.565 78.605 84.795 ;
        RECT 66.490 84.150 67.830 84.175 ;
        RECT 79.425 84.150 83.310 95.945 ;
        RECT 84.065 95.435 89.165 95.460 ;
        RECT 84.045 95.205 125.935 95.435 ;
        RECT 84.065 95.180 89.165 95.205 ;
        RECT 83.785 88.060 84.015 95.000 ;
        RECT 83.690 85.060 84.110 88.060 ;
        RECT 83.785 85.000 84.015 85.060 ;
        RECT 91.850 84.795 97.745 95.205 ;
        RECT 104.075 94.390 104.305 95.000 ;
        RECT 105.415 94.390 105.645 95.000 ;
        RECT 104.075 87.560 105.645 94.390 ;
        RECT 104.010 85.520 105.710 87.560 ;
        RECT 104.010 85.060 104.370 85.520 ;
        RECT 105.350 85.060 105.710 85.520 ;
        RECT 104.075 85.000 104.305 85.060 ;
        RECT 105.415 85.000 105.645 85.060 ;
        RECT 113.110 84.795 119.005 95.205 ;
        RECT 125.705 94.940 125.935 95.205 ;
        RECT 125.610 91.940 126.030 94.940 ;
        RECT 126.410 94.735 127.115 95.945 ;
        RECT 126.410 94.010 135.800 94.735 ;
        RECT 125.705 85.000 125.935 91.940 ;
        RECT 125.735 84.795 125.905 85.000 ;
        RECT 84.045 84.565 125.905 84.795 ;
        RECT 57.205 83.420 83.310 84.150 ;
        RECT 57.260 83.410 57.875 83.420 ;
        RECT 66.835 74.920 83.310 83.420 ;
        RECT 84.110 83.415 103.655 84.565 ;
        RECT 106.055 83.415 125.600 84.565 ;
        RECT 83.785 83.185 125.655 83.415 ;
        RECT 83.785 82.920 84.015 83.185 ;
        RECT 83.690 79.920 84.110 82.920 ;
        RECT 66.835 73.690 67.830 74.920 ;
        RECT 68.635 74.415 73.735 74.430 ;
        RECT 68.635 74.185 78.585 74.415 ;
        RECT 68.635 74.170 77.605 74.185 ;
        RECT 66.805 72.095 67.865 73.690 ;
        RECT 68.395 73.675 68.625 73.980 ;
        RECT 68.280 73.040 68.640 73.675 ;
        RECT 68.395 72.980 68.625 73.040 ;
        RECT 70.000 72.775 77.605 74.170 ;
        RECT 78.635 73.920 78.865 73.980 ;
        RECT 78.570 73.040 78.930 73.920 ;
        RECT 78.635 72.980 78.865 73.040 ;
        RECT 68.675 72.545 78.585 72.775 ;
        RECT 79.425 72.095 83.310 74.920 ;
        RECT 83.785 72.980 84.015 79.920 ;
        RECT 83.815 72.775 84.015 72.980 ;
        RECT 91.680 72.775 97.575 83.185 ;
        RECT 104.075 82.920 104.305 82.980 ;
        RECT 105.415 82.920 105.645 82.980 ;
        RECT 104.010 82.400 104.370 82.920 ;
        RECT 105.350 82.400 105.710 82.920 ;
        RECT 104.010 80.420 105.710 82.400 ;
        RECT 104.075 73.995 105.645 80.420 ;
        RECT 104.010 73.470 105.710 73.995 ;
        RECT 104.010 73.040 104.370 73.470 ;
        RECT 105.350 73.040 105.710 73.470 ;
        RECT 104.075 72.980 104.305 73.040 ;
        RECT 105.415 72.980 105.645 73.040 ;
        RECT 113.195 72.775 119.090 83.185 ;
        RECT 125.705 76.040 125.935 82.980 ;
        RECT 125.610 73.635 126.030 76.040 ;
        RECT 125.705 72.980 125.935 73.635 ;
        RECT 83.815 72.545 125.655 72.775 ;
        RECT 126.410 72.095 130.205 94.010 ;
        RECT 131.090 93.615 131.570 93.645 ;
        RECT 131.080 93.385 131.580 93.615 ;
        RECT 133.550 93.405 134.150 93.725 ;
        RECT 133.600 93.385 134.100 93.405 ;
        RECT 130.645 90.090 130.875 93.335 ;
        RECT 131.785 93.245 132.015 93.335 ;
        RECT 131.710 90.090 132.090 93.245 ;
        RECT 130.645 88.245 132.090 90.090 ;
        RECT 133.165 90.090 133.395 93.335 ;
        RECT 134.305 93.035 134.535 93.335 ;
        RECT 134.230 90.090 134.610 93.035 ;
        RECT 130.645 77.105 132.015 88.245 ;
        RECT 130.645 73.375 130.875 77.105 ;
        RECT 131.785 73.375 132.015 77.105 ;
        RECT 133.165 88.035 134.610 90.090 ;
        RECT 133.165 77.105 134.535 88.035 ;
        RECT 133.165 73.375 133.395 77.105 ;
        RECT 134.305 73.375 134.535 77.105 ;
        RECT 131.080 73.095 131.580 73.325 ;
        RECT 133.600 73.095 134.100 73.325 ;
        RECT 131.090 73.065 131.570 73.095 ;
        RECT 133.610 73.065 134.090 73.095 ;
        RECT 134.995 72.095 135.800 94.010 ;
        RECT 259.640 92.950 272.635 93.710 ;
        RECT 243.610 90.800 246.665 90.830 ;
        RECT 240.490 90.145 246.665 90.800 ;
        RECT 240.535 87.750 241.045 90.145 ;
        RECT 242.280 89.760 242.780 89.825 ;
        RECT 241.840 89.530 242.840 89.760 ;
        RECT 241.450 89.030 241.680 89.480 ;
        RECT 242.280 89.465 242.780 89.530 ;
        RECT 241.435 88.530 241.695 89.030 ;
        RECT 241.450 88.520 241.680 88.530 ;
        RECT 242.280 88.470 242.780 88.535 ;
        RECT 243.000 88.520 243.230 89.480 ;
        RECT 241.840 88.240 242.840 88.470 ;
        RECT 242.280 88.175 242.780 88.240 ;
        RECT 243.610 87.750 246.665 90.145 ;
        RECT 259.670 89.515 260.180 92.950 ;
        RECT 260.635 89.880 262.680 92.690 ;
        RECT 269.630 89.880 271.675 92.690 ;
        RECT 264.660 89.515 265.170 89.545 ;
        RECT 271.895 89.515 272.605 92.950 ;
        RECT 240.535 87.070 246.665 87.750 ;
        RECT 240.535 84.625 241.045 87.070 ;
        RECT 243.610 87.050 246.665 87.070 ;
        RECT 259.640 88.675 272.605 89.515 ;
        RECT 259.640 87.480 265.170 88.675 ;
        RECT 265.630 88.215 267.145 88.275 ;
        RECT 270.910 88.215 271.610 88.280 ;
        RECT 265.570 87.965 267.675 88.215 ;
        RECT 269.565 87.965 271.670 88.215 ;
        RECT 265.630 87.900 267.145 87.965 ;
        RECT 270.910 87.900 271.610 87.965 ;
        RECT 271.895 87.480 272.605 88.675 ;
        RECT 259.640 87.050 272.605 87.480 ;
        RECT 243.610 86.655 272.605 87.050 ;
        RECT 242.280 86.565 242.780 86.630 ;
        RECT 241.840 86.335 242.840 86.565 ;
        RECT 241.450 85.835 241.680 86.285 ;
        RECT 242.280 86.270 242.780 86.335 ;
        RECT 241.435 85.335 241.695 85.835 ;
        RECT 241.450 85.325 241.680 85.335 ;
        RECT 242.280 85.275 242.780 85.340 ;
        RECT 243.000 85.325 243.230 86.285 ;
        RECT 243.610 85.475 246.660 86.655 ;
        RECT 264.640 86.635 272.605 86.655 ;
        RECT 264.660 86.605 265.170 86.635 ;
        RECT 247.145 86.140 248.145 86.210 ;
        RECT 270.125 86.140 271.125 86.210 ;
        RECT 247.035 85.890 249.140 86.140 ;
        RECT 269.030 85.890 271.135 86.140 ;
        RECT 247.145 85.850 248.145 85.890 ;
        RECT 270.125 85.850 271.125 85.890 ;
        RECT 271.665 85.500 272.605 86.635 ;
        RECT 252.530 85.475 253.635 85.500 ;
        RECT 243.610 85.450 253.635 85.475 ;
        RECT 271.515 85.470 272.605 85.500 ;
        RECT 256.140 85.450 272.605 85.470 ;
        RECT 241.840 85.045 242.840 85.275 ;
        RECT 242.280 84.980 242.780 85.045 ;
        RECT 243.610 84.805 272.605 85.450 ;
        RECT 243.610 84.625 272.635 84.805 ;
        RECT 240.535 83.815 272.635 84.625 ;
        RECT 240.535 81.240 241.045 83.815 ;
        RECT 246.780 83.370 251.780 83.435 ;
        RECT 241.840 83.140 251.840 83.370 ;
        RECT 241.450 82.640 241.680 83.090 ;
        RECT 246.780 83.075 251.780 83.140 ;
        RECT 241.435 82.140 241.695 82.640 ;
        RECT 241.450 82.130 241.680 82.140 ;
        RECT 246.780 82.080 251.780 82.145 ;
        RECT 252.000 82.130 252.230 83.090 ;
        RECT 241.840 81.850 251.840 82.080 ;
        RECT 246.780 81.785 251.780 81.850 ;
        RECT 252.530 81.240 272.635 83.815 ;
        RECT 240.535 80.725 272.635 81.240 ;
        RECT 229.620 78.120 234.745 78.140 ;
        RECT 229.560 77.995 234.805 78.120 ;
        RECT 229.560 77.440 234.855 77.995 ;
        RECT 229.620 77.420 234.855 77.440 ;
        RECT 66.805 69.690 135.800 72.095 ;
        RECT 229.655 74.970 230.430 77.420 ;
        RECT 232.915 76.980 233.315 77.045 ;
        RECT 231.375 76.750 233.375 76.980 ;
        RECT 230.940 75.740 231.170 76.700 ;
        RECT 232.915 76.685 233.315 76.750 ;
        RECT 233.580 76.250 233.810 76.700 ;
        RECT 231.435 75.690 231.835 75.755 ;
        RECT 233.565 75.750 233.825 76.250 ;
        RECT 233.580 75.740 233.810 75.750 ;
        RECT 231.375 75.460 233.375 75.690 ;
        RECT 231.435 75.395 231.835 75.460 ;
        RECT 234.205 74.970 234.855 77.420 ;
        RECT 229.655 74.325 234.855 74.970 ;
        RECT 229.655 71.790 230.430 74.325 ;
        RECT 232.915 73.785 233.315 73.850 ;
        RECT 231.375 73.555 233.375 73.785 ;
        RECT 230.940 72.545 231.170 73.505 ;
        RECT 232.915 73.490 233.315 73.555 ;
        RECT 233.580 73.055 233.810 73.505 ;
        RECT 231.435 72.495 231.835 72.560 ;
        RECT 233.565 72.555 233.825 73.055 ;
        RECT 233.580 72.545 233.810 72.555 ;
        RECT 231.375 72.265 233.375 72.495 ;
        RECT 231.435 72.200 231.835 72.265 ;
        RECT 234.205 71.790 234.855 74.325 ;
        RECT 229.655 71.145 234.855 71.790 ;
        RECT 192.915 67.515 224.630 68.900 ;
        RECT 229.655 68.585 230.430 71.145 ;
        RECT 232.915 70.590 233.315 70.655 ;
        RECT 231.375 70.360 233.375 70.590 ;
        RECT 230.940 69.350 231.170 70.310 ;
        RECT 232.915 70.295 233.315 70.360 ;
        RECT 233.580 69.860 233.810 70.310 ;
        RECT 231.435 69.300 231.835 69.365 ;
        RECT 233.565 69.360 233.825 69.860 ;
        RECT 233.580 69.350 233.810 69.360 ;
        RECT 231.375 69.070 233.375 69.300 ;
        RECT 231.435 69.005 231.835 69.070 ;
        RECT 234.205 68.585 234.855 71.145 ;
        RECT 229.655 67.940 234.855 68.585 ;
        RECT 72.220 59.945 72.875 59.960 ;
        RECT 72.220 59.900 77.565 59.945 ;
        RECT 48.305 57.905 63.315 59.490 ;
        RECT 72.200 59.330 77.565 59.900 ;
        RECT 38.535 55.215 39.310 55.245 ;
        RECT 48.315 55.215 49.390 57.905 ;
        RECT 49.980 57.160 59.990 57.390 ;
        RECT 49.635 56.015 49.995 57.015 ;
        RECT 49.700 55.955 49.930 56.015 ;
        RECT 51.545 55.760 58.290 57.160 ;
        RECT 60.040 56.895 60.270 56.955 ;
        RECT 59.925 56.015 60.285 56.895 ;
        RECT 60.040 55.955 60.270 56.015 ;
        RECT 49.990 55.750 58.290 55.760 ;
        RECT 49.980 55.520 59.990 55.750 ;
        RECT 49.990 55.500 53.635 55.520 ;
        RECT 60.735 55.215 63.310 57.905 ;
        RECT 72.200 56.350 72.895 59.330 ;
        RECT 73.425 58.860 73.885 59.090 ;
        RECT 74.215 58.860 74.675 59.090 ;
        RECT 75.005 58.860 75.465 59.090 ;
        RECT 75.795 58.860 76.255 59.090 ;
        RECT 73.145 58.215 73.375 58.655 ;
        RECT 73.080 57.715 73.440 58.215 ;
        RECT 73.145 57.655 73.375 57.715 ;
        RECT 73.585 57.450 73.765 58.860 ;
        RECT 74.335 58.855 74.515 58.860 ;
        RECT 73.935 57.655 74.165 58.655 ;
        RECT 74.340 57.455 74.505 58.855 ;
        RECT 74.725 58.595 74.955 58.655 ;
        RECT 74.660 58.095 75.020 58.595 ;
        RECT 74.725 57.655 74.955 58.095 ;
        RECT 74.335 57.450 74.515 57.455 ;
        RECT 75.160 57.450 75.340 58.860 ;
        RECT 75.515 57.655 75.745 58.655 ;
        RECT 75.920 57.450 76.100 58.860 ;
        RECT 76.305 58.215 76.535 58.655 ;
        RECT 76.240 57.715 76.600 58.215 ;
        RECT 76.305 57.655 76.535 57.715 ;
        RECT 73.425 57.220 73.885 57.450 ;
        RECT 74.215 57.220 74.675 57.450 ;
        RECT 75.005 57.220 75.465 57.450 ;
        RECT 75.795 57.220 76.255 57.450 ;
        RECT 72.220 56.290 72.875 56.350 ;
        RECT 38.535 55.185 63.310 55.215 ;
        RECT 38.495 54.095 63.310 55.185 ;
        RECT 73.425 56.075 73.675 57.220 ;
        RECT 73.425 55.805 74.075 56.075 ;
        RECT 73.425 54.895 73.675 55.805 ;
        RECT 38.495 51.310 39.330 54.095 ;
        RECT 39.980 53.345 59.940 53.575 ;
        RECT 39.700 53.080 39.930 53.140 ;
        RECT 38.535 50.280 39.310 51.310 ;
        RECT 39.605 51.200 39.995 53.080 ;
        RECT 39.700 51.140 39.930 51.200 ;
        RECT 44.490 50.935 56.735 53.345 ;
        RECT 59.990 53.080 60.220 53.140 ;
        RECT 59.925 51.200 60.285 53.080 ;
        RECT 59.990 51.140 60.220 51.200 ;
        RECT 39.980 50.705 59.940 50.935 ;
        RECT 39.990 50.655 45.090 50.705 ;
        RECT 60.735 50.280 63.310 54.095 ;
        RECT 70.555 54.645 73.675 54.895 ;
        RECT 69.185 53.820 69.590 53.880 ;
        RECT 69.165 50.795 69.610 53.820 ;
        RECT 70.555 52.970 70.805 54.645 ;
        RECT 74.215 54.405 74.465 57.220 ;
        RECT 75.005 55.460 75.255 57.220 ;
        RECT 74.610 55.190 75.255 55.460 ;
        RECT 73.335 54.155 74.465 54.405 ;
        RECT 75.005 54.405 75.255 55.190 ;
        RECT 75.795 54.895 76.045 57.220 ;
        RECT 76.825 56.420 77.565 59.330 ;
        RECT 192.930 57.165 194.570 67.515 ;
        RECT 195.240 67.060 195.850 67.110 ;
        RECT 207.285 67.060 207.850 67.090 ;
        RECT 195.230 66.830 207.850 67.060 ;
        RECT 76.845 56.360 77.545 56.420 ;
        RECT 165.370 55.890 194.570 57.165 ;
        RECT 75.795 54.645 78.935 54.895 ;
        RECT 75.005 54.155 76.155 54.405 ;
        RECT 70.345 52.740 70.805 52.970 ;
        RECT 70.065 52.520 70.295 52.580 ;
        RECT 70.000 52.120 70.360 52.520 ;
        RECT 70.065 51.580 70.295 52.120 ;
        RECT 70.855 52.040 71.085 52.580 ;
        RECT 70.790 51.640 71.150 52.040 ;
        RECT 70.855 51.580 71.085 51.640 ;
        RECT 70.345 51.190 70.805 51.420 ;
        RECT 71.595 50.795 72.280 53.880 ;
        RECT 73.335 52.970 73.585 54.155 ;
        RECT 73.125 52.740 73.585 52.970 ;
        RECT 72.845 52.040 73.075 52.580 ;
        RECT 73.635 52.520 73.865 52.580 ;
        RECT 73.570 52.120 73.930 52.520 ;
        RECT 72.780 51.640 73.140 52.040 ;
        RECT 72.845 51.580 73.075 51.640 ;
        RECT 73.635 51.580 73.865 52.120 ;
        RECT 73.125 51.190 73.585 51.420 ;
        RECT 73.135 51.110 73.575 51.190 ;
        RECT 74.380 50.795 75.065 53.895 ;
        RECT 75.905 52.970 76.155 54.155 ;
        RECT 75.905 52.740 76.365 52.970 ;
        RECT 75.625 52.520 75.855 52.580 ;
        RECT 75.560 52.120 75.920 52.520 ;
        RECT 75.625 51.580 75.855 52.120 ;
        RECT 76.415 52.040 76.645 52.580 ;
        RECT 76.350 51.640 76.710 52.040 ;
        RECT 76.415 51.580 76.645 51.640 ;
        RECT 75.905 51.190 76.365 51.420 ;
        RECT 77.200 50.795 77.885 53.855 ;
        RECT 78.685 52.970 78.935 54.645 ;
        RECT 79.900 53.830 80.280 53.890 ;
        RECT 78.685 52.740 79.145 52.970 ;
        RECT 78.405 52.040 78.635 52.580 ;
        RECT 79.195 52.520 79.425 52.580 ;
        RECT 79.130 52.120 79.490 52.520 ;
        RECT 78.340 51.640 78.700 52.040 ;
        RECT 78.405 51.580 78.635 51.640 ;
        RECT 79.195 51.580 79.425 52.120 ;
        RECT 78.685 51.190 79.145 51.420 ;
        RECT 78.695 51.110 79.135 51.190 ;
        RECT 79.880 50.795 80.300 53.830 ;
        RECT 161.285 51.585 162.005 51.645 ;
        RECT 165.380 51.585 166.255 55.890 ;
        RECT 167.060 55.400 167.680 55.465 ;
        RECT 167.050 55.170 179.620 55.400 ;
        RECT 145.445 51.305 146.585 51.380 ;
        RECT 38.535 50.120 63.310 50.280 ;
        RECT 69.155 50.165 80.300 50.795 ;
        RECT 86.235 50.550 87.240 50.580 ;
        RECT 86.235 50.465 92.790 50.550 ;
        RECT 38.515 49.540 63.310 50.120 ;
        RECT 38.535 49.370 63.310 49.540 ;
        RECT 86.235 49.775 130.265 50.465 ;
        RECT 145.415 50.190 159.315 51.305 ;
        RECT 161.250 50.545 166.255 51.585 ;
        RECT 38.535 49.315 63.295 49.370 ;
        RECT 38.535 49.285 39.720 49.315 ;
        RECT 38.555 39.725 39.720 49.285 ;
        RECT 40.540 48.415 42.900 48.645 ;
        RECT 45.220 48.415 47.580 48.645 ;
        RECT 40.260 48.150 40.490 48.210 ;
        RECT 40.165 46.975 40.585 48.150 ;
        RECT 40.260 45.710 40.490 46.975 ;
        RECT 41.195 45.505 42.155 48.415 ;
        RECT 42.950 46.300 43.180 48.210 ;
        RECT 43.775 46.300 44.340 46.310 ;
        RECT 44.940 46.300 45.170 48.210 ;
        RECT 42.950 45.710 45.170 46.300 ;
        RECT 40.540 45.275 42.900 45.505 ;
        RECT 40.540 44.930 41.040 45.275 ;
        RECT 43.775 45.190 44.340 45.710 ;
        RECT 45.930 45.505 46.890 48.415 ;
        RECT 47.630 46.950 47.860 48.210 ;
        RECT 47.535 45.770 47.955 46.950 ;
        RECT 47.630 45.710 47.860 45.770 ;
        RECT 45.220 45.305 47.580 45.505 ;
        RECT 45.220 45.275 47.610 45.305 ;
        RECT 40.490 44.430 41.090 44.930 ;
        RECT 42.350 43.680 42.950 44.180 ;
        RECT 42.400 43.435 42.900 43.680 ;
        RECT 40.540 43.205 42.900 43.435 ;
        RECT 40.260 41.740 40.490 43.000 ;
        RECT 40.165 40.560 40.585 41.740 ;
        RECT 40.260 40.500 40.490 40.560 ;
        RECT 41.195 40.295 42.155 43.205 ;
        RECT 43.795 43.000 44.295 45.190 ;
        RECT 45.170 44.430 45.770 44.930 ;
        RECT 45.220 43.435 45.720 44.430 ;
        RECT 47.110 44.180 47.610 45.275 ;
        RECT 47.060 43.680 47.660 44.180 ;
        RECT 45.220 43.205 47.580 43.435 ;
        RECT 42.950 42.410 45.170 43.000 ;
        RECT 42.950 40.500 43.180 42.410 ;
        RECT 44.940 40.500 45.170 42.410 ;
        RECT 45.905 40.295 46.865 43.205 ;
        RECT 47.630 42.940 47.860 43.000 ;
        RECT 47.535 41.765 47.955 42.940 ;
        RECT 47.630 40.500 47.860 41.765 ;
        RECT 40.540 40.065 42.900 40.295 ;
        RECT 45.220 40.065 47.580 40.295 ;
        RECT 48.250 39.725 49.125 49.315 ;
        RECT 38.555 39.145 49.225 39.725 ;
        RECT 53.375 39.685 54.165 49.315 ;
        RECT 60.755 49.310 63.295 49.315 ;
        RECT 54.870 48.505 57.230 48.735 ;
        RECT 59.530 48.505 62.140 48.735 ;
        RECT 54.590 46.860 54.820 48.300 ;
        RECT 54.495 45.860 54.915 46.860 ;
        RECT 54.590 45.800 54.820 45.860 ;
        RECT 55.330 45.595 56.585 48.505 ;
        RECT 57.280 48.240 57.510 48.300 ;
        RECT 59.250 48.240 59.480 48.300 ;
        RECT 57.215 47.240 57.575 48.240 ;
        RECT 59.185 47.240 59.545 48.240 ;
        RECT 57.280 45.800 57.510 47.240 ;
        RECT 59.250 45.800 59.480 47.240 ;
        RECT 60.195 45.595 61.235 48.505 ;
        RECT 61.970 48.300 62.140 48.505 ;
        RECT 61.940 48.240 62.170 48.300 ;
        RECT 61.845 47.240 62.265 48.240 ;
        RECT 61.940 45.800 62.170 47.240 ;
        RECT 61.970 45.595 62.140 45.800 ;
        RECT 54.870 45.565 57.230 45.595 ;
        RECT 59.530 45.565 62.140 45.595 ;
        RECT 54.870 45.395 62.140 45.565 ;
        RECT 54.870 45.365 57.230 45.395 ;
        RECT 56.605 43.310 57.230 45.365 ;
        RECT 54.620 43.280 57.230 43.310 ;
        RECT 59.530 45.365 62.140 45.395 ;
        RECT 59.530 43.310 60.155 45.365 ;
        RECT 59.530 43.280 61.890 43.310 ;
        RECT 54.620 43.110 61.890 43.280 ;
        RECT 54.620 43.080 57.230 43.110 ;
        RECT 59.530 43.080 61.890 43.110 ;
        RECT 54.620 42.875 54.790 43.080 ;
        RECT 54.590 42.815 54.820 42.875 ;
        RECT 54.495 41.815 54.915 42.815 ;
        RECT 54.590 40.375 54.820 41.815 ;
        RECT 54.620 40.170 54.790 40.375 ;
        RECT 55.545 40.170 56.585 43.080 ;
        RECT 57.280 42.815 57.510 42.875 ;
        RECT 59.250 42.815 59.480 42.875 ;
        RECT 57.215 41.815 57.575 42.815 ;
        RECT 59.185 41.815 59.545 42.815 ;
        RECT 57.280 40.375 57.510 41.815 ;
        RECT 59.250 40.375 59.480 41.815 ;
        RECT 60.130 40.170 61.170 43.080 ;
        RECT 61.940 41.435 62.170 42.875 ;
        RECT 61.845 40.435 62.265 41.435 ;
        RECT 61.940 40.375 62.170 40.435 ;
        RECT 54.620 39.940 57.230 40.170 ;
        RECT 59.530 39.940 61.890 40.170 ;
        RECT 62.590 39.685 63.295 49.310 ;
        RECT 38.555 39.115 39.720 39.145 ;
        RECT 53.375 39.045 63.295 39.685 ;
        RECT 53.395 38.995 63.295 39.045 ;
        RECT 53.395 38.985 54.145 38.995 ;
        RECT 62.590 38.980 63.295 38.995 ;
        RECT 62.610 38.920 63.275 38.980 ;
        RECT 51.950 38.590 52.340 38.650 ;
        RECT 51.930 38.570 52.360 38.590 ;
        RECT 35.895 38.550 52.360 38.570 ;
        RECT 35.810 38.500 52.360 38.550 ;
        RECT 35.810 38.490 63.375 38.500 ;
        RECT 35.790 38.130 63.375 38.490 ;
        RECT 35.790 38.110 52.360 38.130 ;
        RECT 35.790 35.415 36.290 38.110 ;
        RECT 36.940 37.695 42.900 37.725 ;
        RECT 45.220 37.695 51.180 37.725 ;
        RECT 36.690 37.525 51.180 37.695 ;
        RECT 36.690 37.495 42.900 37.525 ;
        RECT 45.220 37.495 51.180 37.525 ;
        RECT 36.690 37.335 36.860 37.495 ;
        RECT 36.660 37.275 36.890 37.335 ;
        RECT 42.950 37.275 43.180 37.335 ;
        RECT 44.940 37.275 45.170 37.335 ;
        RECT 36.565 36.955 36.985 37.275 ;
        RECT 36.660 36.335 36.890 36.955 ;
        RECT 42.885 36.775 43.245 37.275 ;
        RECT 44.875 36.775 45.235 37.275 ;
        RECT 42.950 36.335 43.180 36.775 ;
        RECT 44.940 36.335 45.170 36.775 ;
        RECT 51.230 36.715 51.460 37.335 ;
        RECT 51.135 36.395 51.555 36.715 ;
        RECT 51.230 36.335 51.460 36.395 ;
        RECT 36.685 36.175 36.860 36.335 ;
        RECT 36.685 36.145 42.900 36.175 ;
        RECT 45.220 36.145 51.180 36.175 ;
        RECT 36.685 35.975 51.180 36.145 ;
        RECT 36.685 35.945 42.900 35.975 ;
        RECT 45.220 35.945 51.180 35.975 ;
        RECT 51.930 35.415 52.360 38.110 ;
        RECT 35.790 35.345 52.360 35.415 ;
        RECT 53.435 35.345 54.220 38.130 ;
        RECT 54.870 37.495 57.030 37.725 ;
        RECT 54.590 37.275 54.820 37.335 ;
        RECT 54.495 36.775 54.915 37.275 ;
        RECT 57.080 36.895 57.310 37.335 ;
        RECT 54.590 36.335 54.820 36.775 ;
        RECT 57.015 36.395 57.375 36.895 ;
        RECT 57.080 36.335 57.310 36.395 ;
        RECT 54.880 36.175 55.780 36.195 ;
        RECT 54.870 35.945 57.030 36.175 ;
        RECT 54.880 35.875 55.780 35.945 ;
        RECT 57.835 35.345 58.900 38.130 ;
        RECT 59.730 37.500 61.890 37.730 ;
        RECT 59.450 37.280 59.680 37.340 ;
        RECT 61.940 37.280 62.170 37.340 ;
        RECT 59.385 36.780 59.745 37.280 ;
        RECT 61.845 36.780 62.265 37.280 ;
        RECT 59.450 36.340 59.680 36.780 ;
        RECT 61.940 36.340 62.170 36.780 ;
        RECT 59.740 36.180 60.640 36.205 ;
        RECT 59.730 35.950 61.890 36.180 ;
        RECT 59.740 35.885 60.640 35.950 ;
        RECT 62.640 35.345 63.365 38.130 ;
        RECT 35.790 34.975 63.435 35.345 ;
        RECT 35.790 34.655 52.360 34.975 ;
        RECT 35.790 31.845 36.290 34.655 ;
        RECT 36.690 34.115 42.900 34.145 ;
        RECT 45.220 34.115 51.180 34.145 ;
        RECT 36.690 33.945 51.180 34.115 ;
        RECT 36.690 33.915 42.900 33.945 ;
        RECT 45.220 33.915 51.180 33.945 ;
        RECT 36.690 33.755 36.860 33.915 ;
        RECT 36.660 33.695 36.890 33.755 ;
        RECT 36.565 33.375 36.985 33.695 ;
        RECT 36.660 32.755 36.890 33.375 ;
        RECT 42.950 33.315 43.180 33.755 ;
        RECT 44.940 33.315 45.170 33.755 ;
        RECT 42.885 32.815 43.245 33.315 ;
        RECT 44.875 32.815 45.235 33.315 ;
        RECT 51.230 33.080 51.460 33.755 ;
        RECT 42.950 32.755 43.180 32.815 ;
        RECT 44.940 32.755 45.170 32.815 ;
        RECT 51.135 32.760 51.555 33.080 ;
        RECT 51.230 32.755 51.460 32.760 ;
        RECT 36.690 32.595 36.860 32.755 ;
        RECT 36.690 32.565 42.900 32.595 ;
        RECT 45.220 32.565 51.180 32.595 ;
        RECT 36.690 32.395 51.180 32.565 ;
        RECT 36.690 32.365 42.900 32.395 ;
        RECT 45.220 32.365 51.180 32.395 ;
        RECT 51.930 31.845 52.360 34.655 ;
        RECT 35.790 31.085 52.360 31.845 ;
        RECT 35.790 28.190 36.290 31.085 ;
        RECT 36.940 30.535 42.900 30.565 ;
        RECT 45.220 30.535 51.430 30.565 ;
        RECT 36.940 30.365 51.430 30.535 ;
        RECT 36.940 30.335 42.900 30.365 ;
        RECT 45.220 30.335 51.430 30.365 ;
        RECT 51.260 30.175 51.430 30.335 ;
        RECT 36.660 30.115 36.890 30.175 ;
        RECT 36.565 29.795 36.985 30.115 ;
        RECT 36.660 29.175 36.890 29.795 ;
        RECT 42.950 29.735 43.180 30.175 ;
        RECT 44.940 29.735 45.170 30.175 ;
        RECT 51.230 30.115 51.460 30.175 ;
        RECT 51.135 29.795 51.555 30.115 ;
        RECT 42.885 29.235 43.245 29.735 ;
        RECT 44.875 29.235 45.235 29.735 ;
        RECT 42.950 29.175 43.180 29.235 ;
        RECT 44.940 29.175 45.170 29.235 ;
        RECT 51.230 29.175 51.460 29.795 ;
        RECT 51.260 29.015 51.430 29.175 ;
        RECT 36.940 28.985 42.900 29.015 ;
        RECT 45.220 28.985 51.430 29.015 ;
        RECT 36.940 28.815 51.430 28.985 ;
        RECT 36.940 28.785 42.900 28.815 ;
        RECT 45.220 28.785 51.430 28.815 ;
        RECT 51.930 28.190 52.360 31.085 ;
        RECT 35.790 27.430 52.360 28.190 ;
        RECT 35.790 24.705 36.290 27.430 ;
        RECT 36.940 26.955 42.900 26.985 ;
        RECT 45.220 26.955 51.430 26.985 ;
        RECT 36.940 26.785 51.430 26.955 ;
        RECT 36.940 26.755 42.900 26.785 ;
        RECT 45.220 26.755 51.430 26.785 ;
        RECT 51.260 26.595 51.430 26.755 ;
        RECT 36.660 25.975 36.890 26.595 ;
        RECT 42.950 26.155 43.180 26.595 ;
        RECT 44.940 26.155 45.170 26.595 ;
        RECT 51.230 26.535 51.460 26.595 ;
        RECT 51.135 26.215 51.555 26.535 ;
        RECT 36.565 25.655 36.985 25.975 ;
        RECT 42.885 25.655 43.245 26.155 ;
        RECT 44.875 25.655 45.235 26.155 ;
        RECT 36.660 25.595 36.890 25.655 ;
        RECT 42.950 25.595 43.180 25.655 ;
        RECT 44.940 25.595 45.170 25.655 ;
        RECT 51.230 25.595 51.460 26.215 ;
        RECT 51.260 25.435 51.430 25.595 ;
        RECT 36.940 25.405 42.900 25.435 ;
        RECT 45.220 25.405 51.430 25.435 ;
        RECT 36.940 25.235 51.430 25.405 ;
        RECT 36.940 25.205 42.900 25.235 ;
        RECT 45.220 25.205 51.430 25.235 ;
        RECT 51.930 24.705 52.360 27.430 ;
        RECT 35.790 23.990 52.360 24.705 ;
        RECT 35.810 23.945 52.360 23.990 ;
        RECT 35.810 23.930 36.270 23.945 ;
        RECT 51.930 23.940 52.360 23.945 ;
        RECT 86.235 31.265 91.800 49.775 ;
        RECT 94.035 49.690 130.265 49.775 ;
        RECT 104.050 49.205 130.265 49.690 ;
        RECT 100.975 49.060 102.975 49.125 ;
        RECT 92.645 48.830 103.425 49.060 ;
        RECT 92.645 47.480 92.875 48.830 ;
        RECT 100.975 48.765 102.975 48.830 ;
        RECT 93.095 48.270 95.095 48.335 ;
        RECT 93.035 48.040 103.035 48.270 ;
        RECT 93.095 47.975 95.095 48.040 ;
        RECT 100.975 47.480 102.975 47.545 ;
        RECT 103.195 47.480 103.425 48.830 ;
        RECT 92.645 47.250 103.425 47.480 ;
        RECT 92.645 45.900 92.875 47.250 ;
        RECT 100.975 47.185 102.975 47.250 ;
        RECT 93.095 46.690 95.095 46.755 ;
        RECT 93.035 46.460 103.035 46.690 ;
        RECT 93.095 46.395 95.095 46.460 ;
        RECT 100.975 45.900 102.975 45.965 ;
        RECT 103.195 45.900 103.425 47.250 ;
        RECT 92.645 45.670 103.425 45.900 ;
        RECT 92.645 44.320 92.875 45.670 ;
        RECT 100.975 45.605 102.975 45.670 ;
        RECT 93.095 45.110 95.095 45.175 ;
        RECT 93.035 44.880 103.035 45.110 ;
        RECT 93.095 44.815 95.095 44.880 ;
        RECT 100.975 44.320 102.975 44.385 ;
        RECT 103.195 44.320 103.425 45.670 ;
        RECT 92.645 44.090 103.425 44.320 ;
        RECT 92.645 42.740 92.875 44.090 ;
        RECT 100.975 44.025 102.975 44.090 ;
        RECT 93.095 43.530 95.095 43.595 ;
        RECT 93.035 43.300 103.035 43.530 ;
        RECT 93.095 43.235 95.095 43.300 ;
        RECT 100.975 42.740 102.975 42.805 ;
        RECT 103.195 42.740 103.425 44.090 ;
        RECT 92.645 42.510 103.425 42.740 ;
        RECT 92.645 41.160 92.875 42.510 ;
        RECT 100.975 42.445 102.975 42.510 ;
        RECT 93.095 41.950 95.095 42.015 ;
        RECT 93.035 41.720 103.035 41.950 ;
        RECT 93.095 41.655 95.095 41.720 ;
        RECT 100.975 41.160 102.975 41.225 ;
        RECT 103.195 41.160 103.425 42.510 ;
        RECT 92.645 40.930 103.425 41.160 ;
        RECT 92.645 39.580 92.875 40.930 ;
        RECT 100.975 40.865 102.975 40.930 ;
        RECT 93.095 40.370 95.095 40.435 ;
        RECT 93.035 40.140 103.035 40.370 ;
        RECT 93.095 40.075 95.095 40.140 ;
        RECT 100.975 39.580 102.975 39.645 ;
        RECT 103.195 39.580 103.425 40.930 ;
        RECT 92.645 39.350 103.425 39.580 ;
        RECT 92.645 38.000 92.875 39.350 ;
        RECT 100.975 39.285 102.975 39.350 ;
        RECT 93.090 38.790 95.090 38.855 ;
        RECT 93.035 38.560 103.035 38.790 ;
        RECT 93.090 38.495 95.090 38.560 ;
        RECT 100.975 38.000 102.975 38.065 ;
        RECT 103.195 38.000 103.425 39.350 ;
        RECT 92.645 37.770 103.425 38.000 ;
        RECT 92.645 36.420 92.875 37.770 ;
        RECT 100.975 37.705 102.975 37.770 ;
        RECT 93.095 37.210 95.095 37.275 ;
        RECT 93.035 36.980 103.035 37.210 ;
        RECT 93.095 36.915 95.095 36.980 ;
        RECT 100.975 36.420 102.975 36.485 ;
        RECT 103.195 36.420 103.425 37.770 ;
        RECT 92.645 36.190 103.425 36.420 ;
        RECT 92.645 34.840 92.875 36.190 ;
        RECT 100.975 36.125 102.975 36.190 ;
        RECT 93.095 35.630 95.095 35.695 ;
        RECT 93.035 35.400 103.035 35.630 ;
        RECT 93.095 35.335 95.095 35.400 ;
        RECT 100.975 34.840 102.975 34.905 ;
        RECT 103.195 34.840 103.425 36.190 ;
        RECT 92.645 34.610 103.425 34.840 ;
        RECT 92.645 33.260 92.875 34.610 ;
        RECT 100.975 34.545 102.975 34.610 ;
        RECT 93.095 34.050 95.095 34.115 ;
        RECT 93.035 33.820 103.035 34.050 ;
        RECT 93.095 33.755 95.095 33.820 ;
        RECT 100.975 33.260 102.975 33.325 ;
        RECT 103.195 33.260 103.425 34.610 ;
        RECT 92.645 33.030 103.425 33.260 ;
        RECT 92.645 31.680 92.875 33.030 ;
        RECT 100.975 32.965 102.975 33.030 ;
        RECT 93.095 32.470 95.095 32.535 ;
        RECT 93.035 32.240 103.035 32.470 ;
        RECT 93.095 32.175 95.095 32.240 ;
        RECT 100.975 31.680 102.975 31.745 ;
        RECT 103.195 31.680 103.425 33.030 ;
        RECT 92.645 31.450 103.425 31.680 ;
        RECT 104.080 48.880 130.210 49.205 ;
        RECT 104.080 40.100 105.260 48.880 ;
        RECT 110.310 46.700 112.415 46.850 ;
        RECT 108.640 40.970 109.615 46.125 ;
        RECT 110.280 45.150 112.415 46.700 ;
        RECT 126.280 46.395 128.440 46.850 ;
        RECT 110.310 44.965 112.415 45.150 ;
        RECT 126.305 45.250 128.410 45.315 ;
        RECT 110.310 43.720 112.415 43.835 ;
        RECT 110.305 42.170 112.440 43.720 ;
        RECT 126.305 43.700 128.440 45.250 ;
        RECT 126.305 43.485 128.410 43.700 ;
        RECT 110.310 42.055 112.415 42.170 ;
        RECT 126.280 41.955 128.440 42.405 ;
        RECT 129.490 41.805 130.210 48.880 ;
        RECT 129.490 41.555 130.230 41.805 ;
        RECT 100.975 31.385 102.975 31.450 ;
        RECT 51.950 23.880 52.340 23.940 ;
        RECT 86.235 17.830 87.240 31.265 ;
        RECT 104.080 30.730 105.055 40.100 ;
        RECT 113.190 39.090 115.740 39.155 ;
        RECT 125.550 39.090 128.050 39.155 ;
        RECT 105.840 38.860 115.800 39.090 ;
        RECT 118.150 38.860 128.110 39.090 ;
        RECT 106.265 38.795 115.740 38.860 ;
        RECT 125.550 38.795 128.050 38.860 ;
        RECT 105.560 38.690 105.790 38.700 ;
        RECT 105.545 37.710 105.805 38.690 ;
        RECT 105.560 37.700 105.790 37.710 ;
        RECT 106.265 37.540 115.315 38.795 ;
        RECT 115.850 38.690 116.080 38.700 ;
        RECT 117.870 38.690 118.100 38.700 ;
        RECT 128.160 38.690 128.390 38.700 ;
        RECT 115.835 37.710 116.095 38.690 ;
        RECT 117.855 37.710 118.115 38.690 ;
        RECT 128.145 37.710 128.405 38.690 ;
        RECT 115.850 37.700 116.080 37.710 ;
        RECT 117.870 37.700 118.100 37.710 ;
        RECT 128.160 37.700 128.390 37.710 ;
        RECT 105.840 37.265 115.800 37.540 ;
        RECT 105.855 37.255 115.785 37.265 ;
        RECT 105.870 36.210 115.730 37.255 ;
        RECT 105.855 36.205 115.785 36.210 ;
        RECT 105.840 35.930 115.800 36.205 ;
        RECT 118.150 35.930 128.110 37.540 ;
        RECT 105.560 35.760 105.790 35.770 ;
        RECT 105.545 34.780 105.805 35.760 ;
        RECT 105.560 34.770 105.790 34.780 ;
        RECT 106.265 34.610 115.315 35.930 ;
        RECT 115.850 35.760 116.080 35.770 ;
        RECT 117.870 35.760 118.100 35.770 ;
        RECT 128.160 35.760 128.390 35.770 ;
        RECT 115.835 34.780 116.095 35.760 ;
        RECT 117.855 34.780 118.115 35.760 ;
        RECT 128.145 34.780 128.405 35.760 ;
        RECT 115.850 34.770 116.080 34.780 ;
        RECT 117.870 34.770 118.100 34.780 ;
        RECT 128.160 34.770 128.390 34.780 ;
        RECT 105.840 33.000 115.800 34.610 ;
        RECT 118.150 33.000 128.110 34.610 ;
        RECT 105.560 32.830 105.790 32.840 ;
        RECT 105.545 31.850 105.805 32.830 ;
        RECT 105.560 31.840 105.790 31.850 ;
        RECT 106.265 31.680 115.365 33.000 ;
        RECT 115.850 32.830 116.080 32.840 ;
        RECT 117.870 32.830 118.100 32.840 ;
        RECT 128.160 32.830 128.390 32.840 ;
        RECT 115.835 31.850 116.095 32.830 ;
        RECT 117.855 31.850 118.115 32.830 ;
        RECT 128.145 31.850 128.405 32.830 ;
        RECT 115.850 31.840 116.080 31.850 ;
        RECT 117.870 31.840 118.100 31.850 ;
        RECT 128.160 31.840 128.390 31.850 ;
        RECT 105.840 31.450 115.800 31.680 ;
        RECT 118.150 31.450 128.110 31.680 ;
        RECT 105.560 29.580 107.560 29.635 ;
        RECT 108.780 29.580 110.940 29.680 ;
        RECT 88.020 29.450 90.125 29.580 ;
        RECT 87.990 28.020 90.150 29.450 ;
        RECT 105.515 29.330 107.620 29.580 ;
        RECT 108.780 29.330 110.945 29.580 ;
        RECT 126.305 29.435 128.410 29.580 ;
        RECT 105.560 29.275 107.560 29.330 ;
        RECT 108.780 29.230 110.940 29.330 ;
        RECT 88.020 27.850 90.125 28.020 ;
        RECT 105.515 27.935 107.620 28.100 ;
        RECT 88.020 26.535 90.125 26.620 ;
        RECT 87.990 25.105 90.150 26.535 ;
        RECT 105.490 26.505 107.650 27.935 ;
        RECT 108.810 27.930 110.915 28.100 ;
        RECT 126.280 28.055 128.440 29.435 ;
        RECT 108.780 26.550 110.940 27.930 ;
        RECT 126.305 27.850 128.410 28.055 ;
        RECT 105.515 26.370 107.620 26.505 ;
        RECT 108.810 26.370 110.915 26.550 ;
        RECT 126.305 26.430 128.410 26.620 ;
        RECT 88.020 24.890 90.125 25.105 ;
        RECT 105.515 25.015 107.620 25.140 ;
        RECT 88.020 23.590 90.125 23.660 ;
        RECT 87.990 22.160 90.150 23.590 ;
        RECT 105.490 23.585 107.650 25.015 ;
        RECT 108.810 24.985 110.915 25.140 ;
        RECT 126.280 25.050 128.440 26.430 ;
        RECT 108.780 23.605 110.940 24.985 ;
        RECT 126.305 24.890 128.410 25.050 ;
        RECT 105.515 23.410 107.620 23.585 ;
        RECT 108.810 23.410 110.915 23.605 ;
        RECT 126.305 23.515 128.410 23.660 ;
        RECT 88.020 21.930 90.125 22.160 ;
        RECT 105.515 22.050 107.620 22.180 ;
        RECT 88.020 20.480 90.125 20.700 ;
        RECT 105.490 20.620 107.650 22.050 ;
        RECT 108.810 21.975 110.915 22.180 ;
        RECT 126.280 22.135 128.440 23.515 ;
        RECT 87.990 19.200 90.150 20.480 ;
        RECT 105.515 20.450 107.620 20.620 ;
        RECT 108.780 20.595 110.940 21.975 ;
        RECT 126.305 21.930 128.410 22.135 ;
        RECT 108.810 20.450 110.915 20.595 ;
        RECT 126.305 20.520 128.410 20.700 ;
        RECT 107.485 19.220 108.980 19.270 ;
        RECT 88.020 18.970 90.125 19.200 ;
        RECT 105.515 18.970 110.915 19.220 ;
        RECT 126.280 19.140 128.440 20.520 ;
        RECT 126.305 18.970 128.410 19.140 ;
        RECT 107.485 18.920 108.980 18.970 ;
        RECT 129.490 17.830 130.210 41.555 ;
        RECT 145.445 28.805 146.585 50.190 ;
        RECT 152.260 49.840 157.360 49.855 ;
        RECT 147.370 49.610 157.370 49.840 ;
        RECT 152.260 49.595 157.360 49.610 ;
        RECT 146.980 48.465 147.210 49.560 ;
        RECT 157.530 48.465 157.760 49.560 ;
        RECT 146.980 42.260 157.760 48.465 ;
        RECT 146.980 40.680 147.210 42.260 ;
        RECT 157.530 40.720 157.760 42.260 ;
        RECT 146.980 38.310 147.215 40.680 ;
        RECT 147.380 40.550 152.480 40.565 ;
        RECT 147.370 40.320 157.370 40.550 ;
        RECT 147.380 40.305 152.480 40.320 ;
        RECT 147.380 38.640 152.480 38.655 ;
        RECT 147.370 38.410 157.370 38.640 ;
        RECT 147.380 38.395 152.480 38.410 ;
        RECT 157.530 38.320 157.765 40.720 ;
        RECT 146.980 37.110 147.210 38.310 ;
        RECT 157.530 37.110 157.760 38.320 ;
        RECT 146.980 32.460 157.760 37.110 ;
        RECT 146.915 30.905 157.760 32.460 ;
        RECT 158.255 30.965 159.285 50.190 ;
        RECT 161.285 44.935 162.005 50.545 ;
        RECT 162.400 49.905 163.640 50.135 ;
        RECT 162.400 49.640 162.630 49.905 ;
        RECT 163.690 49.640 163.920 49.700 ;
        RECT 162.340 45.760 162.700 49.640 ;
        RECT 163.620 47.640 164.025 49.640 ;
        RECT 162.400 45.495 162.630 45.760 ;
        RECT 163.690 45.700 163.920 47.640 ;
        RECT 162.400 45.265 163.640 45.495 ;
        RECT 164.360 44.935 166.255 50.545 ;
        RECT 166.770 49.025 167.000 54.965 ;
        RECT 166.705 45.025 167.065 49.025 ;
        RECT 166.770 44.965 167.000 45.025 ;
        RECT 161.285 44.215 166.255 44.935 ;
        RECT 167.265 44.760 167.730 55.170 ;
        RECT 168.060 54.905 168.290 54.965 ;
        RECT 167.990 50.905 168.350 54.905 ;
        RECT 168.060 44.965 168.290 50.905 ;
        RECT 168.570 44.760 169.035 55.170 ;
        RECT 169.350 49.025 169.580 54.965 ;
        RECT 169.285 45.025 169.645 49.025 ;
        RECT 169.350 44.965 169.580 45.025 ;
        RECT 169.905 44.760 170.370 55.170 ;
        RECT 170.640 54.910 170.870 54.965 ;
        RECT 170.575 50.910 170.935 54.910 ;
        RECT 170.640 44.965 170.870 50.910 ;
        RECT 171.210 44.760 171.675 55.170 ;
        RECT 171.930 49.025 172.160 54.965 ;
        RECT 171.865 45.025 172.225 49.025 ;
        RECT 171.930 44.965 172.160 45.025 ;
        RECT 172.480 44.760 172.945 55.170 ;
        RECT 173.220 54.910 173.450 54.965 ;
        RECT 173.155 50.910 173.515 54.910 ;
        RECT 173.220 44.965 173.450 50.910 ;
        RECT 173.725 44.760 174.190 55.170 ;
        RECT 174.510 49.025 174.740 54.965 ;
        RECT 174.445 45.025 174.805 49.025 ;
        RECT 174.510 44.965 174.740 45.025 ;
        RECT 175.030 44.760 175.495 55.170 ;
        RECT 175.800 54.905 176.030 54.965 ;
        RECT 175.735 50.905 176.095 54.905 ;
        RECT 175.800 44.965 176.030 50.905 ;
        RECT 176.335 44.760 176.800 55.170 ;
        RECT 177.090 49.025 177.320 54.965 ;
        RECT 177.025 45.025 177.385 49.025 ;
        RECT 177.090 44.965 177.320 45.025 ;
        RECT 177.605 44.760 178.070 55.170 ;
        RECT 178.380 54.910 178.610 54.965 ;
        RECT 178.315 50.910 178.675 54.910 ;
        RECT 178.380 44.965 178.610 50.910 ;
        RECT 178.880 44.760 179.345 55.170 ;
        RECT 179.670 49.025 179.900 54.965 ;
        RECT 179.605 45.025 179.965 49.025 ;
        RECT 179.670 44.965 179.900 45.025 ;
        RECT 167.050 44.530 179.620 44.760 ;
        RECT 161.285 44.185 162.005 44.215 ;
        RECT 165.380 44.115 166.255 44.215 ;
        RECT 180.270 44.115 181.475 55.890 ;
        RECT 182.125 55.400 182.660 55.445 ;
        RECT 182.115 55.170 188.235 55.400 ;
        RECT 181.835 49.025 182.065 54.965 ;
        RECT 181.770 45.025 182.130 49.025 ;
        RECT 181.835 44.965 182.065 45.025 ;
        RECT 182.390 44.760 182.855 55.170 ;
        RECT 183.125 54.905 183.355 54.965 ;
        RECT 183.055 50.905 183.415 54.905 ;
        RECT 183.125 44.965 183.355 50.905 ;
        RECT 183.665 44.760 184.130 55.170 ;
        RECT 184.415 49.025 184.645 54.965 ;
        RECT 184.350 45.025 184.710 49.025 ;
        RECT 184.415 44.965 184.645 45.025 ;
        RECT 184.935 44.760 185.400 55.170 ;
        RECT 185.705 54.910 185.935 54.965 ;
        RECT 185.640 50.910 186.000 54.910 ;
        RECT 185.705 44.965 185.935 50.910 ;
        RECT 186.240 44.760 186.705 55.170 ;
        RECT 186.995 49.025 187.225 54.965 ;
        RECT 186.930 45.025 187.290 49.025 ;
        RECT 186.995 44.965 187.225 45.025 ;
        RECT 187.485 44.760 187.950 55.170 ;
        RECT 188.285 54.900 188.515 54.965 ;
        RECT 188.220 50.900 188.580 54.900 ;
        RECT 188.945 52.445 194.570 55.890 ;
        RECT 188.285 44.965 188.515 50.900 ;
        RECT 188.945 50.825 194.575 52.445 ;
        RECT 188.945 50.760 194.580 50.825 ;
        RECT 182.115 44.530 188.235 44.760 ;
        RECT 188.945 44.115 190.070 50.760 ;
        RECT 192.950 50.725 194.580 50.760 ;
        RECT 190.735 50.305 191.265 50.365 ;
        RECT 190.725 50.075 192.975 50.305 ;
        RECT 190.445 48.930 190.675 49.870 ;
        RECT 190.380 44.930 190.740 48.930 ;
        RECT 190.445 44.870 190.675 44.930 ;
        RECT 190.965 44.665 191.365 50.075 ;
        RECT 191.735 49.810 191.965 49.870 ;
        RECT 191.670 47.095 192.030 49.810 ;
        RECT 191.735 44.870 191.965 47.095 ;
        RECT 192.265 44.665 192.665 50.075 ;
        RECT 193.025 48.930 193.255 49.870 ;
        RECT 192.960 44.930 193.320 48.930 ;
        RECT 193.025 44.870 193.255 44.930 ;
        RECT 190.725 44.435 192.975 44.665 ;
        RECT 165.380 44.085 190.070 44.115 ;
        RECT 165.380 43.505 190.220 44.085 ;
        RECT 165.335 42.875 190.220 43.505 ;
        RECT 165.335 32.875 166.365 42.875 ;
        RECT 170.085 42.825 174.390 42.875 ;
        RECT 170.225 42.810 174.390 42.825 ;
        RECT 166.995 42.515 168.585 42.565 ;
        RECT 166.995 42.285 177.035 42.515 ;
        RECT 166.765 37.640 166.995 42.080 ;
        RECT 166.700 33.640 167.060 37.640 ;
        RECT 166.765 33.580 166.995 33.640 ;
        RECT 167.275 33.375 167.725 42.285 ;
        RECT 168.055 42.020 168.285 42.080 ;
        RECT 167.990 38.020 168.350 42.020 ;
        RECT 168.055 33.580 168.285 38.020 ;
        RECT 168.610 33.375 169.060 42.285 ;
        RECT 169.345 37.640 169.575 42.080 ;
        RECT 169.280 33.640 169.640 37.640 ;
        RECT 169.345 33.580 169.575 33.640 ;
        RECT 169.895 33.375 170.345 42.285 ;
        RECT 170.635 42.020 170.865 42.080 ;
        RECT 170.570 38.020 170.930 42.020 ;
        RECT 170.635 33.580 170.865 38.020 ;
        RECT 171.185 33.375 171.635 42.285 ;
        RECT 171.925 37.640 172.155 42.080 ;
        RECT 171.860 33.640 172.220 37.640 ;
        RECT 171.925 33.580 172.155 33.640 ;
        RECT 172.500 33.375 172.950 42.285 ;
        RECT 173.215 42.045 173.445 42.080 ;
        RECT 173.150 38.045 173.510 42.045 ;
        RECT 173.215 33.580 173.445 38.045 ;
        RECT 173.725 33.375 174.175 42.285 ;
        RECT 174.505 37.640 174.735 42.080 ;
        RECT 174.440 33.640 174.800 37.640 ;
        RECT 174.505 33.580 174.735 33.640 ;
        RECT 175.045 33.375 175.495 42.285 ;
        RECT 175.795 42.025 176.025 42.080 ;
        RECT 175.730 38.025 176.090 42.025 ;
        RECT 175.795 33.580 176.025 38.025 ;
        RECT 176.330 33.375 176.780 42.285 ;
        RECT 177.085 37.640 177.315 42.080 ;
        RECT 177.740 40.785 190.220 42.875 ;
        RECT 177.020 33.640 177.380 37.640 ;
        RECT 177.740 34.940 181.810 40.785 ;
        RECT 182.505 40.290 183.210 40.350 ;
        RECT 182.495 40.060 184.745 40.290 ;
        RECT 182.215 36.845 182.445 39.855 ;
        RECT 182.150 35.915 182.510 36.845 ;
        RECT 182.215 35.855 182.445 35.915 ;
        RECT 182.700 35.650 183.165 40.060 ;
        RECT 183.320 40.055 183.930 40.060 ;
        RECT 183.505 39.795 183.735 39.855 ;
        RECT 183.440 38.865 183.800 39.795 ;
        RECT 183.505 35.855 183.735 38.865 ;
        RECT 184.100 35.650 184.565 40.060 ;
        RECT 185.495 39.925 190.220 40.785 ;
        RECT 193.700 41.050 194.580 50.725 ;
        RECT 194.950 45.685 195.180 66.625 ;
        RECT 194.885 41.685 195.245 45.685 ;
        RECT 194.950 41.625 195.180 41.685 ;
        RECT 195.490 41.420 195.880 66.830 ;
        RECT 196.240 66.610 196.470 66.625 ;
        RECT 196.140 62.610 196.500 66.610 ;
        RECT 196.240 41.625 196.470 62.610 ;
        RECT 196.800 41.420 197.190 66.830 ;
        RECT 197.530 45.680 197.760 66.625 ;
        RECT 197.465 41.680 197.825 45.680 ;
        RECT 197.530 41.625 197.760 41.680 ;
        RECT 198.105 41.420 198.495 66.830 ;
        RECT 198.820 66.610 199.050 66.625 ;
        RECT 198.755 62.610 199.115 66.610 ;
        RECT 198.820 41.625 199.050 62.610 ;
        RECT 199.410 41.420 199.800 66.830 ;
        RECT 200.110 45.690 200.340 66.625 ;
        RECT 200.050 41.690 200.410 45.690 ;
        RECT 200.110 41.625 200.340 41.690 ;
        RECT 200.690 41.420 201.080 66.830 ;
        RECT 201.400 66.570 201.630 66.625 ;
        RECT 201.325 62.570 201.685 66.570 ;
        RECT 201.400 41.625 201.630 62.570 ;
        RECT 201.995 41.420 202.385 66.830 ;
        RECT 202.690 45.675 202.920 66.625 ;
        RECT 202.640 41.675 203.000 45.675 ;
        RECT 202.690 41.625 202.920 41.675 ;
        RECT 203.255 41.420 203.645 66.830 ;
        RECT 203.980 66.570 204.210 66.625 ;
        RECT 203.930 62.570 204.290 66.570 ;
        RECT 203.980 41.625 204.210 62.570 ;
        RECT 204.500 41.420 204.890 66.830 ;
        RECT 205.270 45.675 205.500 66.625 ;
        RECT 205.200 41.675 205.560 45.675 ;
        RECT 205.270 41.625 205.500 41.675 ;
        RECT 205.805 41.420 206.195 66.830 ;
        RECT 206.560 66.550 206.790 66.625 ;
        RECT 206.510 62.550 206.870 66.550 ;
        RECT 206.560 41.625 206.790 62.550 ;
        RECT 207.065 41.435 207.455 66.830 ;
        RECT 207.850 45.680 208.080 66.625 ;
        RECT 208.575 65.510 209.300 67.515 ;
        RECT 210.080 67.060 210.645 67.115 ;
        RECT 210.070 66.830 222.640 67.060 ;
        RECT 207.775 41.680 208.135 45.680 ;
        RECT 208.475 42.795 209.395 65.510 ;
        RECT 209.790 45.670 210.020 66.625 ;
        RECT 207.850 41.625 208.080 41.680 ;
        RECT 207.065 41.420 207.790 41.435 ;
        RECT 195.230 41.190 207.800 41.420 ;
        RECT 207.350 41.175 207.790 41.190 ;
        RECT 193.700 40.790 195.655 41.050 ;
        RECT 193.700 40.785 195.685 40.790 ;
        RECT 197.055 40.785 198.240 40.790 ;
        RECT 202.290 40.785 203.475 40.790 ;
        RECT 208.575 40.785 209.300 42.795 ;
        RECT 209.700 41.670 210.060 45.670 ;
        RECT 209.790 41.625 210.020 41.670 ;
        RECT 210.380 41.430 210.770 66.830 ;
        RECT 211.080 66.560 211.310 66.625 ;
        RECT 211.020 62.560 211.380 66.560 ;
        RECT 211.080 41.625 211.310 62.560 ;
        RECT 210.080 41.420 210.770 41.430 ;
        RECT 211.655 41.420 212.045 66.830 ;
        RECT 212.370 45.670 212.600 66.625 ;
        RECT 212.295 41.670 212.655 45.670 ;
        RECT 212.370 41.625 212.600 41.670 ;
        RECT 212.930 41.420 213.320 66.830 ;
        RECT 213.660 66.560 213.890 66.625 ;
        RECT 213.595 62.560 213.955 66.560 ;
        RECT 213.660 41.625 213.890 62.560 ;
        RECT 214.190 41.420 214.580 66.830 ;
        RECT 214.950 45.670 215.180 66.625 ;
        RECT 214.885 41.670 215.245 45.670 ;
        RECT 214.950 41.625 215.180 41.670 ;
        RECT 215.470 41.420 215.860 66.830 ;
        RECT 216.240 66.580 216.470 66.625 ;
        RECT 216.190 62.580 216.550 66.580 ;
        RECT 216.240 41.625 216.470 62.580 ;
        RECT 216.790 41.420 217.180 66.830 ;
        RECT 217.530 45.695 217.760 66.625 ;
        RECT 217.435 41.695 217.795 45.695 ;
        RECT 217.530 41.625 217.760 41.695 ;
        RECT 218.095 41.420 218.485 66.830 ;
        RECT 218.820 66.560 219.050 66.625 ;
        RECT 218.745 62.560 219.105 66.560 ;
        RECT 218.820 41.625 219.050 62.560 ;
        RECT 219.340 41.420 219.730 66.830 ;
        RECT 220.110 45.670 220.340 66.625 ;
        RECT 220.050 41.670 220.410 45.670 ;
        RECT 220.110 41.625 220.340 41.670 ;
        RECT 220.680 41.420 221.070 66.830 ;
        RECT 221.400 66.560 221.630 66.625 ;
        RECT 221.320 62.560 221.680 66.560 ;
        RECT 221.400 41.625 221.630 62.560 ;
        RECT 221.955 41.420 222.345 66.830 ;
        RECT 222.690 45.670 222.920 66.625 ;
        RECT 222.620 41.670 222.980 45.670 ;
        RECT 222.690 41.625 222.920 41.670 ;
        RECT 210.070 41.190 222.640 41.420 ;
        RECT 210.080 41.170 210.520 41.190 ;
        RECT 223.265 40.785 224.560 67.515 ;
        RECT 193.700 39.925 224.560 40.785 ;
        RECT 184.795 36.845 185.025 39.855 ;
        RECT 185.495 39.675 224.560 39.925 ;
        RECT 185.495 38.850 194.580 39.675 ;
        RECT 195.205 39.305 195.975 39.365 ;
        RECT 197.260 39.305 198.030 39.410 ;
        RECT 199.855 39.305 200.625 39.380 ;
        RECT 202.465 39.305 203.235 39.395 ;
        RECT 205.045 39.305 205.815 39.380 ;
        RECT 195.205 39.075 207.800 39.305 ;
        RECT 195.205 39.065 195.975 39.075 ;
        RECT 184.730 35.915 185.090 36.845 ;
        RECT 185.495 36.080 190.220 38.850 ;
        RECT 190.880 38.415 191.935 38.530 ;
        RECT 190.880 38.185 192.960 38.415 ;
        RECT 190.720 37.685 190.950 37.980 ;
        RECT 190.650 37.040 191.020 37.685 ;
        RECT 190.720 36.980 190.950 37.040 ;
        RECT 191.365 36.775 192.330 38.185 ;
        RECT 193.010 37.525 193.240 37.980 ;
        RECT 192.945 37.040 193.305 37.525 ;
        RECT 193.010 36.980 193.240 37.040 ;
        RECT 191.000 36.545 192.960 36.775 ;
        RECT 193.700 36.080 194.580 38.850 ;
        RECT 184.795 35.855 185.025 35.915 ;
        RECT 182.495 35.420 183.455 35.650 ;
        RECT 183.785 35.420 184.745 35.650 ;
        RECT 185.495 34.940 194.580 36.080 ;
        RECT 177.740 34.195 194.580 34.940 ;
        RECT 177.085 33.580 177.315 33.640 ;
        RECT 167.045 33.145 168.005 33.375 ;
        RECT 168.335 33.145 169.295 33.375 ;
        RECT 169.625 33.145 170.585 33.375 ;
        RECT 170.915 33.145 171.875 33.375 ;
        RECT 172.205 33.145 173.165 33.375 ;
        RECT 173.495 33.145 174.455 33.375 ;
        RECT 174.785 33.145 175.745 33.375 ;
        RECT 176.075 33.145 177.035 33.375 ;
        RECT 177.740 32.875 179.120 34.195 ;
        RECT 165.335 31.975 179.120 32.875 ;
        RECT 165.660 31.925 179.120 31.975 ;
        RECT 177.740 31.895 179.120 31.925 ;
        RECT 161.195 30.975 174.540 30.985 ;
        RECT 160.255 30.965 174.540 30.975 ;
        RECT 146.915 29.460 147.275 30.905 ;
        RECT 146.980 29.400 147.210 29.460 ;
        RECT 157.530 29.400 157.760 30.905 ;
        RECT 158.225 29.740 174.540 30.965 ;
        RECT 158.225 29.685 174.525 29.740 ;
        RECT 152.260 29.350 157.360 29.365 ;
        RECT 147.370 29.120 157.370 29.350 ;
        RECT 152.260 29.105 157.360 29.120 ;
        RECT 158.225 28.805 161.945 29.685 ;
        RECT 162.800 29.350 167.900 29.365 ;
        RECT 162.790 29.120 172.790 29.350 ;
        RECT 162.800 29.105 167.900 29.120 ;
        RECT 145.420 28.705 161.945 28.805 ;
        RECT 145.420 28.410 161.885 28.705 ;
        RECT 162.400 28.635 162.630 29.070 ;
        RECT 145.420 25.990 161.905 28.410 ;
        RECT 145.455 19.270 146.230 25.990 ;
        RECT 146.930 25.205 147.490 25.245 ;
        RECT 146.920 24.975 159.490 25.205 ;
        RECT 146.640 21.875 146.870 24.815 ;
        RECT 146.575 19.875 146.935 21.875 ;
        RECT 146.640 19.815 146.870 19.875 ;
        RECT 147.090 19.655 147.595 24.975 ;
        RECT 147.930 24.755 148.160 24.815 ;
        RECT 147.865 22.755 148.225 24.755 ;
        RECT 147.930 19.815 148.160 22.755 ;
        RECT 148.400 19.655 148.905 24.975 ;
        RECT 149.220 21.875 149.450 24.815 ;
        RECT 149.155 19.875 149.515 21.875 ;
        RECT 149.220 19.815 149.450 19.875 ;
        RECT 149.745 19.655 150.250 24.975 ;
        RECT 150.510 24.755 150.740 24.815 ;
        RECT 150.445 22.755 150.805 24.755 ;
        RECT 150.510 19.815 150.740 22.755 ;
        RECT 151.025 19.655 151.530 24.975 ;
        RECT 151.800 21.875 152.030 24.815 ;
        RECT 151.735 19.875 152.095 21.875 ;
        RECT 151.800 19.815 152.030 19.875 ;
        RECT 152.325 19.655 152.830 24.975 ;
        RECT 153.090 24.760 153.320 24.815 ;
        RECT 153.025 22.760 153.385 24.760 ;
        RECT 153.090 19.815 153.320 22.760 ;
        RECT 153.620 19.655 154.125 24.975 ;
        RECT 154.380 21.875 154.610 24.815 ;
        RECT 154.315 19.875 154.675 21.875 ;
        RECT 154.380 19.815 154.610 19.875 ;
        RECT 154.900 19.655 155.405 24.975 ;
        RECT 155.670 24.755 155.900 24.815 ;
        RECT 155.605 22.755 155.965 24.755 ;
        RECT 155.670 19.815 155.900 22.755 ;
        RECT 156.145 19.655 156.650 24.975 ;
        RECT 156.960 21.875 157.190 24.815 ;
        RECT 156.895 19.875 157.255 21.875 ;
        RECT 156.960 19.815 157.190 19.875 ;
        RECT 157.475 19.655 157.980 24.975 ;
        RECT 158.250 24.755 158.480 24.815 ;
        RECT 158.185 22.755 158.545 24.755 ;
        RECT 158.250 19.815 158.480 22.755 ;
        RECT 158.740 19.655 159.245 24.975 ;
        RECT 159.540 21.870 159.770 24.815 ;
        RECT 159.475 19.870 159.835 21.870 ;
        RECT 160.215 20.895 161.905 25.990 ;
        RECT 162.325 27.280 162.705 28.635 ;
        RECT 172.950 27.280 173.180 29.070 ;
        RECT 162.325 24.635 173.180 27.280 ;
        RECT 162.400 21.075 173.180 24.635 ;
        RECT 159.540 19.815 159.770 19.870 ;
        RECT 146.920 19.425 159.490 19.655 ;
        RECT 160.255 19.270 161.885 20.895 ;
        RECT 162.400 20.110 162.630 21.075 ;
        RECT 172.950 20.110 173.180 21.075 ;
        RECT 162.800 20.060 167.900 20.075 ;
        RECT 162.790 19.830 172.790 20.060 ;
        RECT 162.800 19.815 167.900 19.830 ;
        RECT 173.565 19.270 174.515 29.685 ;
        RECT 193.700 20.075 194.580 34.195 ;
        RECT 194.950 24.925 195.180 38.870 ;
        RECT 194.895 20.925 195.255 24.925 ;
        RECT 194.950 20.870 195.180 20.925 ;
        RECT 195.475 20.665 195.865 39.065 ;
        RECT 196.240 38.825 196.470 38.870 ;
        RECT 196.185 34.825 196.545 38.825 ;
        RECT 196.240 20.870 196.470 34.825 ;
        RECT 196.785 20.665 197.175 39.075 ;
        RECT 197.530 24.930 197.760 38.870 ;
        RECT 197.440 20.930 197.800 24.930 ;
        RECT 197.530 20.870 197.760 20.930 ;
        RECT 198.045 20.665 198.435 39.075 ;
        RECT 198.820 38.850 199.050 38.870 ;
        RECT 198.715 34.850 199.075 38.850 ;
        RECT 198.820 20.870 199.050 34.850 ;
        RECT 199.335 20.665 199.725 39.075 ;
        RECT 200.110 24.920 200.340 38.870 ;
        RECT 200.040 20.920 200.400 24.920 ;
        RECT 200.110 20.870 200.340 20.920 ;
        RECT 200.625 20.665 201.015 39.075 ;
        RECT 201.400 38.850 201.630 38.870 ;
        RECT 201.335 34.850 201.695 38.850 ;
        RECT 201.400 20.870 201.630 34.850 ;
        RECT 201.950 20.665 202.340 39.075 ;
        RECT 202.690 24.920 202.920 38.870 ;
        RECT 202.630 20.920 202.990 24.920 ;
        RECT 202.690 20.870 202.920 20.920 ;
        RECT 203.225 20.665 203.615 39.075 ;
        RECT 203.980 38.825 204.210 38.870 ;
        RECT 203.930 34.825 204.290 38.825 ;
        RECT 203.980 20.870 204.210 34.825 ;
        RECT 204.485 20.665 204.875 39.075 ;
        RECT 205.270 24.920 205.500 38.870 ;
        RECT 205.190 20.920 205.550 24.920 ;
        RECT 205.270 20.870 205.500 20.920 ;
        RECT 205.855 20.665 206.245 39.075 ;
        RECT 206.560 38.825 206.790 38.870 ;
        RECT 206.505 34.825 206.865 38.825 ;
        RECT 206.560 20.870 206.790 34.825 ;
        RECT 207.100 20.665 207.490 39.075 ;
        RECT 207.850 24.920 208.080 38.870 ;
        RECT 208.535 38.040 209.670 39.675 ;
        RECT 210.245 39.230 211.015 39.305 ;
        RECT 212.435 39.230 213.205 39.335 ;
        RECT 214.910 39.230 215.680 39.335 ;
        RECT 217.610 39.230 218.380 39.335 ;
        RECT 220.145 39.230 220.915 39.350 ;
        RECT 210.245 39.005 222.915 39.230 ;
        RECT 210.345 39.000 222.915 39.005 ;
        RECT 207.770 20.920 208.130 24.920 ;
        RECT 208.525 21.895 209.685 38.040 ;
        RECT 210.065 24.865 210.295 38.795 ;
        RECT 207.850 20.870 208.080 20.920 ;
        RECT 195.230 20.435 207.800 20.665 ;
        RECT 195.965 20.430 207.785 20.435 ;
        RECT 208.535 20.075 209.670 21.895 ;
        RECT 210.015 20.865 210.375 24.865 ;
        RECT 210.065 20.795 210.295 20.865 ;
        RECT 210.615 20.595 211.005 39.000 ;
        RECT 211.355 38.760 211.585 38.795 ;
        RECT 211.300 34.760 211.660 38.760 ;
        RECT 211.355 20.795 211.585 34.760 ;
        RECT 211.875 20.595 212.265 39.000 ;
        RECT 212.645 24.855 212.875 38.795 ;
        RECT 212.585 20.855 212.945 24.855 ;
        RECT 212.645 20.795 212.875 20.855 ;
        RECT 213.210 20.595 213.600 39.000 ;
        RECT 213.935 38.785 214.165 38.795 ;
        RECT 213.880 34.785 214.240 38.785 ;
        RECT 213.935 20.795 214.165 34.785 ;
        RECT 214.520 20.595 214.910 39.000 ;
        RECT 215.225 24.855 215.455 38.795 ;
        RECT 215.185 20.855 215.545 24.855 ;
        RECT 215.225 20.795 215.455 20.855 ;
        RECT 215.795 20.595 216.185 39.000 ;
        RECT 216.515 38.760 216.745 38.795 ;
        RECT 216.430 34.760 216.790 38.760 ;
        RECT 216.515 20.795 216.745 34.760 ;
        RECT 217.100 20.595 217.490 39.000 ;
        RECT 217.805 24.845 218.035 38.795 ;
        RECT 217.745 20.845 218.105 24.845 ;
        RECT 217.805 20.795 218.035 20.845 ;
        RECT 218.375 20.595 218.765 39.000 ;
        RECT 219.095 38.760 219.325 38.795 ;
        RECT 219.030 34.760 219.390 38.760 ;
        RECT 219.095 20.795 219.325 34.760 ;
        RECT 219.670 20.595 220.060 39.000 ;
        RECT 220.385 24.845 220.615 38.795 ;
        RECT 220.325 20.845 220.685 24.845 ;
        RECT 220.385 20.795 220.615 20.845 ;
        RECT 220.960 20.595 221.350 39.000 ;
        RECT 221.675 38.740 221.905 38.795 ;
        RECT 221.625 34.740 221.985 38.740 ;
        RECT 221.675 20.795 221.905 34.740 ;
        RECT 222.220 20.595 222.610 39.000 ;
        RECT 222.965 24.855 223.195 38.795 ;
        RECT 222.905 20.855 223.265 24.855 ;
        RECT 222.965 20.795 223.195 20.855 ;
        RECT 210.430 20.590 222.610 20.595 ;
        RECT 210.345 20.360 222.915 20.590 ;
        RECT 223.580 20.075 224.560 39.675 ;
        RECT 229.655 65.360 230.430 67.940 ;
        RECT 232.915 67.395 233.315 67.460 ;
        RECT 231.375 67.165 233.375 67.395 ;
        RECT 230.940 66.155 231.170 67.115 ;
        RECT 232.915 67.100 233.315 67.165 ;
        RECT 233.580 66.665 233.810 67.115 ;
        RECT 231.435 66.105 231.835 66.170 ;
        RECT 233.565 66.165 233.825 66.665 ;
        RECT 233.580 66.155 233.810 66.165 ;
        RECT 231.375 65.875 233.375 66.105 ;
        RECT 231.435 65.810 231.835 65.875 ;
        RECT 234.205 65.360 234.855 67.940 ;
        RECT 229.655 64.715 234.855 65.360 ;
        RECT 229.655 62.175 230.430 64.715 ;
        RECT 231.435 64.200 231.835 64.265 ;
        RECT 231.375 63.970 233.375 64.200 ;
        RECT 230.940 62.960 231.170 63.920 ;
        RECT 231.435 63.905 231.835 63.970 ;
        RECT 233.580 63.910 233.810 63.920 ;
        RECT 233.565 63.410 233.825 63.910 ;
        RECT 232.915 62.910 233.315 62.975 ;
        RECT 233.580 62.960 233.810 63.410 ;
        RECT 231.375 62.680 233.375 62.910 ;
        RECT 232.915 62.615 233.315 62.680 ;
        RECT 234.205 62.175 234.855 64.715 ;
        RECT 229.655 61.530 234.855 62.175 ;
        RECT 229.655 58.950 230.430 61.530 ;
        RECT 231.430 61.005 231.830 61.070 ;
        RECT 231.370 60.775 233.370 61.005 ;
        RECT 230.935 59.765 231.165 60.725 ;
        RECT 231.430 60.710 231.830 60.775 ;
        RECT 233.575 60.715 233.805 60.725 ;
        RECT 233.560 60.215 233.820 60.715 ;
        RECT 232.910 59.715 233.310 59.780 ;
        RECT 233.575 59.765 233.805 60.215 ;
        RECT 231.370 59.485 233.370 59.715 ;
        RECT 232.910 59.420 233.310 59.485 ;
        RECT 234.205 58.950 234.855 61.530 ;
        RECT 229.655 58.305 234.855 58.950 ;
        RECT 229.655 55.790 230.430 58.305 ;
        RECT 231.430 57.810 231.830 57.875 ;
        RECT 231.370 57.580 233.370 57.810 ;
        RECT 230.935 56.570 231.165 57.530 ;
        RECT 231.430 57.515 231.830 57.580 ;
        RECT 233.575 57.520 233.805 57.530 ;
        RECT 233.560 57.020 233.820 57.520 ;
        RECT 232.910 56.520 233.310 56.585 ;
        RECT 233.575 56.570 233.805 57.020 ;
        RECT 231.370 56.290 233.370 56.520 ;
        RECT 232.910 56.225 233.310 56.290 ;
        RECT 234.205 55.790 234.855 58.305 ;
        RECT 229.655 55.145 234.855 55.790 ;
        RECT 229.655 52.585 230.430 55.145 ;
        RECT 231.430 54.615 231.830 54.680 ;
        RECT 231.370 54.385 233.370 54.615 ;
        RECT 230.935 53.375 231.165 54.335 ;
        RECT 231.430 54.320 231.830 54.385 ;
        RECT 233.575 54.325 233.805 54.335 ;
        RECT 233.560 53.825 233.820 54.325 ;
        RECT 232.910 53.325 233.310 53.390 ;
        RECT 233.575 53.375 233.805 53.825 ;
        RECT 231.370 53.095 233.370 53.325 ;
        RECT 232.910 53.030 233.310 53.095 ;
        RECT 234.205 52.585 234.855 55.145 ;
        RECT 229.655 51.940 234.855 52.585 ;
        RECT 229.655 49.405 230.430 51.940 ;
        RECT 231.430 51.420 231.830 51.485 ;
        RECT 231.370 51.190 233.370 51.420 ;
        RECT 230.935 50.180 231.165 51.140 ;
        RECT 231.430 51.125 231.830 51.190 ;
        RECT 233.575 51.130 233.805 51.140 ;
        RECT 233.560 50.630 233.820 51.130 ;
        RECT 232.910 50.130 233.310 50.195 ;
        RECT 233.575 50.180 233.805 50.630 ;
        RECT 231.370 49.900 233.370 50.130 ;
        RECT 232.910 49.835 233.310 49.900 ;
        RECT 234.205 49.405 234.855 51.940 ;
        RECT 229.655 48.760 234.855 49.405 ;
        RECT 229.655 46.155 230.430 48.760 ;
        RECT 231.430 48.225 231.830 48.290 ;
        RECT 231.370 47.995 233.370 48.225 ;
        RECT 230.935 46.985 231.165 47.945 ;
        RECT 231.430 47.930 231.830 47.995 ;
        RECT 233.575 47.935 233.805 47.945 ;
        RECT 233.560 47.435 233.820 47.935 ;
        RECT 232.910 46.935 233.310 47.000 ;
        RECT 233.575 46.985 233.805 47.435 ;
        RECT 231.370 46.705 233.370 46.935 ;
        RECT 232.910 46.640 233.310 46.705 ;
        RECT 234.205 46.155 234.855 48.760 ;
        RECT 229.655 45.510 234.855 46.155 ;
        RECT 229.655 43.040 230.430 45.510 ;
        RECT 231.430 45.030 231.830 45.095 ;
        RECT 231.370 44.800 233.370 45.030 ;
        RECT 234.205 44.870 234.855 45.510 ;
        RECT 230.935 43.790 231.165 44.750 ;
        RECT 231.430 44.735 231.830 44.800 ;
        RECT 233.575 44.740 233.805 44.750 ;
        RECT 233.560 44.240 233.820 44.740 ;
        RECT 234.200 44.285 234.855 44.870 ;
        RECT 232.910 43.740 233.310 43.805 ;
        RECT 233.575 43.790 233.805 44.240 ;
        RECT 231.370 43.510 233.370 43.740 ;
        RECT 232.910 43.445 233.310 43.510 ;
        RECT 234.205 43.040 234.855 44.285 ;
        RECT 229.655 42.395 234.855 43.040 ;
        RECT 229.655 39.815 230.430 42.395 ;
        RECT 231.430 41.835 231.830 41.900 ;
        RECT 231.370 41.605 233.370 41.835 ;
        RECT 230.935 40.595 231.165 41.555 ;
        RECT 231.430 41.540 231.830 41.605 ;
        RECT 233.575 41.545 233.805 41.555 ;
        RECT 233.560 41.045 233.820 41.545 ;
        RECT 232.910 40.545 233.310 40.610 ;
        RECT 233.575 40.595 233.805 41.045 ;
        RECT 231.370 40.315 233.370 40.545 ;
        RECT 232.910 40.250 233.310 40.315 ;
        RECT 234.205 39.815 234.855 42.395 ;
        RECT 229.655 39.170 234.855 39.815 ;
        RECT 229.655 36.610 230.430 39.170 ;
        RECT 231.430 38.640 231.830 38.705 ;
        RECT 231.370 38.410 233.370 38.640 ;
        RECT 230.935 37.400 231.165 38.360 ;
        RECT 231.430 38.345 231.830 38.410 ;
        RECT 233.575 38.350 233.805 38.360 ;
        RECT 233.560 37.850 233.820 38.350 ;
        RECT 232.910 37.350 233.310 37.415 ;
        RECT 233.575 37.400 233.805 37.850 ;
        RECT 231.370 37.120 233.370 37.350 ;
        RECT 232.910 37.055 233.310 37.120 ;
        RECT 234.205 36.610 234.855 39.170 ;
        RECT 229.655 35.965 234.855 36.610 ;
        RECT 229.655 33.405 230.430 35.965 ;
        RECT 231.430 35.445 231.830 35.510 ;
        RECT 231.370 35.215 233.370 35.445 ;
        RECT 230.935 34.205 231.165 35.165 ;
        RECT 231.430 35.150 231.830 35.215 ;
        RECT 233.575 35.155 233.805 35.165 ;
        RECT 233.560 34.655 233.820 35.155 ;
        RECT 232.910 34.155 233.310 34.220 ;
        RECT 233.575 34.205 233.805 34.655 ;
        RECT 231.370 33.925 233.370 34.155 ;
        RECT 232.910 33.860 233.310 33.925 ;
        RECT 234.205 33.405 234.855 35.965 ;
        RECT 229.655 32.760 234.855 33.405 ;
        RECT 229.655 30.245 230.430 32.760 ;
        RECT 231.430 32.250 231.830 32.315 ;
        RECT 231.370 32.020 233.370 32.250 ;
        RECT 230.935 31.010 231.165 31.970 ;
        RECT 231.430 31.955 231.830 32.020 ;
        RECT 233.575 31.960 233.805 31.970 ;
        RECT 233.560 31.460 233.820 31.960 ;
        RECT 232.910 30.960 233.310 31.025 ;
        RECT 233.575 31.010 233.805 31.460 ;
        RECT 231.370 30.730 233.370 30.960 ;
        RECT 232.910 30.665 233.310 30.730 ;
        RECT 234.205 30.245 234.855 32.760 ;
        RECT 229.655 29.600 234.855 30.245 ;
        RECT 229.655 27.035 230.430 29.600 ;
        RECT 231.430 29.055 231.830 29.120 ;
        RECT 231.370 28.825 233.370 29.055 ;
        RECT 230.935 27.815 231.165 28.775 ;
        RECT 231.430 28.760 231.830 28.825 ;
        RECT 233.575 28.765 233.805 28.775 ;
        RECT 233.565 28.265 233.825 28.765 ;
        RECT 232.910 27.765 233.310 27.830 ;
        RECT 233.575 27.815 233.805 28.265 ;
        RECT 231.370 27.535 233.370 27.765 ;
        RECT 232.910 27.470 233.310 27.535 ;
        RECT 234.205 27.035 234.855 29.600 ;
        RECT 229.655 26.390 234.855 27.035 ;
        RECT 229.655 23.825 230.430 26.390 ;
        RECT 232.910 25.860 233.310 25.925 ;
        RECT 231.370 25.630 233.370 25.860 ;
        RECT 230.935 24.620 231.165 25.580 ;
        RECT 232.910 25.565 233.310 25.630 ;
        RECT 233.575 25.130 233.805 25.580 ;
        RECT 231.430 24.570 231.830 24.635 ;
        RECT 233.560 24.630 233.820 25.130 ;
        RECT 233.575 24.620 233.805 24.630 ;
        RECT 231.370 24.340 233.370 24.570 ;
        RECT 231.430 24.275 231.830 24.340 ;
        RECT 234.205 23.825 234.855 26.390 ;
        RECT 229.655 23.180 234.855 23.825 ;
        RECT 229.655 20.595 230.430 23.180 ;
        RECT 232.910 22.670 233.310 22.735 ;
        RECT 231.370 22.440 233.370 22.670 ;
        RECT 230.935 21.430 231.165 22.390 ;
        RECT 232.910 22.375 233.310 22.440 ;
        RECT 233.575 21.940 233.805 22.390 ;
        RECT 231.430 21.380 231.830 21.445 ;
        RECT 233.560 21.440 233.820 21.940 ;
        RECT 233.575 21.430 233.805 21.440 ;
        RECT 231.370 21.150 233.370 21.380 ;
        RECT 231.430 21.085 231.830 21.150 ;
        RECT 234.205 20.595 234.855 23.180 ;
        RECT 238.750 22.925 239.415 25.020 ;
        RECT 229.655 20.575 234.855 20.595 ;
        RECT 238.745 20.575 239.415 22.925 ;
        RECT 193.700 20.015 224.560 20.075 ;
        RECT 145.420 18.405 174.550 19.270 ;
        RECT 193.700 18.845 224.590 20.015 ;
        RECT 229.615 19.895 234.860 20.575 ;
        RECT 229.675 19.875 234.800 19.895 ;
        RECT 193.715 18.800 224.460 18.845 ;
        RECT 193.715 18.770 194.495 18.800 ;
        RECT 145.455 18.395 146.230 18.405 ;
        RECT 86.205 17.170 130.240 17.830 ;
        RECT 86.315 17.160 130.160 17.170 ;
        RECT 238.745 13.095 239.410 20.575 ;
        RECT 240.535 20.275 241.045 80.725 ;
        RECT 252.530 80.680 272.635 80.725 ;
        RECT 252.530 80.670 272.520 80.680 ;
        RECT 246.780 80.175 251.780 80.240 ;
        RECT 241.840 79.945 251.840 80.175 ;
        RECT 241.450 79.445 241.680 79.895 ;
        RECT 246.780 79.880 251.780 79.945 ;
        RECT 241.435 78.945 241.695 79.445 ;
        RECT 241.450 78.935 241.680 78.945 ;
        RECT 246.780 78.885 251.780 78.950 ;
        RECT 252.000 78.935 252.230 79.895 ;
        RECT 241.840 78.655 251.840 78.885 ;
        RECT 246.780 78.590 251.780 78.655 ;
        RECT 252.530 78.215 257.175 80.670 ;
        RECT 257.490 78.615 257.760 80.270 ;
        RECT 243.685 78.195 257.175 78.215 ;
        RECT 241.900 76.980 242.300 77.045 ;
        RECT 241.840 76.750 242.840 76.980 ;
        RECT 241.450 76.250 241.680 76.700 ;
        RECT 241.900 76.685 242.300 76.750 ;
        RECT 243.630 76.740 257.175 78.195 ;
        RECT 257.500 78.075 257.750 78.615 ;
        RECT 241.435 75.750 241.695 76.250 ;
        RECT 241.450 75.740 241.680 75.750 ;
        RECT 242.380 75.690 242.780 75.755 ;
        RECT 243.000 75.740 243.230 76.700 ;
        RECT 241.840 75.460 242.840 75.690 ;
        RECT 242.380 75.395 242.780 75.460 ;
        RECT 241.900 73.785 242.300 73.850 ;
        RECT 241.840 73.555 242.840 73.785 ;
        RECT 241.450 73.055 241.680 73.505 ;
        RECT 241.900 73.490 242.300 73.555 ;
        RECT 241.435 72.555 241.695 73.055 ;
        RECT 241.450 72.545 241.680 72.555 ;
        RECT 242.380 72.495 242.780 72.560 ;
        RECT 243.000 72.545 243.230 73.505 ;
        RECT 241.840 72.265 242.840 72.495 ;
        RECT 242.380 72.200 242.780 72.265 ;
        RECT 241.900 70.590 242.300 70.655 ;
        RECT 241.840 70.360 242.840 70.590 ;
        RECT 241.450 69.860 241.680 70.310 ;
        RECT 241.900 70.295 242.300 70.360 ;
        RECT 241.435 69.360 241.695 69.860 ;
        RECT 241.450 69.350 241.680 69.360 ;
        RECT 242.380 69.300 242.780 69.365 ;
        RECT 243.000 69.350 243.230 70.310 ;
        RECT 241.840 69.070 242.840 69.300 ;
        RECT 242.380 69.005 242.780 69.070 ;
        RECT 241.900 67.395 242.300 67.460 ;
        RECT 241.840 67.165 242.840 67.395 ;
        RECT 241.450 66.665 241.680 67.115 ;
        RECT 241.900 67.100 242.300 67.165 ;
        RECT 241.435 66.165 241.695 66.665 ;
        RECT 241.450 66.155 241.680 66.165 ;
        RECT 242.380 66.105 242.780 66.170 ;
        RECT 243.000 66.155 243.230 67.115 ;
        RECT 241.840 65.875 242.840 66.105 ;
        RECT 243.685 66.085 244.865 76.740 ;
        RECT 242.380 65.810 242.780 65.875 ;
        RECT 243.680 64.780 246.590 66.085 ;
        RECT 243.730 64.665 246.510 64.780 ;
        RECT 244.380 64.200 244.780 64.265 ;
        RECT 241.840 63.970 244.840 64.200 ;
        RECT 241.450 63.910 241.680 63.920 ;
        RECT 241.435 63.410 241.695 63.910 ;
        RECT 244.380 63.905 244.780 63.970 ;
        RECT 241.450 62.960 241.680 63.410 ;
        RECT 244.380 62.910 244.780 62.975 ;
        RECT 245.000 62.960 245.230 63.920 ;
        RECT 241.840 62.680 244.840 62.910 ;
        RECT 244.380 62.615 244.780 62.680 ;
        RECT 244.380 61.005 244.780 61.070 ;
        RECT 241.840 60.775 244.840 61.005 ;
        RECT 241.450 60.715 241.680 60.725 ;
        RECT 241.435 60.215 241.695 60.715 ;
        RECT 244.380 60.710 244.780 60.775 ;
        RECT 241.450 59.765 241.680 60.215 ;
        RECT 244.380 59.715 244.780 59.780 ;
        RECT 245.000 59.765 245.230 60.725 ;
        RECT 241.840 59.485 244.840 59.715 ;
        RECT 244.380 59.420 244.780 59.485 ;
        RECT 244.380 57.810 244.780 57.875 ;
        RECT 241.840 57.580 244.840 57.810 ;
        RECT 241.450 57.520 241.680 57.530 ;
        RECT 241.435 57.020 241.695 57.520 ;
        RECT 244.380 57.515 244.780 57.580 ;
        RECT 241.450 56.570 241.680 57.020 ;
        RECT 241.900 56.520 242.300 56.585 ;
        RECT 245.000 56.570 245.230 57.530 ;
        RECT 241.840 56.290 244.840 56.520 ;
        RECT 241.900 56.225 242.300 56.290 ;
        RECT 244.380 54.615 244.780 54.680 ;
        RECT 241.840 54.385 244.840 54.615 ;
        RECT 241.450 54.325 241.680 54.335 ;
        RECT 241.435 53.825 241.695 54.325 ;
        RECT 244.380 54.320 244.780 54.385 ;
        RECT 241.450 53.375 241.680 53.825 ;
        RECT 244.380 53.325 244.780 53.390 ;
        RECT 245.000 53.375 245.230 54.335 ;
        RECT 241.840 53.095 244.840 53.325 ;
        RECT 244.380 53.030 244.780 53.095 ;
        RECT 244.380 51.420 244.780 51.485 ;
        RECT 241.840 51.190 244.840 51.420 ;
        RECT 241.450 51.130 241.680 51.140 ;
        RECT 241.435 50.630 241.695 51.130 ;
        RECT 244.380 51.125 244.780 51.190 ;
        RECT 241.450 50.180 241.680 50.630 ;
        RECT 244.380 50.130 244.780 50.195 ;
        RECT 245.000 50.180 245.230 51.140 ;
        RECT 241.840 49.900 244.840 50.130 ;
        RECT 244.380 49.835 244.780 49.900 ;
        RECT 244.380 48.225 244.780 48.290 ;
        RECT 241.840 47.995 244.840 48.225 ;
        RECT 241.450 47.935 241.680 47.945 ;
        RECT 241.435 47.435 241.695 47.935 ;
        RECT 244.380 47.930 244.780 47.995 ;
        RECT 241.450 46.985 241.680 47.435 ;
        RECT 241.900 46.935 242.300 47.000 ;
        RECT 245.000 46.985 245.230 47.945 ;
        RECT 241.840 46.705 244.840 46.935 ;
        RECT 241.900 46.640 242.300 46.705 ;
        RECT 244.380 45.030 244.780 45.095 ;
        RECT 241.840 44.800 244.840 45.030 ;
        RECT 241.450 44.740 241.680 44.750 ;
        RECT 241.435 44.240 241.695 44.740 ;
        RECT 244.380 44.735 244.780 44.800 ;
        RECT 241.450 43.790 241.680 44.240 ;
        RECT 244.380 43.740 244.780 43.805 ;
        RECT 245.000 43.790 245.230 44.750 ;
        RECT 241.840 43.510 244.840 43.740 ;
        RECT 244.380 43.445 244.780 43.510 ;
        RECT 244.380 41.835 244.780 41.900 ;
        RECT 241.840 41.605 244.840 41.835 ;
        RECT 241.450 41.545 241.680 41.555 ;
        RECT 241.435 41.045 241.695 41.545 ;
        RECT 244.380 41.540 244.780 41.605 ;
        RECT 241.450 40.595 241.680 41.045 ;
        RECT 244.380 40.545 244.780 40.610 ;
        RECT 245.000 40.595 245.230 41.555 ;
        RECT 241.840 40.315 244.840 40.545 ;
        RECT 244.380 40.250 244.780 40.315 ;
        RECT 244.380 38.640 244.780 38.705 ;
        RECT 241.840 38.410 244.840 38.640 ;
        RECT 241.450 38.350 241.680 38.360 ;
        RECT 241.435 37.850 241.695 38.350 ;
        RECT 244.380 38.345 244.780 38.410 ;
        RECT 241.450 37.400 241.680 37.850 ;
        RECT 241.900 37.350 242.300 37.415 ;
        RECT 245.000 37.400 245.230 38.360 ;
        RECT 241.840 37.120 244.840 37.350 ;
        RECT 241.900 37.055 242.300 37.120 ;
        RECT 244.380 35.445 244.780 35.510 ;
        RECT 241.840 35.215 244.840 35.445 ;
        RECT 241.450 35.155 241.680 35.165 ;
        RECT 241.435 34.655 241.695 35.155 ;
        RECT 244.380 35.150 244.780 35.215 ;
        RECT 241.450 34.205 241.680 34.655 ;
        RECT 244.380 34.155 244.780 34.220 ;
        RECT 245.000 34.205 245.230 35.165 ;
        RECT 241.840 33.925 244.840 34.155 ;
        RECT 244.380 33.860 244.780 33.925 ;
        RECT 244.380 32.250 244.780 32.315 ;
        RECT 241.840 32.020 244.840 32.250 ;
        RECT 241.450 31.960 241.680 31.970 ;
        RECT 241.435 31.460 241.695 31.960 ;
        RECT 244.380 31.955 244.780 32.020 ;
        RECT 241.450 31.010 241.680 31.460 ;
        RECT 244.380 30.960 244.780 31.025 ;
        RECT 245.000 31.010 245.230 31.970 ;
        RECT 241.840 30.730 244.840 30.960 ;
        RECT 244.380 30.665 244.780 30.730 ;
        RECT 244.380 29.055 244.780 29.120 ;
        RECT 241.840 28.825 244.840 29.055 ;
        RECT 241.450 28.765 241.680 28.775 ;
        RECT 241.435 28.265 241.695 28.765 ;
        RECT 244.380 28.760 244.780 28.825 ;
        RECT 241.450 27.815 241.680 28.265 ;
        RECT 241.900 27.765 242.300 27.830 ;
        RECT 245.000 27.815 245.230 28.775 ;
        RECT 241.840 27.535 244.840 27.765 ;
        RECT 241.900 27.470 242.300 27.535 ;
        RECT 245.505 27.065 246.510 64.665 ;
        RECT 243.695 27.050 246.555 27.065 ;
        RECT 241.900 25.860 242.300 25.925 ;
        RECT 241.840 25.630 242.840 25.860 ;
        RECT 243.610 25.680 246.555 27.050 ;
        RECT 241.450 25.130 241.680 25.580 ;
        RECT 241.900 25.565 242.300 25.630 ;
        RECT 241.435 24.630 241.695 25.130 ;
        RECT 241.450 24.620 241.680 24.630 ;
        RECT 242.380 24.570 242.780 24.635 ;
        RECT 243.000 24.620 243.230 25.580 ;
        RECT 241.840 24.340 242.840 24.570 ;
        RECT 242.380 24.275 242.780 24.340 ;
        RECT 241.915 22.670 242.315 22.735 ;
        RECT 241.855 22.440 242.855 22.670 ;
        RECT 241.465 21.940 241.695 22.390 ;
        RECT 241.915 22.375 242.315 22.440 ;
        RECT 241.450 21.440 241.710 21.940 ;
        RECT 241.465 21.430 241.695 21.440 ;
        RECT 242.395 21.380 242.795 21.445 ;
        RECT 243.015 21.430 243.245 22.390 ;
        RECT 241.855 21.150 242.855 21.380 ;
        RECT 242.395 21.085 242.795 21.150 ;
        RECT 243.610 20.280 244.865 25.680 ;
        RECT 256.220 20.475 257.175 76.740 ;
        RECT 257.500 52.845 257.750 53.235 ;
        RECT 257.490 51.190 257.760 52.845 ;
        RECT 257.500 51.130 257.750 51.190 ;
        RECT 257.490 48.325 257.760 49.980 ;
        RECT 257.500 47.835 257.750 48.325 ;
        RECT 257.500 22.555 257.750 22.995 ;
        RECT 257.490 20.900 257.760 22.555 ;
        RECT 257.500 20.890 257.750 20.900 ;
        RECT 258.045 20.475 258.615 80.670 ;
        RECT 258.970 78.615 259.240 80.270 ;
        RECT 258.980 78.075 259.230 78.615 ;
        RECT 258.980 52.845 259.230 53.235 ;
        RECT 258.970 51.190 259.240 52.845 ;
        RECT 258.980 51.130 259.230 51.190 ;
        RECT 258.970 48.325 259.240 49.980 ;
        RECT 258.980 47.835 259.230 48.325 ;
        RECT 258.980 22.555 259.230 22.995 ;
        RECT 258.970 20.900 259.240 22.555 ;
        RECT 258.980 20.890 259.230 20.900 ;
        RECT 259.530 20.475 260.100 80.670 ;
        RECT 260.450 78.615 260.720 80.270 ;
        RECT 260.460 78.075 260.710 78.615 ;
        RECT 260.460 52.845 260.710 53.235 ;
        RECT 260.450 51.190 260.720 52.845 ;
        RECT 260.460 51.130 260.710 51.190 ;
        RECT 260.450 48.325 260.720 49.980 ;
        RECT 260.460 47.835 260.710 48.325 ;
        RECT 260.460 22.555 260.710 22.995 ;
        RECT 260.450 20.900 260.720 22.555 ;
        RECT 260.460 20.890 260.710 20.900 ;
        RECT 261.200 20.475 261.810 80.670 ;
        RECT 256.220 20.280 261.810 20.475 ;
        RECT 243.610 20.275 261.810 20.280 ;
        RECT 240.535 19.335 261.810 20.275 ;
        RECT 240.535 19.325 240.780 19.335 ;
        RECT 261.200 19.315 261.810 19.335 ;
        RECT 238.695 12.430 239.465 13.095 ;
      LAYER met2 ;
        RECT 14.810 214.365 31.790 215.620 ;
        RECT 14.810 154.025 16.085 214.365 ;
        RECT 30.660 157.630 31.720 214.365 ;
        RECT 32.805 158.220 57.060 159.245 ;
        RECT 16.565 154.460 16.925 156.560 ;
        RECT 33.765 156.545 34.025 156.880 ;
        RECT 55.655 156.660 55.975 157.260 ;
        RECT 29.940 156.245 34.025 156.545 ;
        RECT 29.940 154.460 30.200 156.245 ;
        RECT 34.120 155.740 35.385 156.125 ;
        RECT 53.790 155.695 55.590 156.160 ;
        RECT 56.440 155.410 57.015 158.220 ;
        RECT 32.800 154.720 57.055 155.410 ;
        RECT 32.800 154.525 57.090 154.720 ;
        RECT 32.800 154.385 57.095 154.525 ;
        RECT 11.440 153.980 16.085 154.025 ;
        RECT 11.440 152.945 31.720 153.980 ;
        RECT 11.440 152.935 14.920 152.945 ;
        RECT 55.075 146.940 57.095 154.385 ;
        RECT 55.075 144.920 57.140 146.940 ;
        RECT 57.495 141.520 60.120 141.550 ;
        RECT 11.465 138.895 60.120 141.520 ;
        RECT 57.495 138.865 60.120 138.895 ;
        RECT 96.515 138.835 96.915 138.885 ;
        RECT 90.890 138.475 96.915 138.835 ;
        RECT 96.515 136.415 96.915 138.475 ;
        RECT 103.475 129.615 106.120 130.145 ;
        RECT 91.375 125.155 92.875 125.515 ;
        RECT 55.295 122.865 56.490 122.900 ;
        RECT 55.295 122.790 82.745 122.865 ;
        RECT 55.295 120.715 90.805 122.790 ;
        RECT 55.295 120.685 82.745 120.715 ;
        RECT 26.885 44.930 27.705 120.380 ;
        RECT 55.295 98.580 56.490 120.685 ;
        RECT 57.485 120.305 57.785 120.345 ;
        RECT 57.485 120.085 60.135 120.305 ;
        RECT 57.485 119.945 57.785 120.085 ;
        RECT 59.835 119.945 60.135 120.085 ;
        RECT 62.345 120.085 67.425 120.395 ;
        RECT 62.345 120.035 62.645 120.085 ;
        RECT 64.775 120.035 65.075 120.085 ;
        RECT 67.125 120.035 67.425 120.085 ;
        RECT 69.635 120.085 72.285 120.395 ;
        RECT 69.635 120.035 69.935 120.085 ;
        RECT 71.985 120.035 72.285 120.085 ;
        RECT 74.495 120.085 77.145 120.395 ;
        RECT 74.495 120.035 74.795 120.085 ;
        RECT 76.845 120.035 77.145 120.085 ;
        RECT 79.355 120.035 79.655 120.685 ;
        RECT 57.985 119.550 58.245 119.600 ;
        RECT 59.375 119.550 59.635 119.600 ;
        RECT 57.985 119.045 59.635 119.550 ;
        RECT 57.985 114.500 58.245 119.045 ;
        RECT 59.375 114.500 59.635 119.045 ;
        RECT 60.425 119.560 60.685 119.600 ;
        RECT 61.815 119.560 62.075 119.610 ;
        RECT 60.425 119.055 62.075 119.560 ;
        RECT 60.425 114.500 60.685 119.055 ;
        RECT 61.815 114.510 62.075 119.055 ;
        RECT 65.270 119.575 65.530 119.625 ;
        RECT 66.665 119.575 66.925 119.625 ;
        RECT 65.270 119.070 66.925 119.575 ;
        RECT 65.270 114.525 65.530 119.070 ;
        RECT 66.665 114.525 66.925 119.070 ;
        RECT 67.710 119.565 67.970 119.615 ;
        RECT 69.085 119.565 69.345 119.615 ;
        RECT 67.710 119.060 69.345 119.565 ;
        RECT 67.710 114.515 67.970 119.060 ;
        RECT 69.085 114.515 69.345 119.060 ;
        RECT 70.145 119.560 70.405 119.610 ;
        RECT 71.520 119.560 71.780 119.610 ;
        RECT 70.145 119.055 71.780 119.560 ;
        RECT 70.145 114.510 70.405 119.055 ;
        RECT 71.520 114.510 71.780 119.055 ;
        RECT 72.570 119.565 72.830 119.610 ;
        RECT 73.950 119.565 74.210 119.610 ;
        RECT 72.570 119.060 74.210 119.565 ;
        RECT 75.005 119.560 75.265 119.610 ;
        RECT 76.380 119.560 76.640 119.610 ;
        RECT 72.570 114.510 72.830 119.060 ;
        RECT 73.950 114.510 74.210 119.060 ;
        RECT 74.995 119.055 76.640 119.560 ;
        RECT 75.005 114.510 75.265 119.055 ;
        RECT 76.380 114.510 76.640 119.055 ;
        RECT 77.430 119.605 77.690 119.610 ;
        RECT 78.815 119.605 79.075 119.610 ;
        RECT 77.430 119.100 79.075 119.605 ;
        RECT 77.430 114.510 77.690 119.100 ;
        RECT 78.815 114.510 79.075 119.100 ;
        RECT 92.375 117.830 92.875 125.155 ;
        RECT 104.405 120.030 127.170 120.040 ;
        RECT 104.405 118.640 127.330 120.030 ;
        RECT 125.070 118.635 127.330 118.640 ;
        RECT 80.700 117.330 105.785 117.830 ;
        RECT 80.700 104.990 81.100 117.330 ;
        RECT 105.525 116.730 105.785 117.330 ;
        RECT 125.815 117.230 126.075 117.830 ;
        RECT 125.815 116.730 128.750 117.230 ;
        RECT 83.245 113.350 83.505 113.950 ;
        RECT 81.860 112.850 83.505 113.350 ;
        RECT 103.525 113.350 103.805 113.950 ;
        RECT 103.525 112.850 127.640 113.350 ;
        RECT 81.860 109.520 82.360 112.850 ;
        RECT 83.345 110.555 102.215 111.575 ;
        RECT 107.320 110.425 126.790 111.700 ;
        RECT 81.860 109.470 82.630 109.520 ;
        RECT 127.140 109.470 127.640 112.850 ;
        RECT 81.860 108.970 105.785 109.470 ;
        RECT 82.130 108.920 82.630 108.970 ;
        RECT 83.280 104.990 83.540 105.590 ;
        RECT 80.700 104.490 83.540 104.990 ;
        RECT 82.980 103.175 101.730 103.710 ;
        RECT 102.110 101.200 102.490 108.970 ;
        RECT 104.235 105.730 105.015 108.635 ;
        RECT 105.525 108.370 105.785 108.970 ;
        RECT 125.815 108.970 127.640 109.470 ;
        RECT 125.815 108.370 126.075 108.970 ;
        RECT 126.390 105.730 127.325 108.555 ;
        RECT 103.570 104.990 103.830 105.590 ;
        RECT 104.235 105.500 127.325 105.730 ;
        RECT 104.270 105.245 127.325 105.500 ;
        RECT 127.220 104.990 127.720 105.040 ;
        RECT 128.250 104.990 128.750 116.730 ;
        RECT 103.570 104.490 128.750 104.990 ;
        RECT 127.220 104.440 127.720 104.490 ;
        RECT 102.110 100.820 131.520 101.200 ;
        RECT 57.485 98.230 57.785 100.045 ;
        RECT 59.915 99.965 60.215 100.015 ;
        RECT 62.265 99.965 62.565 100.015 ;
        RECT 59.915 99.655 62.565 99.965 ;
        RECT 57.430 97.630 57.815 98.230 ;
        RECT 34.090 97.055 34.900 97.130 ;
        RECT 64.695 97.055 64.995 100.015 ;
        RECT 67.205 99.965 67.505 100.015 ;
        RECT 69.555 99.965 69.855 100.015 ;
        RECT 67.205 99.655 69.855 99.965 ;
        RECT 72.065 99.965 72.365 100.015 ;
        RECT 74.415 99.965 74.715 100.015 ;
        RECT 72.065 99.655 74.715 99.965 ;
        RECT 76.925 99.965 77.225 100.015 ;
        RECT 79.275 99.965 79.575 100.015 ;
        RECT 76.925 99.655 79.575 99.965 ;
        RECT 34.090 96.795 64.995 97.055 ;
        RECT 34.090 50.965 34.900 96.795 ;
        RECT 58.330 90.830 58.590 96.795 ;
        RECT 73.335 95.130 78.335 95.510 ;
        RECT 84.115 95.130 89.115 95.510 ;
        RECT 58.295 86.890 58.615 87.990 ;
        RECT 44.435 74.120 73.685 74.480 ;
        RECT 66.855 73.390 67.815 73.740 ;
        RECT 68.330 73.390 68.590 73.725 ;
        RECT 66.855 72.990 68.590 73.390 ;
        RECT 78.620 73.410 78.880 94.990 ;
        RECT 125.660 91.890 125.980 94.990 ;
        RECT 131.140 93.335 131.520 100.820 ;
        RECT 133.600 93.355 134.100 93.775 ;
        RECT 131.760 88.195 132.040 93.295 ;
        RECT 217.340 93.230 238.120 93.625 ;
        RECT 83.740 85.010 84.060 88.110 ;
        RECT 134.280 87.985 134.560 93.085 ;
        RECT 83.740 79.870 84.060 82.970 ;
        RECT 104.060 80.370 104.320 87.610 ;
        RECT 105.400 80.370 105.660 87.610 ;
        RECT 217.340 81.450 217.735 93.230 ;
        RECT 237.725 92.020 238.120 93.230 ;
        RECT 244.650 92.305 261.660 92.630 ;
        RECT 244.650 92.300 259.700 92.305 ;
        RECT 237.705 91.675 238.140 92.020 ;
        RECT 237.725 91.650 238.120 91.675 ;
        RECT 244.650 89.775 244.910 92.300 ;
        RECT 260.615 89.940 261.660 92.305 ;
        RECT 270.650 90.450 271.695 92.630 ;
        RECT 270.650 89.940 273.120 90.450 ;
        RECT 271.650 89.935 273.120 89.940 ;
        RECT 242.230 89.515 244.910 89.775 ;
        RECT 241.385 88.880 241.745 88.980 ;
        RECT 235.415 88.580 241.745 88.880 ;
        RECT 195.235 81.055 217.735 81.450 ;
        RECT 104.060 73.410 104.320 74.045 ;
        RECT 105.400 73.410 105.660 74.045 ;
        RECT 125.660 73.795 125.980 76.090 ;
        RECT 125.610 73.635 126.030 73.795 ;
        RECT 78.620 72.990 134.235 73.410 ;
        RECT 66.855 72.115 67.815 72.990 ;
        RECT 66.855 72.050 135.695 72.115 ;
        RECT 136.865 72.050 139.745 72.100 ;
        RECT 66.855 71.945 139.745 72.050 ;
        RECT 66.865 71.605 139.745 71.945 ;
        RECT 59.625 70.045 139.745 71.605 ;
        RECT 59.625 69.650 135.695 70.045 ;
        RECT 136.865 69.995 139.745 70.045 ;
        RECT 59.625 69.600 67.535 69.650 ;
        RECT 59.635 59.600 63.415 69.600 ;
        RECT 76.255 59.965 77.580 69.650 ;
        RECT 72.410 59.950 78.030 59.965 ;
        RECT 59.635 59.510 63.420 59.600 ;
        RECT 48.365 58.960 63.430 59.510 ;
        RECT 72.250 59.310 78.030 59.950 ;
        RECT 48.365 58.500 63.420 58.960 ;
        RECT 48.365 57.885 63.260 58.500 ;
        RECT 49.685 55.965 49.945 57.885 ;
        RECT 37.870 55.450 53.585 55.810 ;
        RECT 38.545 54.095 59.740 55.235 ;
        RECT 38.545 51.260 39.280 54.095 ;
        RECT 39.620 51.150 39.975 53.130 ;
        RECT 59.975 51.410 60.235 56.945 ;
        RECT 58.215 51.150 60.235 51.410 ;
        RECT 34.090 50.605 45.040 50.965 ;
        RECT 34.090 50.600 38.180 50.605 ;
        RECT 34.090 50.595 34.900 50.600 ;
        RECT 38.565 49.490 57.925 50.170 ;
        RECT 40.215 46.920 40.535 48.200 ;
        RECT 43.825 45.140 44.290 46.360 ;
        RECT 47.585 45.720 47.905 47.000 ;
        RECT 40.540 44.930 41.040 44.980 ;
        RECT 45.220 44.930 45.720 44.980 ;
        RECT 26.885 44.430 45.720 44.930 ;
        RECT 40.540 44.380 41.040 44.430 ;
        RECT 45.220 44.380 45.720 44.430 ;
        RECT 30.925 44.180 31.965 44.230 ;
        RECT 42.400 44.180 42.900 44.230 ;
        RECT 47.110 44.180 47.610 44.230 ;
        RECT 30.910 43.680 47.610 44.180 ;
        RECT 30.925 43.625 31.965 43.680 ;
        RECT 42.400 43.630 42.900 43.680 ;
        RECT 47.110 43.630 47.610 43.680 ;
        RECT 40.215 40.510 40.535 41.790 ;
        RECT 47.585 41.715 47.905 42.990 ;
        RECT 48.300 39.745 49.075 49.490 ;
        RECT 38.715 39.125 49.165 39.745 ;
        RECT 53.425 39.705 54.115 49.490 ;
        RECT 58.215 49.250 58.545 51.150 ;
        RECT 60.785 49.320 63.260 57.885 ;
        RECT 72.250 56.300 72.845 59.310 ;
        RECT 70.590 55.465 70.960 55.470 ;
        RECT 70.590 55.460 72.175 55.465 ;
        RECT 73.130 55.460 73.390 58.265 ;
        RECT 74.710 58.045 74.970 59.310 ;
        RECT 73.665 56.075 74.040 56.105 ;
        RECT 76.290 56.075 76.550 58.265 ;
        RECT 76.875 56.370 77.515 59.310 ;
        RECT 73.665 55.805 93.725 56.075 ;
        RECT 73.665 55.775 74.040 55.805 ;
        RECT 74.615 55.460 74.980 55.490 ;
        RECT 70.590 55.190 74.980 55.460 ;
        RECT 69.215 50.815 69.560 53.870 ;
        RECT 73.620 52.575 73.880 55.190 ;
        RECT 74.615 55.160 74.980 55.190 ;
        RECT 70.245 52.570 73.880 52.575 ;
        RECT 70.050 52.315 73.880 52.570 ;
        RECT 70.050 52.070 70.310 52.315 ;
        RECT 70.840 51.870 71.100 52.090 ;
        RECT 72.830 51.870 73.090 52.090 ;
        RECT 73.620 52.070 73.880 52.315 ;
        RECT 75.610 52.570 75.870 55.805 ;
        RECT 75.610 52.310 79.440 52.570 ;
        RECT 75.610 52.070 75.870 52.310 ;
        RECT 70.840 51.640 73.090 51.870 ;
        RECT 70.840 50.815 71.100 51.640 ;
        RECT 72.830 51.590 73.090 51.640 ;
        RECT 76.400 51.820 76.660 52.090 ;
        RECT 78.390 51.820 78.650 52.090 ;
        RECT 79.180 52.070 79.440 52.310 ;
        RECT 76.400 51.590 78.650 51.820 ;
        RECT 73.185 51.060 73.525 51.440 ;
        RECT 76.400 50.815 76.660 51.590 ;
        RECT 78.745 51.060 79.085 51.440 ;
        RECT 79.930 50.815 80.250 53.880 ;
        RECT 69.215 50.715 80.250 50.815 ;
        RECT 69.215 50.685 80.240 50.715 ;
        RECT 69.160 50.145 80.240 50.685 ;
        RECT 57.265 48.990 59.495 49.250 ;
        RECT 54.545 45.810 54.865 46.910 ;
        RECT 54.545 41.765 54.865 42.865 ;
        RECT 57.265 41.765 57.525 48.990 ;
        RECT 59.235 41.765 59.495 48.990 ;
        RECT 61.895 47.190 62.215 48.290 ;
        RECT 61.895 40.385 62.215 41.485 ;
        RECT 62.640 39.705 63.245 49.320 ;
        RECT 53.425 38.995 63.245 39.705 ;
        RECT 53.470 38.975 63.245 38.995 ;
        RECT 62.640 38.930 63.245 38.975 ;
        RECT 51.980 38.590 52.310 38.640 ;
        RECT 35.955 38.540 52.310 38.590 ;
        RECT 35.840 38.520 52.310 38.540 ;
        RECT 35.840 38.500 63.315 38.520 ;
        RECT 69.195 38.500 70.510 50.145 ;
        RECT 86.225 49.890 92.840 50.500 ;
        RECT 35.840 38.110 70.510 38.500 ;
        RECT 35.840 38.090 52.310 38.110 ;
        RECT 35.840 35.435 36.240 38.090 ;
        RECT 36.615 36.905 36.935 37.325 ;
        RECT 42.935 36.725 43.195 38.090 ;
        RECT 44.925 36.725 45.185 38.090 ;
        RECT 51.185 36.345 51.505 36.765 ;
        RECT 51.980 35.435 52.310 38.090 ;
        RECT 35.840 35.365 52.310 35.435 ;
        RECT 53.485 35.365 54.170 38.110 ;
        RECT 54.545 36.725 54.865 37.325 ;
        RECT 54.930 35.825 55.730 36.245 ;
        RECT 57.065 35.365 57.325 36.945 ;
        RECT 57.885 35.365 58.850 38.110 ;
        RECT 59.435 36.730 59.695 38.110 ;
        RECT 61.895 36.730 62.215 37.330 ;
        RECT 62.690 37.305 70.510 38.110 ;
        RECT 59.790 35.835 60.590 36.255 ;
        RECT 62.690 35.365 63.315 37.305 ;
        RECT 35.840 34.955 63.375 35.365 ;
        RECT 35.840 34.635 52.310 34.955 ;
        RECT 35.840 31.865 36.240 34.635 ;
        RECT 36.615 33.325 36.935 33.745 ;
        RECT 42.935 31.865 43.195 33.365 ;
        RECT 44.925 31.865 45.185 33.365 ;
        RECT 51.185 32.710 51.505 33.130 ;
        RECT 51.980 31.865 52.310 34.635 ;
        RECT 35.840 31.065 52.310 31.865 ;
        RECT 35.840 28.210 36.240 31.065 ;
        RECT 36.615 29.745 36.935 30.165 ;
        RECT 42.935 28.210 43.195 29.785 ;
        RECT 44.925 28.210 45.185 29.785 ;
        RECT 51.185 29.745 51.505 30.165 ;
        RECT 51.980 28.210 52.310 31.065 ;
        RECT 35.840 27.410 52.310 28.210 ;
        RECT 35.840 24.725 36.240 27.410 ;
        RECT 36.615 25.605 36.935 26.025 ;
        RECT 42.935 24.725 43.195 26.205 ;
        RECT 44.925 24.725 45.185 26.205 ;
        RECT 51.185 26.165 51.505 26.585 ;
        RECT 51.980 24.725 52.310 27.410 ;
        RECT 35.840 24.465 52.310 24.725 ;
        RECT 35.725 23.925 52.310 24.465 ;
        RECT 38.670 20.920 44.060 23.925 ;
        RECT 51.980 23.890 52.310 23.925 ;
        RECT 86.265 31.315 91.850 49.890 ;
        RECT 93.045 48.285 93.725 55.805 ;
        RECT 104.560 50.350 130.230 50.355 ;
        RECT 93.985 49.740 130.230 50.350 ;
        RECT 100.925 48.815 103.025 49.075 ;
        RECT 93.045 48.025 95.145 48.285 ;
        RECT 93.045 46.705 93.725 48.025 ;
        RECT 102.345 47.495 103.025 48.815 ;
        RECT 100.925 47.235 103.025 47.495 ;
        RECT 93.045 46.445 95.145 46.705 ;
        RECT 93.045 45.125 93.725 46.445 ;
        RECT 102.345 45.915 103.025 47.235 ;
        RECT 100.925 45.655 103.025 45.915 ;
        RECT 93.045 44.865 95.145 45.125 ;
        RECT 93.045 43.545 93.725 44.865 ;
        RECT 102.345 44.335 103.025 45.655 ;
        RECT 100.925 44.075 103.025 44.335 ;
        RECT 93.045 43.285 95.145 43.545 ;
        RECT 93.045 41.965 93.725 43.285 ;
        RECT 102.345 42.755 103.025 44.075 ;
        RECT 100.925 42.495 103.025 42.755 ;
        RECT 93.045 41.705 95.145 41.965 ;
        RECT 93.045 40.385 93.725 41.705 ;
        RECT 102.345 41.175 103.025 42.495 ;
        RECT 100.925 40.915 103.025 41.175 ;
        RECT 93.045 40.125 95.145 40.385 ;
        RECT 93.045 38.805 93.725 40.125 ;
        RECT 102.345 39.595 103.025 40.915 ;
        RECT 104.205 48.930 130.230 49.740 ;
        RECT 104.205 40.150 105.310 48.930 ;
        RECT 108.620 45.915 109.640 48.930 ;
        RECT 126.230 46.445 128.490 46.800 ;
        RECT 108.620 41.030 109.635 45.915 ;
        RECT 126.230 42.005 128.490 42.355 ;
        RECT 129.525 41.555 130.230 48.930 ;
        RECT 132.030 40.735 132.290 69.650 ;
        RECT 195.235 69.645 195.705 81.055 ;
        RECT 229.590 78.480 232.970 82.260 ;
        RECT 229.570 78.130 232.970 78.480 ;
        RECT 228.445 78.090 232.970 78.130 ;
        RECT 228.445 77.470 234.795 78.090 ;
        RECT 228.445 75.705 230.450 77.470 ;
        RECT 235.415 76.995 235.865 88.580 ;
        RECT 243.590 88.485 244.295 88.825 ;
        RECT 242.230 88.225 244.295 88.485 ;
        RECT 272.760 88.230 273.120 89.935 ;
        RECT 243.590 87.015 244.295 88.225 ;
        RECT 245.490 87.950 267.195 88.225 ;
        RECT 270.860 87.950 273.120 88.230 ;
        RECT 245.490 87.945 264.910 87.950 ;
        RECT 245.490 86.580 245.750 87.945 ;
        RECT 242.230 86.320 245.750 86.580 ;
        RECT 272.760 86.160 273.120 87.950 ;
        RECT 246.730 85.900 248.195 86.160 ;
        RECT 270.075 85.900 273.120 86.160 ;
        RECT 241.385 85.685 241.745 85.785 ;
        RECT 236.425 85.385 241.745 85.685 ;
        RECT 243.610 85.290 244.315 85.855 ;
        RECT 242.230 85.030 244.315 85.290 ;
        RECT 243.610 84.435 244.315 85.030 ;
        RECT 243.610 84.345 246.150 84.435 ;
        RECT 243.635 83.880 246.150 84.345 ;
        RECT 246.730 83.385 247.095 85.900 ;
        RECT 247.400 83.900 253.305 84.460 ;
        RECT 246.730 83.125 251.830 83.385 ;
        RECT 241.385 82.490 241.745 82.590 ;
        RECT 238.490 82.190 241.745 82.490 ;
        RECT 252.535 82.095 253.305 83.900 ;
        RECT 246.730 81.835 253.305 82.095 ;
        RECT 252.535 80.765 253.305 81.835 ;
        RECT 272.760 80.220 273.120 85.900 ;
        RECT 246.730 79.930 254.865 80.220 ;
        RECT 241.385 79.295 241.745 79.395 ;
        RECT 239.880 78.995 241.745 79.295 ;
        RECT 252.510 78.900 253.260 79.230 ;
        RECT 246.730 78.640 253.260 78.900 ;
        RECT 252.510 78.165 253.260 78.640 ;
        RECT 243.635 77.420 253.260 78.165 ;
        RECT 232.865 76.735 242.350 76.995 ;
        RECT 233.515 76.090 233.875 76.200 ;
        RECT 237.675 76.090 238.175 76.135 ;
        RECT 241.385 76.090 241.745 76.200 ;
        RECT 233.380 75.800 241.745 76.090 ;
        RECT 243.635 75.705 244.690 77.420 ;
        RECT 228.445 75.445 231.885 75.705 ;
        RECT 242.330 75.445 244.690 75.705 ;
        RECT 228.445 72.510 230.450 75.445 ;
        RECT 236.450 73.800 236.950 73.940 ;
        RECT 232.865 73.540 242.350 73.800 ;
        RECT 233.515 72.895 233.875 73.005 ;
        RECT 235.885 72.895 236.335 72.915 ;
        RECT 241.385 72.895 241.745 73.005 ;
        RECT 233.400 72.605 241.745 72.895 ;
        RECT 243.635 72.510 244.690 75.445 ;
        RECT 228.445 72.250 231.885 72.510 ;
        RECT 242.330 72.250 244.690 72.510 ;
        RECT 195.215 69.225 195.725 69.645 ;
        RECT 228.445 69.315 230.450 72.250 ;
        RECT 238.515 70.605 238.965 70.695 ;
        RECT 232.865 70.345 242.350 70.605 ;
        RECT 233.515 69.700 233.875 69.810 ;
        RECT 238.525 69.700 238.975 69.790 ;
        RECT 241.385 69.700 241.745 69.810 ;
        RECT 233.385 69.410 241.745 69.700 ;
        RECT 238.525 69.380 238.975 69.410 ;
        RECT 243.635 69.315 244.690 72.250 ;
        RECT 195.235 69.200 195.705 69.225 ;
        RECT 228.445 69.055 231.885 69.315 ;
        RECT 242.330 69.055 244.690 69.315 ;
        RECT 228.445 68.920 230.450 69.055 ;
        RECT 192.975 67.495 230.450 68.920 ;
        RECT 192.980 57.185 194.520 67.495 ;
        RECT 195.290 66.800 195.800 67.195 ;
        RECT 196.190 66.635 196.590 67.495 ;
        RECT 198.750 66.635 199.150 67.495 ;
        RECT 201.340 66.635 201.740 67.495 ;
        RECT 203.930 66.635 204.330 67.495 ;
        RECT 206.515 66.635 206.915 67.495 ;
        RECT 207.320 67.165 210.590 67.185 ;
        RECT 207.320 66.805 210.595 67.165 ;
        RECT 207.320 66.790 210.590 66.805 ;
        RECT 207.335 66.780 207.800 66.790 ;
        RECT 211.070 66.635 211.470 67.495 ;
        RECT 213.610 66.635 214.010 67.495 ;
        RECT 216.195 66.635 216.595 67.495 ;
        RECT 218.725 66.635 219.125 67.495 ;
        RECT 221.230 66.635 221.630 67.495 ;
        RECT 196.190 66.200 221.630 66.635 ;
        RECT 196.190 62.560 196.450 66.200 ;
        RECT 198.805 62.560 199.065 66.200 ;
        RECT 201.375 62.520 201.635 66.200 ;
        RECT 203.980 62.520 204.240 66.200 ;
        RECT 206.560 62.500 206.820 66.200 ;
        RECT 165.430 55.870 194.520 57.185 ;
        RECT 165.430 51.605 166.205 55.870 ;
        RECT 167.110 55.140 167.630 55.535 ;
        RECT 168.035 54.960 168.345 55.870 ;
        RECT 170.615 54.960 170.925 55.870 ;
        RECT 173.190 54.960 173.500 55.870 ;
        RECT 175.785 54.960 176.095 55.870 ;
        RECT 178.340 54.960 178.650 55.870 ;
        RECT 168.035 54.645 178.650 54.960 ;
        RECT 168.035 54.485 178.625 54.645 ;
        RECT 145.085 50.170 159.255 51.325 ;
        RECT 161.310 50.525 166.205 51.605 ;
        RECT 168.040 50.855 168.300 54.485 ;
        RECT 170.625 50.860 170.885 54.485 ;
        RECT 173.205 50.860 173.465 54.485 ;
        RECT 175.785 50.855 176.045 54.485 ;
        RECT 178.365 50.860 178.625 54.485 ;
        RECT 152.310 49.545 162.650 49.905 ;
        RECT 164.410 49.690 166.205 50.525 ;
        RECT 162.390 47.475 162.650 49.545 ;
        RECT 163.670 49.200 166.205 49.690 ;
        RECT 163.670 47.590 163.975 49.200 ;
        RECT 162.380 45.710 162.665 47.475 ;
        RECT 164.410 44.955 166.205 49.200 ;
        RECT 166.755 45.420 167.015 49.075 ;
        RECT 169.335 45.420 169.595 49.075 ;
        RECT 171.915 45.420 172.175 49.075 ;
        RECT 174.495 45.420 174.755 49.075 ;
        RECT 177.075 45.420 177.335 49.075 ;
        RECT 179.655 45.420 179.915 49.075 ;
        RECT 166.755 44.975 179.915 45.420 ;
        RECT 161.390 44.240 166.205 44.955 ;
        RECT 165.430 43.995 166.205 44.240 ;
        RECT 165.430 43.555 170.275 43.995 ;
        RECT 115.510 40.475 132.290 40.735 ;
        RECT 165.385 42.825 170.275 43.555 ;
        RECT 100.925 39.335 103.025 39.595 ;
        RECT 93.040 38.545 95.140 38.805 ;
        RECT 93.045 37.225 93.725 38.545 ;
        RECT 102.345 38.015 103.025 39.335 ;
        RECT 115.510 39.105 115.770 40.475 ;
        RECT 129.505 39.480 130.210 40.045 ;
        RECT 132.030 39.105 132.290 40.475 ;
        RECT 147.430 40.255 152.430 40.615 ;
        RECT 113.140 38.845 115.770 39.105 ;
        RECT 125.500 38.845 132.290 39.105 ;
        RECT 147.435 38.705 147.950 40.255 ;
        RECT 115.785 38.640 116.145 38.660 ;
        RECT 100.925 37.755 103.025 38.015 ;
        RECT 93.045 36.965 95.145 37.225 ;
        RECT 93.045 35.645 93.725 36.965 ;
        RECT 102.345 36.435 103.025 37.755 ;
        RECT 100.925 36.175 103.025 36.435 ;
        RECT 93.045 35.385 95.145 35.645 ;
        RECT 93.045 34.065 93.725 35.385 ;
        RECT 102.345 34.855 103.025 36.175 ;
        RECT 100.925 34.595 103.025 34.855 ;
        RECT 105.495 34.770 105.855 38.640 ;
        RECT 115.770 37.760 116.160 38.640 ;
        RECT 115.785 37.700 116.145 37.760 ;
        RECT 93.045 33.805 95.145 34.065 ;
        RECT 93.045 32.485 93.725 33.805 ;
        RECT 102.345 33.275 103.025 34.595 ;
        RECT 100.925 33.015 103.025 33.275 ;
        RECT 93.045 32.225 95.145 32.485 ;
        RECT 86.265 17.785 87.205 31.315 ;
        RECT 93.045 29.805 93.725 32.225 ;
        RECT 102.345 31.695 103.025 33.015 ;
        RECT 105.495 31.695 105.855 32.840 ;
        RECT 115.785 31.900 116.145 35.810 ;
        RECT 117.805 34.730 118.165 38.640 ;
        RECT 128.080 37.760 128.470 38.640 ;
        RECT 128.095 37.700 128.455 37.760 ;
        RECT 100.925 31.435 105.855 31.695 ;
        RECT 93.045 29.100 107.610 29.805 ;
        RECT 117.805 29.635 118.165 32.875 ;
        RECT 128.095 31.900 128.455 35.790 ;
        RECT 129.505 32.915 130.210 38.470 ;
        RECT 147.430 38.345 152.430 38.705 ;
        RECT 165.385 32.895 166.315 42.825 ;
        RECT 167.045 42.235 168.535 42.615 ;
        RECT 171.885 42.085 172.350 44.975 ;
        RECT 180.320 43.995 181.425 55.870 ;
        RECT 182.175 55.125 182.610 55.510 ;
        RECT 183.105 54.960 183.420 55.870 ;
        RECT 185.650 54.960 185.965 55.870 ;
        RECT 188.210 54.960 188.530 55.870 ;
        RECT 183.105 54.460 188.530 54.960 ;
        RECT 183.105 50.855 183.365 54.460 ;
        RECT 185.690 50.860 185.950 54.460 ;
        RECT 188.270 50.850 188.530 54.460 ;
        RECT 188.995 50.875 194.520 55.870 ;
        RECT 188.995 50.740 194.530 50.875 ;
        RECT 181.820 45.420 182.080 49.075 ;
        RECT 184.400 45.420 184.660 49.075 ;
        RECT 186.980 45.420 187.240 49.075 ;
        RECT 181.820 44.975 187.240 45.420 ;
        RECT 174.230 42.825 182.405 43.995 ;
        RECT 173.200 42.085 173.460 42.095 ;
        RECT 168.040 41.625 176.040 42.085 ;
        RECT 168.040 37.970 168.300 41.625 ;
        RECT 170.620 37.970 170.880 41.625 ;
        RECT 173.200 37.995 173.460 41.625 ;
        RECT 175.780 37.975 176.040 41.625 ;
        RECT 166.750 34.035 167.010 37.690 ;
        RECT 169.330 34.035 169.590 37.690 ;
        RECT 171.910 34.035 172.170 37.690 ;
        RECT 174.490 34.035 174.750 37.690 ;
        RECT 177.070 34.040 177.330 37.690 ;
        RECT 180.220 34.730 181.760 42.825 ;
        RECT 182.555 40.030 183.160 40.455 ;
        RECT 183.490 38.815 183.750 44.975 ;
        RECT 188.995 44.120 190.020 50.740 ;
        RECT 190.785 50.035 191.215 50.415 ;
        RECT 190.430 45.325 190.690 48.980 ;
        RECT 191.720 47.045 191.980 50.740 ;
        RECT 192.980 50.735 194.530 50.740 ;
        RECT 192.995 45.325 193.270 49.045 ;
        RECT 190.430 44.880 193.270 45.325 ;
        RECT 186.125 44.075 190.020 44.120 ;
        RECT 185.570 42.565 190.020 44.075 ;
        RECT 182.200 36.460 182.460 36.895 ;
        RECT 184.780 36.460 185.040 36.895 ;
        RECT 182.200 35.865 185.040 36.460 ;
        RECT 183.355 34.040 183.835 35.865 ;
        RECT 185.570 34.475 186.555 42.565 ;
        RECT 190.930 38.135 191.885 38.580 ;
        RECT 190.700 37.345 190.970 37.735 ;
        RECT 192.995 37.570 193.270 44.880 ;
        RECT 193.750 41.100 194.530 50.735 ;
        RECT 194.935 42.095 195.195 45.735 ;
        RECT 197.515 42.095 197.775 45.730 ;
        RECT 200.100 42.095 200.360 45.740 ;
        RECT 202.690 42.095 202.950 45.725 ;
        RECT 205.250 42.095 205.510 45.725 ;
        RECT 207.825 42.095 208.085 45.730 ;
        RECT 208.525 42.745 209.345 65.560 ;
        RECT 211.070 62.510 211.330 66.200 ;
        RECT 213.645 62.510 213.905 66.200 ;
        RECT 216.240 62.530 216.500 66.200 ;
        RECT 218.795 62.510 219.055 66.200 ;
        RECT 221.370 62.510 221.630 66.200 ;
        RECT 223.315 67.175 230.450 67.495 ;
        RECT 239.905 67.410 240.305 67.450 ;
        RECT 209.750 42.095 210.010 45.720 ;
        RECT 212.345 42.095 212.605 45.720 ;
        RECT 214.935 42.095 215.195 45.720 ;
        RECT 217.485 42.095 217.745 45.745 ;
        RECT 220.100 42.095 220.360 45.720 ;
        RECT 222.670 42.095 222.930 45.720 ;
        RECT 194.935 41.635 222.930 42.095 ;
        RECT 193.750 40.840 195.605 41.100 ;
        RECT 193.750 39.675 195.635 40.840 ;
        RECT 193.750 39.645 195.605 39.675 ;
        RECT 190.700 34.040 190.975 37.345 ;
        RECT 192.995 36.990 193.255 37.570 ;
        RECT 176.630 34.035 192.615 34.040 ;
        RECT 166.745 33.575 192.615 34.035 ;
        RECT 110.475 29.630 118.165 29.635 ;
        RECT 108.730 29.280 118.165 29.630 ;
        RECT 110.475 29.275 118.165 29.280 ;
        RECT 86.265 17.780 89.040 17.785 ;
        RECT 129.505 17.780 130.210 31.165 ;
        RECT 146.965 29.730 147.225 32.510 ;
        RECT 165.385 31.925 179.060 32.895 ;
        RECT 165.720 31.905 179.060 31.925 ;
        RECT 86.265 17.210 130.210 17.780 ;
        RECT 86.310 15.460 89.040 17.210 ;
        RECT 129.505 16.470 130.210 17.210 ;
        RECT 141.165 29.410 147.225 29.730 ;
        RECT 163.475 29.690 174.490 31.005 ;
        RECT 141.165 29.405 145.240 29.410 ;
        RECT 116.850 11.325 117.760 11.375 ;
        RECT 141.165 11.325 142.360 29.405 ;
        RECT 152.310 29.055 167.850 29.415 ;
        RECT 145.475 28.460 160.465 28.515 ;
        RECT 145.475 25.985 161.855 28.460 ;
        RECT 143.205 25.295 143.655 25.345 ;
        RECT 143.205 24.925 147.440 25.295 ;
        RECT 143.205 24.875 143.655 24.925 ;
        RECT 147.915 24.805 148.265 25.985 ;
        RECT 150.450 24.805 150.800 25.985 ;
        RECT 153.015 24.805 153.365 25.985 ;
        RECT 155.620 24.805 155.970 25.985 ;
        RECT 158.205 24.805 158.555 25.985 ;
        RECT 147.915 24.625 158.555 24.805 ;
        RECT 147.915 24.485 158.495 24.625 ;
        RECT 147.915 22.705 148.175 24.485 ;
        RECT 150.495 22.705 150.755 24.485 ;
        RECT 153.075 22.710 153.335 24.485 ;
        RECT 155.655 22.705 155.915 24.485 ;
        RECT 158.235 22.705 158.495 24.485 ;
        RECT 146.625 20.125 146.885 21.925 ;
        RECT 149.205 20.125 149.465 21.925 ;
        RECT 151.785 20.125 152.045 21.925 ;
        RECT 154.365 20.125 154.625 21.925 ;
        RECT 156.945 20.125 157.205 21.925 ;
        RECT 159.525 20.125 159.785 21.920 ;
        RECT 160.265 20.845 161.855 25.985 ;
        RECT 162.375 24.585 162.655 28.685 ;
        RECT 146.625 19.765 167.850 20.125 ;
        RECT 145.480 18.385 159.960 19.290 ;
        RECT 160.575 12.710 161.615 19.765 ;
        RECT 173.615 19.290 174.465 29.690 ;
        RECT 162.425 19.040 174.490 19.290 ;
        RECT 162.425 18.385 174.495 19.040 ;
        RECT 192.150 18.670 192.615 33.575 ;
        RECT 193.750 18.795 194.530 39.645 ;
        RECT 195.255 39.015 195.925 39.415 ;
        RECT 196.235 38.815 196.775 41.635 ;
        RECT 197.515 41.630 197.775 41.635 ;
        RECT 197.105 39.700 198.190 40.840 ;
        RECT 197.310 39.060 197.980 39.460 ;
        RECT 198.795 38.900 199.335 41.635 ;
        RECT 199.680 39.675 200.765 40.815 ;
        RECT 199.905 39.030 200.575 39.430 ;
        RECT 201.400 38.900 201.940 41.635 ;
        RECT 202.690 41.625 202.950 41.635 ;
        RECT 202.340 39.700 203.425 40.840 ;
        RECT 202.515 39.045 203.185 39.445 ;
        RECT 198.765 38.815 199.335 38.900 ;
        RECT 201.385 38.815 201.940 38.900 ;
        RECT 204.040 38.875 204.580 41.635 ;
        RECT 205.250 41.625 205.510 41.635 ;
        RECT 204.785 39.655 205.870 40.795 ;
        RECT 205.095 39.030 205.765 39.430 ;
        RECT 203.980 38.815 204.580 38.875 ;
        RECT 206.505 38.815 207.045 41.635 ;
        RECT 207.825 41.630 208.085 41.635 ;
        RECT 209.750 41.620 210.010 41.635 ;
        RECT 207.400 41.445 207.740 41.485 ;
        RECT 210.130 41.445 210.470 41.480 ;
        RECT 207.395 41.120 210.470 41.445 ;
        RECT 207.490 39.700 210.890 40.730 ;
        RECT 210.295 38.955 210.965 39.355 ;
        RECT 211.430 38.815 211.970 41.635 ;
        RECT 212.345 41.620 212.605 41.635 ;
        RECT 212.490 39.720 213.400 40.795 ;
        RECT 212.485 38.985 213.155 39.385 ;
        RECT 213.950 38.835 214.490 41.635 ;
        RECT 214.935 41.620 215.195 41.635 ;
        RECT 215.000 39.675 215.910 40.750 ;
        RECT 214.960 38.985 215.630 39.385 ;
        RECT 213.930 38.815 214.490 38.835 ;
        RECT 216.575 38.815 217.115 41.635 ;
        RECT 217.680 39.720 218.590 40.795 ;
        RECT 217.660 38.985 218.330 39.385 ;
        RECT 219.095 38.815 219.635 41.635 ;
        RECT 220.100 41.620 220.360 41.635 ;
        RECT 220.125 39.700 221.035 40.775 ;
        RECT 220.195 39.000 220.865 39.400 ;
        RECT 221.395 38.815 221.935 41.635 ;
        RECT 222.670 41.620 222.930 41.635 ;
        RECT 223.315 40.835 224.510 67.175 ;
        RECT 222.290 39.655 224.510 40.835 ;
        RECT 196.235 38.415 221.935 38.815 ;
        RECT 196.235 34.775 196.495 38.415 ;
        RECT 198.765 34.800 199.025 38.415 ;
        RECT 201.385 34.800 201.645 38.415 ;
        RECT 203.980 34.775 204.240 38.415 ;
        RECT 206.555 34.775 206.815 38.415 ;
        RECT 194.945 21.235 195.205 24.975 ;
        RECT 197.490 21.235 197.750 24.980 ;
        RECT 200.090 21.235 200.350 24.970 ;
        RECT 202.680 21.235 202.940 24.970 ;
        RECT 205.240 21.235 205.500 24.970 ;
        RECT 207.820 21.235 208.080 24.970 ;
        RECT 208.575 21.845 209.635 38.090 ;
        RECT 211.350 34.710 211.610 38.415 ;
        RECT 213.930 34.735 214.190 38.415 ;
        RECT 216.480 34.710 216.740 38.415 ;
        RECT 219.080 34.710 219.340 38.415 ;
        RECT 221.675 34.690 221.935 38.415 ;
        RECT 210.065 21.235 210.325 24.915 ;
        RECT 212.635 21.235 212.895 24.905 ;
        RECT 215.235 21.235 215.495 24.905 ;
        RECT 217.795 21.235 218.055 24.895 ;
        RECT 220.375 21.235 220.635 24.895 ;
        RECT 222.955 21.235 223.215 24.905 ;
        RECT 194.945 20.875 223.215 21.235 ;
        RECT 198.835 20.870 200.350 20.875 ;
        RECT 202.680 20.870 202.940 20.875 ;
        RECT 205.240 20.870 205.500 20.875 ;
        RECT 207.820 20.870 208.080 20.875 ;
        RECT 170.300 15.450 174.495 18.385 ;
        RECT 192.125 18.645 193.025 18.670 ;
        RECT 198.835 18.645 200.145 20.870 ;
        RECT 210.065 20.815 210.325 20.875 ;
        RECT 212.635 20.805 212.895 20.875 ;
        RECT 215.235 20.805 215.495 20.875 ;
        RECT 217.795 20.795 218.055 20.875 ;
        RECT 220.375 20.795 220.635 20.875 ;
        RECT 222.955 20.805 223.215 20.875 ;
        RECT 223.630 20.065 224.510 39.655 ;
        RECT 229.570 66.120 230.450 67.175 ;
        RECT 232.865 67.150 242.350 67.410 ;
        RECT 233.515 66.505 233.875 66.615 ;
        RECT 236.845 66.505 237.280 66.520 ;
        RECT 241.385 66.505 241.745 66.615 ;
        RECT 233.425 66.215 241.745 66.505 ;
        RECT 236.845 66.200 237.280 66.215 ;
        RECT 243.635 66.120 244.690 69.055 ;
        RECT 229.570 65.860 231.885 66.120 ;
        RECT 242.330 65.860 244.690 66.120 ;
        RECT 229.570 64.215 230.450 65.860 ;
        RECT 243.635 65.780 244.690 65.860 ;
        RECT 243.635 65.365 246.525 65.780 ;
        RECT 243.680 65.110 246.525 65.365 ;
        RECT 243.680 64.715 246.545 65.110 ;
        RECT 245.470 64.215 246.545 64.715 ;
        RECT 229.570 63.955 231.885 64.215 ;
        RECT 229.570 61.020 230.450 63.955 ;
        RECT 234.165 63.860 234.820 63.980 ;
        RECT 244.330 63.955 246.545 64.215 ;
        RECT 233.505 63.570 241.745 63.860 ;
        RECT 233.515 63.460 233.875 63.570 ;
        RECT 234.165 63.495 234.820 63.570 ;
        RECT 241.385 63.460 241.745 63.570 ;
        RECT 232.865 62.680 233.365 62.925 ;
        RECT 232.860 62.665 233.365 62.680 ;
        RECT 229.570 60.760 231.880 61.020 ;
        RECT 229.570 57.825 230.450 60.760 ;
        RECT 229.570 57.565 231.880 57.825 ;
        RECT 229.570 54.630 230.450 57.565 ;
        RECT 232.860 56.535 233.360 62.665 ;
        RECT 244.330 60.760 244.830 62.925 ;
        RECT 233.500 60.375 241.745 60.665 ;
        RECT 233.510 60.265 233.870 60.375 ;
        RECT 241.385 60.265 241.745 60.375 ;
        RECT 244.330 57.565 244.830 59.730 ;
        RECT 233.510 57.180 241.745 57.470 ;
        RECT 233.510 57.070 233.870 57.180 ;
        RECT 241.385 57.070 241.745 57.180 ;
        RECT 237.700 56.535 238.150 56.625 ;
        RECT 232.860 56.275 242.350 56.535 ;
        RECT 245.470 54.635 246.545 63.955 ;
        RECT 244.760 54.630 246.545 54.635 ;
        RECT 229.570 54.370 231.880 54.630 ;
        RECT 244.330 54.375 246.545 54.630 ;
        RECT 244.330 54.370 244.830 54.375 ;
        RECT 229.570 51.435 230.450 54.370 ;
        RECT 234.185 54.275 234.840 54.355 ;
        RECT 233.510 53.985 241.745 54.275 ;
        RECT 233.510 53.875 233.870 53.985 ;
        RECT 234.185 53.870 234.840 53.985 ;
        RECT 241.385 53.875 241.745 53.985 ;
        RECT 229.570 51.175 231.880 51.435 ;
        RECT 229.570 48.240 230.450 51.175 ;
        RECT 229.570 47.980 231.880 48.240 ;
        RECT 229.570 45.045 230.450 47.980 ;
        RECT 232.860 46.950 233.360 53.340 ;
        RECT 244.330 51.175 244.830 53.340 ;
        RECT 233.510 50.790 241.745 51.080 ;
        RECT 233.510 50.680 233.870 50.790 ;
        RECT 241.385 50.680 241.745 50.790 ;
        RECT 244.330 47.980 244.830 50.145 ;
        RECT 233.510 47.595 241.745 47.885 ;
        RECT 233.510 47.485 233.870 47.595 ;
        RECT 241.385 47.485 241.745 47.595 ;
        RECT 235.910 46.950 236.310 46.990 ;
        RECT 232.860 46.690 242.350 46.950 ;
        RECT 245.470 45.045 246.545 54.375 ;
        RECT 229.570 44.785 231.880 45.045 ;
        RECT 229.570 41.850 230.450 44.785 ;
        RECT 234.150 44.690 234.805 44.820 ;
        RECT 244.330 44.785 246.545 45.045 ;
        RECT 233.510 44.400 241.745 44.690 ;
        RECT 233.510 44.290 233.870 44.400 ;
        RECT 234.150 44.335 234.805 44.400 ;
        RECT 241.385 44.290 241.745 44.400 ;
        RECT 229.570 41.590 231.880 41.850 ;
        RECT 229.570 38.655 230.450 41.590 ;
        RECT 229.570 38.395 231.880 38.655 ;
        RECT 229.570 35.460 230.450 38.395 ;
        RECT 232.860 37.365 233.360 43.755 ;
        RECT 244.330 41.590 244.830 43.755 ;
        RECT 233.510 41.205 241.745 41.495 ;
        RECT 233.510 41.095 233.870 41.205 ;
        RECT 241.385 41.095 241.745 41.205 ;
        RECT 244.330 38.395 244.830 40.560 ;
        RECT 233.510 38.010 241.745 38.300 ;
        RECT 233.510 37.900 233.870 38.010 ;
        RECT 241.385 37.900 241.745 38.010 ;
        RECT 238.530 37.365 238.965 37.405 ;
        RECT 232.860 37.105 242.350 37.365 ;
        RECT 238.530 37.070 238.965 37.105 ;
        RECT 245.470 35.460 246.545 44.785 ;
        RECT 229.570 35.200 231.880 35.460 ;
        RECT 229.570 32.265 230.450 35.200 ;
        RECT 234.200 35.105 234.855 35.230 ;
        RECT 244.330 35.200 246.545 35.460 ;
        RECT 233.510 34.815 241.745 35.105 ;
        RECT 233.510 34.705 233.870 34.815 ;
        RECT 234.200 34.745 234.855 34.815 ;
        RECT 241.385 34.705 241.745 34.815 ;
        RECT 229.570 32.005 231.880 32.265 ;
        RECT 229.570 29.070 230.450 32.005 ;
        RECT 229.570 28.810 231.880 29.070 ;
        RECT 229.570 24.585 230.450 28.810 ;
        RECT 232.860 27.780 233.360 34.170 ;
        RECT 244.330 32.005 244.830 34.170 ;
        RECT 233.510 31.620 241.745 31.910 ;
        RECT 233.510 31.510 233.870 31.620 ;
        RECT 241.385 31.510 241.745 31.620 ;
        RECT 244.330 28.810 244.830 30.975 ;
        RECT 233.515 28.425 241.745 28.715 ;
        RECT 233.515 28.315 233.875 28.425 ;
        RECT 241.385 28.315 241.745 28.425 ;
        RECT 236.850 27.780 237.270 27.825 ;
        RECT 232.860 27.520 242.350 27.780 ;
        RECT 236.850 27.505 237.270 27.520 ;
        RECT 245.470 26.965 246.545 35.200 ;
        RECT 243.565 26.105 246.545 26.965 ;
        RECT 237.690 25.875 238.090 25.915 ;
        RECT 232.860 25.615 242.350 25.875 ;
        RECT 233.510 24.970 233.870 25.080 ;
        RECT 239.395 24.970 239.795 24.980 ;
        RECT 241.385 24.970 241.745 25.080 ;
        RECT 233.510 24.680 241.745 24.970 ;
        RECT 243.590 24.585 244.550 26.105 ;
        RECT 229.570 24.325 231.880 24.585 ;
        RECT 242.330 24.325 244.550 24.585 ;
        RECT 229.570 21.395 230.450 24.325 ;
        RECT 236.005 22.685 236.405 22.720 ;
        RECT 232.860 22.425 242.365 22.685 ;
        RECT 233.510 21.780 233.870 21.890 ;
        RECT 236.165 21.780 236.775 21.785 ;
        RECT 241.400 21.780 241.760 21.890 ;
        RECT 233.510 21.490 241.760 21.780 ;
        RECT 229.570 21.135 231.880 21.395 ;
        RECT 229.570 20.545 230.450 21.135 ;
        RECT 201.195 18.795 224.540 20.065 ;
        RECT 229.570 19.925 234.850 20.545 ;
        RECT 192.125 18.180 200.145 18.645 ;
        RECT 192.125 13.745 193.025 18.180 ;
        RECT 192.105 12.895 193.045 13.745 ;
        RECT 192.125 12.870 193.025 12.895 ;
        RECT 236.165 12.285 236.775 21.490 ;
        RECT 243.590 21.395 244.550 24.325 ;
        RECT 242.345 21.135 244.550 21.395 ;
        RECT 243.590 20.225 244.550 21.135 ;
        RECT 254.575 21.240 254.865 79.930 ;
        RECT 257.440 79.710 259.290 80.220 ;
        RECT 257.440 78.665 257.810 79.710 ;
        RECT 258.920 78.665 259.290 79.710 ;
        RECT 260.400 80.105 273.120 80.220 ;
        RECT 260.400 79.735 273.125 80.105 ;
        RECT 260.400 78.665 260.770 79.735 ;
        RECT 257.440 48.375 257.810 52.795 ;
        RECT 258.920 48.375 259.290 52.795 ;
        RECT 260.400 48.375 260.770 52.795 ;
        RECT 257.440 21.240 257.810 22.505 ;
        RECT 254.575 20.950 257.810 21.240 ;
        RECT 258.920 21.460 259.290 22.505 ;
        RECT 260.400 21.460 260.770 22.505 ;
        RECT 258.920 20.950 260.770 21.460 ;
        RECT 261.180 20.230 261.825 79.395 ;
        RECT 244.785 20.225 261.830 20.230 ;
        RECT 240.505 19.880 261.830 20.225 ;
        RECT 240.500 19.385 261.830 19.880 ;
        RECT 240.500 15.440 243.780 19.385 ;
        RECT 238.745 12.380 239.415 13.145 ;
        RECT 116.850 11.320 142.400 11.325 ;
        RECT 269.530 11.320 270.725 79.735 ;
        RECT 116.850 10.125 270.725 11.320 ;
        RECT 116.850 10.075 117.760 10.125 ;
      LAYER met3 ;
        RECT 59.865 188.815 91.725 216.590 ;
        RECT 94.345 188.815 126.205 216.600 ;
        RECT 59.865 186.200 126.205 188.815 ;
        RECT 59.865 186.190 96.045 186.200 ;
        RECT 89.370 184.310 96.045 186.190 ;
        RECT 59.860 184.300 96.045 184.310 ;
        RECT 59.860 182.230 126.200 184.300 ;
        RECT 55.605 156.685 56.110 157.240 ;
        RECT 16.515 154.485 16.975 156.535 ;
        RECT 59.860 156.135 91.720 182.230 ;
        RECT 34.070 155.765 35.435 156.100 ;
        RECT 11.460 154.025 12.550 154.050 ;
        RECT 9.385 152.935 12.550 154.025 ;
        RECT 11.460 152.910 12.550 152.935 ;
        RECT 16.565 152.545 16.925 154.485 ;
        RECT 31.065 153.845 31.745 153.870 ;
        RECT 34.070 153.845 34.465 155.765 ;
        RECT 53.740 155.720 91.720 156.135 ;
        RECT 59.860 153.910 91.720 155.720 ;
        RECT 94.340 153.900 126.200 182.230 ;
        RECT 31.065 153.460 34.465 153.845 ;
        RECT 31.065 153.435 31.745 153.460 ;
        RECT 16.450 151.980 17.025 152.545 ;
        RECT 11.485 141.520 14.110 141.545 ;
        RECT 9.705 138.895 14.110 141.520 ;
        RECT 11.485 138.870 14.110 138.895 ;
        RECT 16.450 66.250 17.015 151.980 ;
        RECT 55.100 146.940 57.120 146.965 ;
        RECT 55.100 144.920 141.875 146.940 ;
        RECT 55.100 144.895 57.120 144.920 ;
        RECT 103.425 129.640 106.170 130.120 ;
        RECT 26.835 120.325 27.755 120.355 ;
        RECT 26.835 120.320 55.045 120.325 ;
        RECT 26.835 119.970 57.835 120.320 ;
        RECT 26.835 119.965 55.045 119.970 ;
        RECT 26.835 119.345 27.755 119.965 ;
        RECT 103.475 112.875 103.855 129.640 ;
        RECT 125.020 119.995 127.380 120.005 ;
        RECT 136.905 119.995 166.265 135.285 ;
        RECT 125.020 118.695 166.265 119.995 ;
        RECT 125.020 118.660 127.380 118.695 ;
        RECT 82.080 108.945 82.680 109.495 ;
        RECT 136.905 107.385 166.265 118.695 ;
        RECT 127.170 104.465 127.770 105.015 ;
        RECT 162.090 104.355 165.745 107.385 ;
        RECT 57.380 97.655 57.865 98.205 ;
        RECT 73.285 95.155 89.165 95.485 ;
        RECT 125.610 91.915 126.030 94.965 ;
        RECT 131.710 93.380 134.150 93.785 ;
        RECT 131.710 93.375 133.720 93.380 ;
        RECT 131.710 88.220 132.090 93.375 ;
        RECT 136.905 93.060 166.265 104.355 ;
        RECT 134.230 92.560 166.265 93.060 ;
        RECT 58.245 86.915 58.665 87.965 ;
        RECT 83.690 85.035 84.110 88.085 ;
        RECT 134.230 88.010 134.610 92.560 ;
        RECT 83.690 79.895 84.110 82.945 ;
        RECT 136.905 76.455 166.265 92.560 ;
        RECT 219.445 93.015 238.925 93.020 ;
        RECT 219.445 92.675 238.950 93.015 ;
        RECT 219.445 92.670 238.925 92.675 ;
        RECT 219.445 79.615 219.795 92.670 ;
        RECT 182.125 79.265 219.795 79.615 ;
        RECT 224.205 91.890 237.255 92.235 ;
        RECT 224.205 91.210 224.550 91.890 ;
        RECT 236.835 91.210 237.255 91.890 ;
        RECT 237.725 91.480 238.120 92.045 ;
        RECT 44.455 74.480 44.815 74.505 ;
        RECT 40.395 74.120 44.815 74.480 ;
        RECT 44.455 74.095 44.815 74.120 ;
        RECT 125.610 73.590 126.030 76.065 ;
        RECT 136.815 70.020 139.795 72.075 ;
        RECT 16.450 65.685 69.230 66.250 ;
        RECT 37.890 55.810 38.250 55.835 ;
        RECT 36.205 55.450 38.250 55.810 ;
        RECT 37.890 55.425 38.250 55.450 ;
        RECT 68.590 55.480 69.230 65.685 ;
        RECT 167.060 55.510 167.415 59.780 ;
        RECT 70.610 55.480 70.940 55.495 ;
        RECT 68.590 55.180 70.940 55.480 ;
        RECT 70.610 55.165 70.940 55.180 ;
        RECT 167.060 55.165 167.680 55.510 ;
        RECT 182.125 55.485 182.430 79.265 ;
        RECT 190.735 76.550 191.125 76.555 ;
        RECT 224.205 76.550 224.545 91.210 ;
        RECT 234.515 91.120 234.870 91.145 ;
        RECT 228.130 90.755 234.875 91.120 ;
        RECT 237.705 91.105 238.140 91.480 ;
        RECT 237.725 91.095 238.120 91.105 ;
        RECT 234.515 90.730 234.870 90.755 ;
        RECT 236.450 85.335 236.950 85.735 ;
        RECT 229.540 80.275 233.020 82.235 ;
        RECT 190.735 76.210 224.545 76.550 ;
        RECT 182.125 55.150 182.660 55.485 ;
        RECT 39.570 51.670 40.025 53.105 ;
        RECT 39.570 51.175 44.340 51.670 ;
        RECT 39.580 51.170 44.340 51.175 ;
        RECT 40.165 46.945 40.585 48.175 ;
        RECT 43.775 45.165 44.340 51.170 ;
        RECT 53.170 47.945 62.265 48.265 ;
        RECT 47.535 46.245 47.955 46.975 ;
        RECT 47.535 45.745 49.270 46.245 ;
        RECT 30.875 43.650 32.015 44.205 ;
        RECT 40.165 41.035 40.585 41.765 ;
        RECT 47.535 41.740 47.955 42.965 ;
        RECT 48.770 41.035 49.270 45.745 ;
        RECT 53.170 42.840 53.490 47.945 ;
        RECT 61.845 47.215 62.265 47.945 ;
        RECT 54.495 45.835 54.915 46.885 ;
        RECT 53.170 42.520 54.915 42.840 ;
        RECT 40.165 40.535 49.270 41.035 ;
        RECT 36.560 36.930 37.300 37.300 ;
        RECT 40.165 37.280 40.585 40.535 ;
        RECT 47.530 38.715 47.960 39.035 ;
        RECT 40.120 36.950 40.635 37.280 ;
        RECT 47.580 36.615 47.910 38.715 ;
        RECT 54.495 36.750 54.915 42.520 ;
        RECT 61.845 40.410 62.265 41.460 ;
        RECT 61.845 36.755 62.265 37.540 ;
        RECT 51.135 36.615 51.555 36.740 ;
        RECT 35.330 36.270 51.555 36.615 ;
        RECT 35.330 33.720 35.700 36.270 ;
        RECT 54.880 35.850 55.780 36.220 ;
        RECT 59.740 35.860 60.640 36.230 ;
        RECT 59.740 33.725 60.060 35.860 ;
        RECT 52.900 33.720 60.060 33.725 ;
        RECT 35.330 33.405 60.060 33.720 ;
        RECT 35.330 33.350 37.195 33.405 ;
        RECT 35.330 26.000 35.700 33.350 ;
        RECT 50.805 32.735 51.555 33.105 ;
        RECT 52.915 30.140 53.285 33.405 ;
        RECT 36.565 29.770 37.265 30.140 ;
        RECT 51.135 29.770 53.285 30.140 ;
        RECT 50.895 26.190 51.580 26.560 ;
        RECT 35.330 25.630 36.985 26.000 ;
        RECT 38.620 20.945 44.110 23.025 ;
        RECT 19.635 18.705 22.875 18.730 ;
        RECT 19.630 15.455 36.565 18.705 ;
        RECT 73.135 16.750 73.575 51.415 ;
        RECT 78.695 38.985 79.135 51.415 ;
        RECT 190.735 50.390 191.125 76.210 ;
        RECT 236.475 73.490 236.925 85.335 ;
        RECT 238.515 82.140 238.965 82.540 ;
        RECT 237.715 76.185 238.135 76.205 ;
        RECT 237.700 75.750 238.150 76.185 ;
        RECT 237.715 75.730 238.135 75.750 ;
        RECT 235.920 72.965 236.290 72.980 ;
        RECT 235.910 72.555 236.310 72.965 ;
        RECT 235.920 72.540 236.290 72.555 ;
        RECT 195.235 69.055 195.705 70.000 ;
        RECT 195.240 67.170 195.705 69.055 ;
        RECT 195.240 66.825 195.850 67.170 ;
        RECT 234.990 60.715 235.290 60.860 ;
        RECT 234.965 60.325 235.315 60.715 ;
        RECT 234.990 51.130 235.290 60.325 ;
        RECT 234.965 50.740 235.315 51.130 ;
        RECT 190.735 50.060 191.265 50.390 ;
        RECT 126.255 46.395 128.465 46.850 ;
        RECT 162.330 45.535 162.715 47.450 ;
        RECT 162.380 42.590 162.700 45.535 ;
        RECT 126.255 41.955 143.655 42.405 ;
        RECT 78.645 38.505 79.185 38.985 ;
        RECT 78.695 38.475 79.135 38.505 ;
        RECT 115.795 37.710 116.135 38.690 ;
        RECT 128.105 37.710 128.445 41.955 ;
        RECT 143.205 25.320 143.655 41.955 ;
        RECT 162.380 42.260 191.245 42.590 ;
        RECT 162.380 28.660 162.700 42.260 ;
        RECT 182.500 40.430 182.840 42.260 ;
        RECT 182.500 40.280 183.210 40.430 ;
        RECT 182.505 40.055 183.210 40.280 ;
        RECT 190.915 39.365 191.245 42.260 ;
        RECT 195.205 39.365 195.975 39.390 ;
        RECT 197.260 39.365 198.030 39.435 ;
        RECT 199.855 39.365 200.625 39.405 ;
        RECT 202.465 39.365 203.235 39.420 ;
        RECT 205.045 39.365 205.815 39.405 ;
        RECT 220.145 39.365 220.915 39.375 ;
        RECT 190.915 39.035 223.250 39.365 ;
        RECT 190.915 38.555 191.245 39.035 ;
        RECT 210.245 38.980 211.015 39.035 ;
        RECT 212.435 39.010 213.205 39.035 ;
        RECT 214.910 39.010 215.680 39.035 ;
        RECT 217.610 39.010 218.380 39.035 ;
        RECT 220.145 39.025 220.915 39.035 ;
        RECT 190.880 38.160 191.935 38.555 ;
        RECT 137.010 24.900 143.705 25.320 ;
        RECT 39.570 16.310 73.575 16.750 ;
        RECT 19.635 15.430 22.875 15.455 ;
        RECT 39.570 5.235 40.470 16.310 ;
        RECT 86.260 15.550 89.085 16.825 ;
        RECT 137.010 15.590 137.910 24.900 ;
        RECT 162.325 24.610 162.705 28.660 ;
        RECT 234.990 21.830 235.290 50.740 ;
        RECT 235.935 46.640 236.285 72.540 ;
        RECT 236.870 65.890 237.255 66.570 ;
        RECT 237.725 56.225 238.125 75.730 ;
        RECT 238.540 70.295 238.940 82.140 ;
        RECT 239.905 78.945 240.305 79.345 ;
        RECT 238.550 68.915 238.950 69.840 ;
        RECT 239.930 67.100 240.280 78.945 ;
        RECT 239.445 57.520 239.745 60.860 ;
        RECT 239.420 57.130 239.770 57.520 ;
        RECT 237.740 47.935 238.040 47.990 ;
        RECT 237.715 47.545 238.065 47.935 ;
        RECT 236.055 41.545 236.355 41.725 ;
        RECT 236.030 41.155 236.380 41.545 ;
        RECT 236.055 31.960 236.355 41.155 ;
        RECT 236.030 31.570 236.380 31.960 ;
        RECT 236.055 22.770 236.355 31.570 ;
        RECT 237.740 28.765 238.040 47.545 ;
        RECT 239.445 38.350 239.745 57.130 ;
        RECT 239.420 37.960 239.770 38.350 ;
        RECT 238.555 37.020 238.940 37.955 ;
        RECT 237.715 28.375 238.065 28.765 ;
        RECT 236.875 27.455 237.245 28.280 ;
        RECT 237.740 25.965 238.040 28.375 ;
        RECT 237.715 25.565 238.065 25.965 ;
        RECT 239.445 25.030 239.745 37.960 ;
        RECT 239.420 24.630 239.770 25.030 ;
        RECT 236.030 22.375 236.380 22.770 ;
        RECT 234.965 21.440 235.315 21.830 ;
        RECT 170.525 15.740 174.155 18.165 ;
        RECT 240.855 15.780 243.640 18.400 ;
        RECT 97.530 14.690 137.910 15.590 ;
        RECT 39.545 4.345 40.495 5.235 ;
        RECT 39.570 4.340 40.470 4.345 ;
        RECT 97.530 2.065 98.430 14.690 ;
        RECT 160.520 12.730 161.640 13.770 ;
        RECT 116.800 10.100 117.810 11.350 ;
        RECT 116.850 9.695 117.755 10.100 ;
        RECT 116.850 3.380 117.750 9.695 ;
        RECT 116.825 2.490 117.775 3.380 ;
        RECT 192.125 2.830 193.025 13.770 ;
        RECT 236.115 12.310 236.825 13.120 ;
        RECT 238.695 12.405 239.465 13.120 ;
        RECT 116.850 2.485 117.750 2.490 ;
        RECT 97.505 1.175 98.455 2.065 ;
        RECT 192.100 1.940 193.050 2.830 ;
        RECT 192.125 1.935 193.025 1.940 ;
        RECT 97.530 1.170 98.430 1.175 ;
      LAYER met4 ;
        RECT 18.090 224.760 18.095 225.000 ;
        RECT 23.305 224.760 23.310 224.905 ;
        RECT 26.370 224.760 26.375 225.010 ;
        RECT 29.130 224.760 29.140 224.975 ;
        RECT 31.890 224.760 31.895 224.905 ;
        RECT 37.105 224.760 37.110 224.990 ;
        RECT 40.170 224.760 40.175 224.975 ;
        RECT 45.690 224.760 45.695 224.950 ;
        RECT 50.905 224.760 50.910 224.845 ;
        RECT 53.970 224.760 53.975 224.930 ;
        RECT 59.490 224.760 59.495 224.905 ;
        RECT 64.705 224.760 64.710 225.000 ;
        RECT 67.770 224.760 67.775 225.000 ;
        RECT 73.290 224.760 73.295 224.990 ;
        RECT 78.505 224.760 78.510 224.995 ;
        RECT 15.030 220.320 15.330 224.760 ;
        RECT 17.795 220.320 18.095 224.760 ;
        RECT 20.550 220.320 20.850 224.760 ;
        RECT 23.305 220.320 23.605 224.760 ;
        RECT 26.075 220.320 26.375 224.760 ;
        RECT 28.840 220.320 29.140 224.760 ;
        RECT 31.595 220.320 31.895 224.760 ;
        RECT 34.350 220.320 34.650 224.760 ;
        RECT 37.105 220.320 37.405 224.760 ;
        RECT 39.875 220.320 40.175 224.760 ;
        RECT 42.630 220.320 42.930 224.760 ;
        RECT 45.395 220.320 45.695 224.760 ;
        RECT 48.150 220.320 48.450 224.760 ;
        RECT 50.905 220.320 51.205 224.760 ;
        RECT 53.675 220.320 53.975 224.760 ;
        RECT 56.430 220.320 56.730 224.760 ;
        RECT 59.195 220.320 59.495 224.760 ;
        RECT 61.950 220.320 62.250 224.760 ;
        RECT 64.705 220.320 65.005 224.760 ;
        RECT 67.475 220.320 67.775 224.760 ;
        RECT 70.230 220.320 70.530 224.760 ;
        RECT 72.995 220.320 73.295 224.760 ;
        RECT 75.750 220.320 76.050 224.760 ;
        RECT 78.505 222.640 78.810 224.760 ;
        RECT 78.505 220.320 78.805 222.640 ;
        RECT 6.000 218.605 79.635 220.320 ;
        RECT 60.260 186.585 89.870 216.195 ;
        RECT 85.155 183.915 88.470 186.585 ;
        RECT 91.225 186.250 91.705 216.530 ;
        RECT 94.740 186.595 124.350 216.205 ;
        RECT 60.255 157.215 89.865 183.915 ;
        RECT 55.650 156.705 89.865 157.215 ;
        RECT 9.410 154.025 10.500 154.030 ;
        RECT 6.000 152.935 10.500 154.025 ;
        RECT 9.410 152.930 10.500 152.935 ;
        RECT 57.985 151.930 58.775 156.705 ;
        RECT 60.255 154.305 89.865 156.705 ;
        RECT 31.075 150.660 58.775 151.930 ;
        RECT 86.685 152.180 89.830 154.305 ;
        RECT 91.220 153.970 91.700 184.250 ;
        RECT 96.770 183.905 99.940 186.595 ;
        RECT 125.705 186.260 126.185 216.540 ;
        RECT 94.735 154.295 124.345 183.905 ;
        RECT 94.785 152.180 97.995 154.295 ;
        RECT 125.700 153.960 126.180 184.240 ;
        RECT 9.730 141.520 12.355 141.525 ;
        RECT 6.000 138.895 12.355 141.520 ;
        RECT 9.730 138.890 12.355 138.895 ;
        RECT 31.075 74.480 32.345 150.660 ;
        RECT 86.685 149.030 97.995 152.180 ;
        RECT 139.830 146.940 141.850 146.945 ;
        RECT 139.830 144.920 173.540 146.940 ;
        RECT 139.830 144.915 141.850 144.920 ;
        RECT 82.125 108.965 82.635 109.475 ;
        RECT 57.425 98.180 57.820 98.185 ;
        RECT 56.625 97.680 57.865 98.180 ;
        RECT 56.625 87.945 57.125 97.680 ;
        RECT 57.425 97.675 57.820 97.680 ;
        RECT 56.625 87.445 58.620 87.945 ;
        RECT 58.290 86.935 58.620 87.445 ;
        RECT 82.130 85.555 82.630 108.965 ;
        RECT 136.925 107.445 137.405 135.225 ;
        RECT 138.760 107.780 165.870 134.890 ;
        RECT 138.760 106.010 141.865 107.780 ;
        RECT 133.595 105.500 141.865 106.010 ;
        RECT 127.215 104.485 127.725 104.995 ;
        RECT 125.655 92.435 125.985 94.945 ;
        RECT 127.220 92.435 127.720 104.485 ;
        RECT 133.595 93.400 134.105 105.500 ;
        RECT 125.655 91.935 127.720 92.435 ;
        RECT 83.735 85.555 84.065 88.065 ;
        RECT 82.130 85.055 84.065 85.555 ;
        RECT 82.130 76.045 82.630 85.055 ;
        RECT 127.220 82.925 127.720 91.935 ;
        RECT 83.735 82.425 127.720 82.925 ;
        RECT 83.735 79.915 84.065 82.425 ;
        RECT 136.925 76.515 137.405 104.295 ;
        RECT 138.760 103.960 141.865 105.500 ;
        RECT 138.760 76.850 165.870 103.960 ;
        RECT 171.520 100.060 173.540 144.920 ;
        RECT 171.520 98.685 315.000 100.060 ;
        RECT 171.595 98.060 315.000 98.685 ;
        RECT 82.130 75.545 125.985 76.045 ;
        RECT 40.420 74.480 40.780 74.485 ;
        RECT 31.075 74.120 40.780 74.480 ;
        RECT 31.075 55.810 32.345 74.120 ;
        RECT 40.420 74.115 40.780 74.120 ;
        RECT 125.655 73.655 125.985 75.545 ;
        RECT 136.860 72.040 139.750 72.055 ;
        RECT 171.595 72.040 173.595 98.060 ;
        RECT 228.155 91.120 228.520 91.125 ;
        RECT 222.600 90.755 228.520 91.120 ;
        RECT 222.600 77.965 222.965 90.755 ;
        RECT 228.155 90.750 228.520 90.755 ;
        RECT 229.595 82.215 232.975 98.060 ;
        RECT 234.510 90.755 236.285 91.120 ;
        RECT 229.585 80.295 232.975 82.215 ;
        RECT 136.860 70.040 173.595 72.040 ;
        RECT 176.940 77.600 222.965 77.965 ;
        RECT 229.595 77.770 232.975 80.295 ;
        RECT 176.940 61.720 177.305 77.600 ;
        RECT 235.920 73.465 236.285 90.755 ;
        RECT 235.915 72.585 236.295 73.465 ;
        RECT 236.890 66.525 237.230 91.550 ;
        RECT 237.730 76.590 238.115 91.485 ;
        RECT 237.710 75.775 238.140 76.590 ;
        RECT 238.575 69.795 238.925 93.020 ;
        RECT 238.570 69.375 238.930 69.795 ;
        RECT 236.890 66.195 237.235 66.525 ;
        RECT 236.890 65.845 237.230 66.195 ;
        RECT 167.060 61.355 177.305 61.720 ;
        RECT 167.060 59.755 167.415 61.355 ;
        RECT 167.055 59.400 167.420 59.755 ;
        RECT 36.230 55.810 36.590 55.815 ;
        RECT 31.075 55.450 36.590 55.810 ;
        RECT 36.230 55.445 36.590 55.450 ;
        RECT 40.210 47.755 49.785 48.155 ;
        RECT 40.210 46.970 40.540 47.755 ;
        RECT 30.920 43.670 31.970 44.185 ;
        RECT 6.000 15.455 27.270 18.705 ;
        RECT 30.925 13.770 31.965 43.670 ;
        RECT 49.285 42.945 49.785 47.755 ;
        RECT 54.540 46.175 54.870 46.865 ;
        RECT 115.800 46.805 128.430 46.810 ;
        RECT 115.800 46.440 128.445 46.805 ;
        RECT 115.800 46.430 128.430 46.440 ;
        RECT 54.540 45.855 63.640 46.175 ;
        RECT 47.580 42.445 49.785 42.945 ;
        RECT 47.580 39.040 47.910 42.445 ;
        RECT 61.890 40.750 62.220 41.440 ;
        RECT 63.320 40.750 63.640 45.855 ;
        RECT 61.890 40.430 63.640 40.750 ;
        RECT 47.575 38.710 47.915 39.040 ;
        RECT 61.890 38.985 62.220 40.430 ;
        RECT 78.690 38.985 79.140 38.990 ;
        RECT 61.890 38.510 79.250 38.985 ;
        RECT 40.165 37.280 40.590 37.285 ;
        RECT 36.610 36.950 52.740 37.280 ;
        RECT 40.165 36.945 40.590 36.950 ;
        RECT 52.410 33.085 52.740 36.950 ;
        RECT 61.890 36.775 62.220 38.510 ;
        RECT 63.705 38.505 79.250 38.510 ;
        RECT 78.690 38.500 79.140 38.505 ;
        RECT 115.800 37.755 116.130 46.430 ;
        RECT 34.850 32.755 52.740 33.085 ;
        RECT 34.850 30.120 35.180 32.755 ;
        RECT 34.850 29.790 36.940 30.120 ;
        RECT 52.410 29.660 52.740 32.755 ;
        RECT 54.925 35.870 55.735 36.200 ;
        RECT 54.925 29.660 55.245 35.870 ;
        RECT 52.410 29.340 55.245 29.660 ;
        RECT 52.410 26.540 52.740 29.340 ;
        RECT 236.895 27.500 237.230 65.845 ;
        RECT 238.575 37.065 238.925 69.375 ;
        RECT 51.175 26.210 52.740 26.540 ;
        RECT 38.670 23.005 44.060 24.080 ;
        RECT 38.665 20.965 44.065 23.005 ;
        RECT 33.290 18.705 36.540 18.710 ;
        RECT 38.670 18.705 44.060 20.965 ;
        RECT 33.290 15.455 243.830 18.705 ;
        RECT 33.290 15.450 36.540 15.455 ;
        RECT 160.545 13.770 161.585 13.775 ;
        RECT 30.925 12.730 161.585 13.770 ;
        RECT 160.545 12.725 161.585 12.730 ;
        RECT 236.160 12.330 236.780 13.100 ;
        RECT 238.740 12.425 239.420 13.100 ;
        RECT 236.165 8.070 236.775 12.330 ;
        RECT 58.890 7.170 236.775 8.070 ;
        RECT 39.570 1.000 40.470 5.240 ;
        RECT 58.890 1.000 59.790 7.170 ;
        RECT 238.745 5.305 239.415 12.425 ;
        RECT 78.210 4.405 239.420 5.305 ;
        RECT 78.210 1.000 79.110 4.405 ;
        RECT 238.745 4.400 239.415 4.405 ;
        RECT 97.530 1.375 98.430 2.070 ;
        RECT 97.525 1.000 98.430 1.375 ;
        RECT 116.850 1.000 117.750 3.385 ;
        RECT 136.170 1.935 193.025 2.835 ;
        RECT 136.170 1.315 137.070 1.935 ;
        RECT 136.165 1.000 137.070 1.315 ;
  END
END tt_um_DalinEM_asic_1
END LIBRARY

