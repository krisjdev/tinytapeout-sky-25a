VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_cw_vref
  CLASS BLOCK ;
  FOREIGN tt_um_cw_vref ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 320.000000 ;
    ANTENNADIFFAREA 9.280000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 1032.322510 ;
    ANTENNADIFFAREA 940.731567 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1728.040771 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    USE POWER ;
    ANTENNAGATEAREA 1032.322510 ;
    ANTENNADIFFAREA 940.731567 ;
    PORT
      LAYER met4 ;
        RECT 177.615 2.590 179.215 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.615 2.590 219.215 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.600 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 180.915 2.590 182.515 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 220.915 2.590 222.515 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.600 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    USE POWER ;
    ANTENNAGATEAREA 2912.000000 ;
    ANTENNADIFFAREA 2005.394531 ;
    PORT
      LAYER met4 ;
        RECT 6.200 5.000 7.800 220.760 ;
    END
  END VAPWR
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  OBS
      LAYER nwell ;
        RECT 3.250 220.980 103.675 223.480 ;
        RECT 3.250 5.750 5.750 220.980 ;
        RECT 8.935 180.290 45.725 212.250 ;
        RECT 48.860 187.290 56.700 210.740 ;
      LAYER pwell ;
        RECT 9.140 168.330 52.250 178.810 ;
      LAYER nwell ;
        RECT 62.865 170.855 99.075 217.105 ;
        RECT 101.175 182.070 103.675 220.980 ;
        RECT 108.240 216.015 153.520 220.985 ;
        RECT 108.240 203.045 153.520 214.015 ;
      LAYER pwell ;
        RECT 108.440 184.690 153.320 201.100 ;
      LAYER nwell ;
        RECT 161.905 200.075 236.345 201.680 ;
      LAYER pwell ;
        RECT 162.100 198.875 163.470 199.685 ;
        RECT 165.780 199.555 167.125 199.785 ;
        RECT 163.480 198.875 165.310 199.555 ;
        RECT 165.780 198.875 167.610 199.555 ;
        RECT 167.620 198.875 173.130 199.685 ;
        RECT 173.140 198.875 174.970 199.685 ;
        RECT 174.990 198.960 175.420 199.745 ;
        RECT 175.925 199.555 177.270 199.785 ;
        RECT 175.440 198.875 177.270 199.555 ;
        RECT 177.280 198.875 182.790 199.685 ;
        RECT 182.800 198.875 184.630 199.685 ;
        RECT 185.585 199.555 186.930 199.785 ;
        RECT 185.100 198.875 186.930 199.555 ;
        RECT 187.870 198.960 188.300 199.745 ;
        RECT 188.320 198.875 193.830 199.685 ;
        RECT 195.245 199.555 196.590 199.785 ;
        RECT 194.760 198.875 196.590 199.555 ;
        RECT 196.600 198.875 200.270 199.685 ;
        RECT 200.750 198.960 201.180 199.745 ;
        RECT 201.200 198.875 203.950 199.685 ;
        RECT 204.905 199.555 206.250 199.785 ;
        RECT 204.420 198.875 206.250 199.555 ;
        RECT 206.260 198.875 211.770 199.685 ;
        RECT 211.780 198.875 213.610 199.685 ;
        RECT 213.630 198.960 214.060 199.745 ;
        RECT 214.565 199.555 215.910 199.785 ;
        RECT 214.080 198.875 215.910 199.555 ;
        RECT 215.920 198.875 221.430 199.685 ;
        RECT 221.440 198.875 223.270 199.685 ;
        RECT 224.225 199.555 225.570 199.785 ;
        RECT 223.740 198.875 225.570 199.555 ;
        RECT 226.510 198.960 226.940 199.745 ;
        RECT 226.960 198.875 232.470 199.685 ;
        RECT 233.425 199.555 234.770 199.785 ;
        RECT 232.940 198.875 234.770 199.555 ;
        RECT 234.780 198.875 236.150 199.685 ;
        RECT 162.240 198.665 162.410 198.875 ;
        RECT 163.620 198.665 163.790 198.875 ;
        RECT 165.455 198.715 165.575 198.825 ;
        RECT 167.300 198.685 167.470 198.875 ;
        RECT 167.760 198.685 167.930 198.875 ;
        RECT 169.140 198.665 169.310 198.855 ;
        RECT 173.280 198.685 173.450 198.875 ;
        RECT 174.660 198.665 174.830 198.855 ;
        RECT 175.580 198.685 175.750 198.875 ;
        RECT 177.420 198.685 177.590 198.875 ;
        RECT 180.180 198.665 180.350 198.855 ;
        RECT 182.940 198.685 183.110 198.875 ;
        RECT 184.775 198.715 184.895 198.825 ;
        RECT 185.240 198.685 185.410 198.875 ;
        RECT 185.700 198.665 185.870 198.855 ;
        RECT 187.090 198.720 187.250 198.830 ;
        RECT 187.535 198.715 187.655 198.825 ;
        RECT 188.460 198.665 188.630 198.875 ;
        RECT 193.980 198.665 194.150 198.855 ;
        RECT 194.900 198.685 195.070 198.875 ;
        RECT 196.740 198.685 196.910 198.875 ;
        RECT 199.500 198.665 199.670 198.855 ;
        RECT 200.415 198.715 200.535 198.825 ;
        RECT 201.340 198.685 201.510 198.875 ;
        RECT 204.095 198.715 204.215 198.825 ;
        RECT 204.560 198.685 204.730 198.875 ;
        RECT 205.020 198.665 205.190 198.855 ;
        RECT 206.400 198.685 206.570 198.875 ;
        RECT 210.540 198.665 210.710 198.855 ;
        RECT 211.920 198.685 212.090 198.875 ;
        RECT 213.295 198.715 213.415 198.825 ;
        RECT 214.220 198.665 214.390 198.875 ;
        RECT 216.060 198.685 216.230 198.875 ;
        RECT 219.740 198.665 219.910 198.855 ;
        RECT 221.580 198.685 221.750 198.875 ;
        RECT 223.415 198.715 223.535 198.825 ;
        RECT 223.880 198.685 224.050 198.875 ;
        RECT 225.260 198.665 225.430 198.855 ;
        RECT 225.730 198.720 225.890 198.830 ;
        RECT 227.100 198.685 227.270 198.875 ;
        RECT 230.780 198.665 230.950 198.855 ;
        RECT 232.615 198.715 232.735 198.825 ;
        RECT 233.080 198.685 233.250 198.875 ;
        RECT 234.455 198.715 234.575 198.825 ;
        RECT 235.840 198.665 236.010 198.875 ;
        RECT 162.100 197.855 163.470 198.665 ;
        RECT 163.480 197.855 168.990 198.665 ;
        RECT 169.000 197.855 174.510 198.665 ;
        RECT 174.520 197.855 180.030 198.665 ;
        RECT 180.040 197.855 185.550 198.665 ;
        RECT 185.560 197.855 187.390 198.665 ;
        RECT 187.870 197.795 188.300 198.580 ;
        RECT 188.320 197.855 193.830 198.665 ;
        RECT 193.840 197.855 199.350 198.665 ;
        RECT 199.360 197.855 204.870 198.665 ;
        RECT 204.880 197.855 210.390 198.665 ;
        RECT 210.400 197.855 213.150 198.665 ;
        RECT 213.630 197.795 214.060 198.580 ;
        RECT 214.080 197.855 219.590 198.665 ;
        RECT 219.600 197.855 225.110 198.665 ;
        RECT 225.120 197.855 230.630 198.665 ;
        RECT 230.640 197.855 234.310 198.665 ;
        RECT 234.780 197.855 236.150 198.665 ;
      LAYER nwell ;
        RECT 161.905 194.635 236.345 197.465 ;
      LAYER pwell ;
        RECT 162.100 193.435 163.470 194.245 ;
        RECT 163.480 193.435 168.990 194.245 ;
        RECT 169.000 193.435 174.510 194.245 ;
        RECT 174.990 193.520 175.420 194.305 ;
        RECT 175.450 193.435 176.800 194.345 ;
        RECT 176.820 193.435 182.330 194.245 ;
        RECT 182.340 193.435 187.850 194.245 ;
        RECT 187.860 193.435 193.370 194.245 ;
        RECT 193.380 193.435 198.890 194.245 ;
        RECT 198.900 193.435 200.730 194.245 ;
        RECT 200.750 193.520 201.180 194.305 ;
        RECT 201.200 193.435 206.710 194.245 ;
        RECT 206.720 193.435 212.230 194.245 ;
        RECT 212.240 193.435 217.750 194.245 ;
        RECT 217.760 193.435 223.270 194.245 ;
        RECT 223.280 193.435 226.030 194.245 ;
        RECT 226.510 193.520 226.940 194.305 ;
        RECT 226.960 193.435 232.470 194.245 ;
        RECT 232.480 193.435 234.310 194.245 ;
        RECT 234.780 193.435 236.150 194.245 ;
        RECT 162.240 193.225 162.410 193.435 ;
        RECT 163.620 193.225 163.790 193.435 ;
        RECT 169.140 193.245 169.310 193.435 ;
        RECT 170.980 193.225 171.150 193.415 ;
        RECT 172.820 193.225 172.990 193.415 ;
        RECT 174.660 193.385 174.830 193.415 ;
        RECT 174.655 193.275 174.830 193.385 ;
        RECT 174.660 193.225 174.830 193.275 ;
        RECT 175.120 193.225 175.290 193.415 ;
        RECT 176.500 193.245 176.670 193.435 ;
        RECT 176.960 193.245 177.130 193.435 ;
        RECT 177.880 193.225 178.050 193.415 ;
        RECT 180.640 193.225 180.810 193.415 ;
        RECT 181.100 193.225 181.270 193.415 ;
        RECT 182.480 193.245 182.650 193.435 ;
        RECT 184.780 193.225 184.950 193.415 ;
        RECT 187.535 193.275 187.655 193.385 ;
        RECT 188.000 193.245 188.170 193.435 ;
        RECT 188.460 193.225 188.630 193.415 ;
        RECT 193.520 193.245 193.690 193.435 ;
        RECT 193.975 193.275 194.095 193.385 ;
        RECT 194.440 193.225 194.610 193.415 ;
        RECT 197.200 193.225 197.370 193.415 ;
        RECT 199.040 193.245 199.210 193.435 ;
        RECT 200.880 193.225 201.050 193.415 ;
        RECT 201.340 193.245 201.510 193.435 ;
        RECT 204.560 193.225 204.730 193.415 ;
        RECT 205.020 193.225 205.190 193.415 ;
        RECT 206.860 193.245 207.030 193.435 ;
        RECT 210.540 193.225 210.710 193.415 ;
        RECT 212.380 193.245 212.550 193.435 ;
        RECT 213.295 193.275 213.415 193.385 ;
        RECT 214.220 193.225 214.390 193.415 ;
        RECT 217.900 193.245 218.070 193.435 ;
        RECT 219.740 193.225 219.910 193.415 ;
        RECT 223.420 193.245 223.590 193.435 ;
        RECT 225.260 193.225 225.430 193.415 ;
        RECT 226.175 193.275 226.295 193.385 ;
        RECT 227.100 193.245 227.270 193.435 ;
        RECT 230.780 193.225 230.950 193.415 ;
        RECT 232.620 193.245 232.790 193.435 ;
        RECT 234.455 193.275 234.575 193.385 ;
        RECT 235.840 193.225 236.010 193.435 ;
        RECT 162.100 192.415 163.470 193.225 ;
        RECT 163.480 192.415 168.990 193.225 ;
        RECT 169.920 192.445 171.290 193.225 ;
        RECT 171.300 192.545 173.130 193.225 ;
        RECT 173.140 192.545 174.970 193.225 ;
        RECT 174.980 192.545 177.720 193.225 ;
        RECT 177.740 192.545 179.570 193.225 ;
        RECT 173.140 192.315 174.485 192.545 ;
        RECT 178.225 192.315 179.570 192.545 ;
        RECT 179.580 192.445 180.950 193.225 ;
        RECT 180.960 192.415 184.630 193.225 ;
        RECT 184.640 192.315 187.390 193.225 ;
        RECT 187.870 192.355 188.300 193.140 ;
        RECT 188.320 192.415 193.830 193.225 ;
        RECT 194.300 192.315 197.050 193.225 ;
        RECT 197.060 192.415 200.730 193.225 ;
        RECT 200.740 192.415 202.110 193.225 ;
        RECT 202.120 192.315 204.870 193.225 ;
        RECT 204.880 192.415 210.390 193.225 ;
        RECT 210.400 192.415 213.150 193.225 ;
        RECT 213.630 192.355 214.060 193.140 ;
        RECT 214.080 192.415 219.590 193.225 ;
        RECT 219.600 192.415 225.110 193.225 ;
        RECT 225.120 192.415 230.630 193.225 ;
        RECT 230.640 192.415 234.310 193.225 ;
        RECT 234.780 192.415 236.150 193.225 ;
      LAYER nwell ;
        RECT 161.905 189.195 236.345 192.025 ;
      LAYER pwell ;
        RECT 162.100 187.995 163.470 188.805 ;
        RECT 163.480 187.995 164.850 188.775 ;
        RECT 164.860 187.995 166.690 188.805 ;
        RECT 166.700 187.995 168.070 188.775 ;
        RECT 168.080 187.995 169.450 188.775 ;
        RECT 169.460 187.995 171.290 188.675 ;
        RECT 171.440 187.995 174.890 188.905 ;
        RECT 174.990 188.080 175.420 188.865 ;
        RECT 175.580 187.995 179.030 188.905 ;
        RECT 179.580 187.995 183.235 188.905 ;
        RECT 183.260 188.225 185.095 188.905 ;
        RECT 183.405 187.995 185.095 188.225 ;
        RECT 186.020 187.995 189.675 188.905 ;
        RECT 190.160 188.225 191.995 188.905 ;
        RECT 190.305 187.995 191.995 188.225 ;
        RECT 192.460 187.995 195.210 188.805 ;
        RECT 195.680 188.675 196.610 188.905 ;
        RECT 195.680 187.995 199.580 188.675 ;
        RECT 200.750 188.080 201.180 188.865 ;
        RECT 201.200 187.995 206.710 188.805 ;
        RECT 206.720 187.995 210.390 188.805 ;
        RECT 211.320 187.995 214.070 188.905 ;
        RECT 214.080 187.995 219.590 188.805 ;
        RECT 219.600 187.995 222.350 188.805 ;
        RECT 222.820 187.995 225.570 188.905 ;
        RECT 226.510 188.080 226.940 188.865 ;
        RECT 226.960 187.995 228.330 188.775 ;
        RECT 228.340 187.995 229.710 188.775 ;
        RECT 229.720 187.995 231.090 188.775 ;
        RECT 231.100 187.995 234.770 188.805 ;
        RECT 234.780 187.995 236.150 188.805 ;
        RECT 162.240 187.785 162.410 187.995 ;
        RECT 163.620 187.785 163.790 187.995 ;
        RECT 165.000 187.785 165.170 187.995 ;
        RECT 166.380 187.785 166.550 187.975 ;
        RECT 166.840 187.805 167.010 187.995 ;
        RECT 167.760 187.785 167.930 187.975 ;
        RECT 168.220 187.805 168.390 187.995 ;
        RECT 170.980 187.805 171.150 187.995 ;
        RECT 173.740 187.785 173.910 187.975 ;
        RECT 174.210 187.830 174.370 187.940 ;
        RECT 174.660 187.805 174.830 187.995 ;
        RECT 178.800 187.975 178.970 187.995 ;
        RECT 175.120 187.785 175.290 187.975 ;
        RECT 177.890 187.830 178.050 187.940 ;
        RECT 178.800 187.805 178.975 187.975 ;
        RECT 179.255 187.835 179.375 187.945 ;
        RECT 179.725 187.805 179.895 187.995 ;
        RECT 178.805 187.785 178.975 187.805 ;
        RECT 181.100 187.785 181.270 187.975 ;
        RECT 182.480 187.785 182.650 187.975 ;
        RECT 183.405 187.805 183.575 187.995 ;
        RECT 183.860 187.785 184.030 187.975 ;
        RECT 185.695 187.940 185.815 187.945 ;
        RECT 185.695 187.835 185.870 187.940 ;
        RECT 185.710 187.830 185.870 187.835 ;
        RECT 186.165 187.805 186.335 187.995 ;
        RECT 186.620 187.785 186.790 187.975 ;
        RECT 188.455 187.835 188.575 187.945 ;
        RECT 188.920 187.785 189.090 187.975 ;
        RECT 189.835 187.835 189.955 187.945 ;
        RECT 190.305 187.785 190.475 187.995 ;
        RECT 192.600 187.805 192.770 187.995 ;
        RECT 194.900 187.785 195.070 187.975 ;
        RECT 195.365 187.945 195.535 187.975 ;
        RECT 195.355 187.835 195.535 187.945 ;
        RECT 195.365 187.785 195.535 187.835 ;
        RECT 196.095 187.805 196.265 187.995 ;
        RECT 199.960 187.785 200.130 187.975 ;
        RECT 200.420 187.785 200.590 187.975 ;
        RECT 201.340 187.805 201.510 187.995 ;
        RECT 205.940 187.785 206.110 187.975 ;
        RECT 206.860 187.805 207.030 187.995 ;
        RECT 208.240 187.785 208.410 187.975 ;
        RECT 209.620 187.785 209.790 187.975 ;
        RECT 210.080 187.785 210.250 187.975 ;
        RECT 210.550 187.840 210.710 187.950 ;
        RECT 211.460 187.785 211.630 187.975 ;
        RECT 212.850 187.830 213.010 187.940 ;
        RECT 213.760 187.805 213.930 187.995 ;
        RECT 214.220 187.785 214.390 187.995 ;
        RECT 215.600 187.785 215.770 187.975 ;
        RECT 217.900 187.785 218.070 187.975 ;
        RECT 219.280 187.785 219.450 187.975 ;
        RECT 219.740 187.945 219.910 187.995 ;
        RECT 219.735 187.835 219.910 187.945 ;
        RECT 219.740 187.805 219.910 187.835 ;
        RECT 220.200 187.785 220.370 187.975 ;
        RECT 222.495 187.835 222.615 187.945 ;
        RECT 222.960 187.805 223.130 187.995 ;
        RECT 225.730 187.840 225.890 187.950 ;
        RECT 227.100 187.805 227.270 187.995 ;
        RECT 229.400 187.805 229.570 187.995 ;
        RECT 230.780 187.805 230.950 187.995 ;
        RECT 231.240 187.805 231.410 187.995 ;
        RECT 232.160 187.785 232.330 187.975 ;
        RECT 233.540 187.785 233.710 187.975 ;
        RECT 234.010 187.830 234.170 187.940 ;
        RECT 235.840 187.785 236.010 187.995 ;
        RECT 162.100 186.975 163.470 187.785 ;
        RECT 163.480 187.005 164.850 187.785 ;
        RECT 164.860 187.005 166.230 187.785 ;
        RECT 166.240 187.005 167.610 187.785 ;
        RECT 167.620 186.875 170.370 187.785 ;
        RECT 170.520 186.875 173.970 187.785 ;
        RECT 174.980 186.875 177.730 187.785 ;
        RECT 178.805 187.555 180.495 187.785 ;
        RECT 178.660 186.875 180.495 187.555 ;
        RECT 180.960 187.005 182.330 187.785 ;
        RECT 182.340 187.005 183.710 187.785 ;
        RECT 183.720 187.105 185.550 187.785 ;
        RECT 184.205 186.875 185.550 187.105 ;
        RECT 186.480 187.005 187.850 187.785 ;
        RECT 187.870 186.915 188.300 187.700 ;
        RECT 188.780 187.005 190.150 187.785 ;
        RECT 190.160 186.875 193.815 187.785 ;
        RECT 193.840 187.005 195.210 187.785 ;
        RECT 195.220 186.875 198.875 187.785 ;
        RECT 198.900 187.005 200.270 187.785 ;
        RECT 200.280 186.975 205.790 187.785 ;
        RECT 205.800 186.975 207.170 187.785 ;
        RECT 207.180 187.005 208.550 187.785 ;
        RECT 208.560 187.005 209.930 187.785 ;
        RECT 209.940 187.005 211.310 187.785 ;
        RECT 211.320 187.005 212.690 187.785 ;
        RECT 213.630 186.915 214.060 187.700 ;
        RECT 214.080 187.005 215.450 187.785 ;
        RECT 215.460 187.005 216.830 187.785 ;
        RECT 216.840 187.005 218.210 187.785 ;
        RECT 218.220 187.005 219.590 187.785 ;
        RECT 220.060 187.615 221.820 187.785 ;
        RECT 220.060 187.570 222.315 187.615 ;
        RECT 220.060 187.535 223.255 187.570 ;
        RECT 224.615 187.535 229.710 187.785 ;
        RECT 220.060 187.105 229.710 187.535 ;
        RECT 221.385 186.935 224.615 187.105 ;
        RECT 222.325 186.890 224.615 186.935 ;
        RECT 223.265 186.855 224.615 186.890 ;
        RECT 227.690 186.875 229.710 187.105 ;
        RECT 229.720 186.875 232.470 187.785 ;
        RECT 232.480 187.005 233.850 187.785 ;
        RECT 234.780 186.975 236.150 187.785 ;
        RECT 227.690 186.855 228.610 186.875 ;
      LAYER nwell ;
        RECT 161.905 183.755 236.345 186.585 ;
      LAYER pwell ;
        RECT 162.100 182.555 163.470 183.365 ;
        RECT 163.940 182.555 165.310 183.335 ;
        RECT 165.320 182.555 166.690 183.335 ;
        RECT 166.715 182.555 170.370 183.465 ;
        RECT 171.300 182.555 174.955 183.465 ;
        RECT 174.990 182.640 175.420 183.425 ;
        RECT 175.580 182.555 179.030 183.465 ;
        RECT 179.580 182.555 180.950 183.335 ;
        RECT 180.960 182.555 182.330 183.335 ;
        RECT 182.340 182.555 183.710 183.335 ;
        RECT 183.720 182.555 185.090 183.335 ;
        RECT 185.100 182.555 186.470 183.335 ;
        RECT 186.480 182.785 188.315 183.465 ;
        RECT 186.625 182.555 188.315 182.785 ;
        RECT 188.780 182.555 192.435 183.465 ;
        RECT 192.460 182.555 196.115 183.465 ;
        RECT 196.140 183.235 197.070 183.465 ;
        RECT 208.545 183.450 209.895 183.485 ;
        RECT 196.140 182.555 200.040 183.235 ;
        RECT 200.750 182.640 201.180 183.425 ;
        RECT 207.605 183.405 209.895 183.450 ;
        RECT 201.200 182.555 202.570 183.335 ;
        RECT 202.580 182.555 203.950 183.335 ;
        RECT 203.960 182.555 205.330 183.365 ;
        RECT 206.665 183.235 209.895 183.405 ;
        RECT 212.970 183.465 213.890 183.485 ;
        RECT 212.970 183.235 214.990 183.465 ;
        RECT 220.045 183.450 221.395 183.485 ;
        RECT 219.105 183.405 221.395 183.450 ;
        RECT 205.340 182.805 214.990 183.235 ;
        RECT 205.340 182.770 208.535 182.805 ;
        RECT 205.340 182.725 207.595 182.770 ;
        RECT 205.340 182.555 207.100 182.725 ;
        RECT 209.895 182.555 214.990 182.805 ;
        RECT 215.000 182.555 216.370 183.335 ;
        RECT 218.165 183.235 221.395 183.405 ;
        RECT 224.470 183.465 225.390 183.485 ;
        RECT 224.470 183.235 226.490 183.465 ;
        RECT 216.840 182.805 226.490 183.235 ;
        RECT 216.840 182.770 220.035 182.805 ;
        RECT 216.840 182.725 219.095 182.770 ;
        RECT 216.840 182.555 218.600 182.725 ;
        RECT 221.395 182.555 226.490 182.805 ;
        RECT 226.510 182.640 226.940 183.425 ;
        RECT 226.960 182.555 228.330 183.335 ;
        RECT 228.340 182.555 229.710 183.335 ;
        RECT 229.720 182.555 231.090 183.335 ;
        RECT 231.100 182.555 232.470 183.335 ;
        RECT 232.480 182.555 233.850 183.335 ;
        RECT 234.780 182.555 236.150 183.365 ;
        RECT 162.240 182.345 162.410 182.555 ;
        RECT 163.615 182.500 163.735 182.505 ;
        RECT 163.615 182.395 163.790 182.500 ;
        RECT 163.630 182.390 163.790 182.395 ;
        RECT 164.080 182.365 164.250 182.555 ;
        RECT 165.460 182.365 165.630 182.555 ;
        RECT 167.760 182.345 167.930 182.535 ;
        RECT 170.055 182.365 170.225 182.555 ;
        RECT 171.445 182.535 171.615 182.555 ;
        RECT 170.530 182.400 170.690 182.510 ;
        RECT 171.440 182.365 171.615 182.535 ;
        RECT 171.440 182.345 171.610 182.365 ;
        RECT 175.120 182.345 175.290 182.535 ;
        RECT 178.800 182.345 178.970 182.555 ;
        RECT 179.255 182.395 179.375 182.505 ;
        RECT 179.720 182.365 179.890 182.555 ;
        RECT 179.995 182.345 180.165 182.535 ;
        RECT 182.020 182.365 182.190 182.555 ;
        RECT 182.480 182.365 182.650 182.555 ;
        RECT 183.860 182.365 184.030 182.555 ;
        RECT 184.135 182.345 184.305 182.535 ;
        RECT 185.240 182.365 185.410 182.555 ;
        RECT 186.625 182.365 186.795 182.555 ;
        RECT 188.455 182.395 188.575 182.505 ;
        RECT 188.925 182.365 189.095 182.555 ;
        RECT 189.195 182.345 189.365 182.535 ;
        RECT 192.605 182.365 192.775 182.555 ;
        RECT 193.055 182.395 193.175 182.505 ;
        RECT 193.795 182.345 193.965 182.535 ;
        RECT 196.555 182.365 196.725 182.555 ;
        RECT 197.670 182.390 197.830 182.500 ;
        RECT 199.500 182.345 199.670 182.535 ;
        RECT 199.960 182.345 200.130 182.535 ;
        RECT 200.415 182.395 200.535 182.505 ;
        RECT 201.340 182.345 201.510 182.535 ;
        RECT 202.260 182.365 202.430 182.555 ;
        RECT 202.720 182.345 202.890 182.535 ;
        RECT 203.640 182.365 203.810 182.555 ;
        RECT 204.100 182.345 204.270 182.555 ;
        RECT 205.480 182.365 205.650 182.555 ;
        RECT 214.220 182.345 214.390 182.535 ;
        RECT 215.140 182.365 215.310 182.555 ;
        RECT 216.515 182.395 216.635 182.505 ;
        RECT 216.980 182.365 217.150 182.555 ;
        RECT 223.880 182.345 224.050 182.535 ;
        RECT 228.020 182.365 228.190 182.555 ;
        RECT 229.400 182.365 229.570 182.555 ;
        RECT 230.780 182.365 230.950 182.555 ;
        RECT 232.160 182.365 232.330 182.555 ;
        RECT 233.540 182.365 233.710 182.555 ;
        RECT 234.010 182.400 234.170 182.510 ;
        RECT 234.460 182.345 234.630 182.535 ;
        RECT 235.840 182.345 236.010 182.555 ;
      LAYER nwell ;
        RECT 101.175 179.570 156.750 182.070 ;
      LAYER pwell ;
        RECT 162.100 181.535 163.470 182.345 ;
        RECT 164.540 181.435 167.990 182.345 ;
        RECT 168.220 181.435 171.670 182.345 ;
        RECT 171.900 181.435 175.350 182.345 ;
        RECT 175.580 181.435 179.030 182.345 ;
        RECT 179.580 181.665 183.480 182.345 ;
        RECT 183.720 181.665 187.620 182.345 ;
        RECT 179.580 181.435 180.510 181.665 ;
        RECT 183.720 181.435 184.650 181.665 ;
        RECT 187.870 181.475 188.300 182.260 ;
        RECT 188.780 181.665 192.680 182.345 ;
        RECT 193.380 181.665 197.280 182.345 ;
        RECT 188.780 181.435 189.710 181.665 ;
        RECT 193.380 181.435 194.310 181.665 ;
        RECT 198.440 181.565 199.810 182.345 ;
        RECT 199.820 181.565 201.190 182.345 ;
        RECT 201.200 181.565 202.570 182.345 ;
        RECT 202.580 181.565 203.950 182.345 ;
        RECT 203.960 182.175 205.720 182.345 ;
        RECT 203.960 182.130 206.215 182.175 ;
        RECT 203.960 182.095 207.155 182.130 ;
        RECT 208.515 182.095 213.610 182.345 ;
        RECT 203.960 181.665 213.610 182.095 ;
        RECT 205.285 181.495 208.515 181.665 ;
        RECT 206.225 181.450 208.515 181.495 ;
        RECT 207.165 181.415 208.515 181.450 ;
        RECT 211.590 181.435 213.610 181.665 ;
        RECT 213.630 181.475 214.060 182.260 ;
        RECT 214.080 182.175 215.840 182.345 ;
        RECT 214.080 182.130 216.335 182.175 ;
        RECT 214.080 182.095 217.275 182.130 ;
        RECT 218.635 182.095 223.730 182.345 ;
        RECT 214.080 181.665 223.730 182.095 ;
        RECT 223.740 182.175 225.500 182.345 ;
        RECT 223.740 182.130 225.995 182.175 ;
        RECT 223.740 182.095 226.935 182.130 ;
        RECT 228.295 182.095 233.390 182.345 ;
        RECT 223.740 181.665 233.390 182.095 ;
        RECT 215.405 181.495 218.635 181.665 ;
        RECT 216.345 181.450 218.635 181.495 ;
        RECT 211.590 181.415 212.510 181.435 ;
        RECT 217.285 181.415 218.635 181.450 ;
        RECT 221.710 181.435 223.730 181.665 ;
        RECT 225.065 181.495 228.295 181.665 ;
        RECT 226.005 181.450 228.295 181.495 ;
        RECT 221.710 181.415 222.630 181.435 ;
        RECT 226.945 181.415 228.295 181.450 ;
        RECT 231.370 181.435 233.390 181.665 ;
        RECT 233.400 181.565 234.770 182.345 ;
        RECT 234.780 181.535 236.150 182.345 ;
        RECT 231.370 181.415 232.290 181.435 ;
        RECT 9.140 147.810 51.970 168.220 ;
      LAYER nwell ;
        RECT 63.050 164.975 97.990 167.475 ;
      LAYER pwell ;
        RECT 9.600 134.835 20.550 138.315 ;
        RECT 23.425 135.385 58.475 143.515 ;
      LAYER nwell ;
        RECT 63.050 135.035 65.550 164.975 ;
        RECT 69.300 160.385 91.740 161.225 ;
        RECT 69.300 139.625 70.140 160.385 ;
      LAYER pwell ;
        RECT 71.090 158.670 89.950 159.435 ;
        RECT 71.090 156.220 71.855 158.670 ;
        RECT 74.305 156.220 75.575 158.670 ;
        RECT 78.025 156.220 79.295 158.670 ;
        RECT 81.745 156.220 83.015 158.670 ;
        RECT 85.465 156.220 86.735 158.670 ;
        RECT 89.185 156.220 89.950 158.670 ;
        RECT 71.090 154.950 89.950 156.220 ;
        RECT 71.090 152.500 71.855 154.950 ;
        RECT 74.305 152.500 75.575 154.950 ;
        RECT 78.025 152.500 79.295 154.950 ;
        RECT 81.745 152.500 83.015 154.950 ;
        RECT 85.465 152.500 86.735 154.950 ;
        RECT 89.185 152.500 89.950 154.950 ;
        RECT 71.090 151.230 89.950 152.500 ;
        RECT 71.090 148.780 71.855 151.230 ;
        RECT 74.305 148.780 75.575 151.230 ;
        RECT 78.025 148.780 79.295 151.230 ;
        RECT 81.745 148.780 83.015 151.230 ;
        RECT 85.465 148.780 86.735 151.230 ;
        RECT 89.185 148.780 89.950 151.230 ;
        RECT 71.090 147.510 89.950 148.780 ;
        RECT 71.090 145.060 71.855 147.510 ;
        RECT 74.305 145.060 75.575 147.510 ;
        RECT 78.025 145.060 79.295 147.510 ;
        RECT 81.745 145.060 83.015 147.510 ;
        RECT 85.465 145.060 86.735 147.510 ;
        RECT 89.185 145.060 89.950 147.510 ;
        RECT 71.090 143.790 89.950 145.060 ;
        RECT 71.090 141.340 71.855 143.790 ;
        RECT 74.305 141.340 75.575 143.790 ;
        RECT 78.025 141.340 79.295 143.790 ;
        RECT 81.745 141.340 83.015 143.790 ;
        RECT 85.465 141.340 86.735 143.790 ;
        RECT 89.185 141.340 89.950 143.790 ;
        RECT 71.090 140.575 89.950 141.340 ;
      LAYER nwell ;
        RECT 90.900 139.625 91.740 160.385 ;
        RECT 69.300 138.785 91.740 139.625 ;
        RECT 95.490 135.035 97.990 164.975 ;
      LAYER pwell ;
        RECT 102.550 158.280 111.160 172.690 ;
        RECT 114.030 166.235 151.540 176.715 ;
      LAYER nwell ;
        RECT 102.350 141.345 111.360 156.335 ;
        RECT 115.985 139.690 149.475 158.060 ;
        RECT 63.050 132.535 97.990 135.035 ;
        RECT 138.080 129.720 145.960 134.690 ;
      LAYER pwell ;
        RECT 138.280 124.290 145.760 128.770 ;
      LAYER nwell ;
        RECT 10.025 41.635 128.935 124.285 ;
      LAYER pwell ;
        RECT 10.225 9.090 74.495 39.430 ;
        RECT 79.865 9.090 128.735 39.430 ;
      LAYER nwell ;
        RECT 135.120 13.460 149.570 109.050 ;
        RECT 154.250 5.750 156.750 179.570 ;
        RECT 161.905 178.315 236.345 181.145 ;
      LAYER pwell ;
        RECT 205.060 178.025 205.980 178.045 ;
        RECT 162.100 177.115 163.470 177.925 ;
        RECT 163.965 177.795 165.310 178.025 ;
        RECT 163.480 177.115 165.310 177.795 ;
        RECT 165.780 177.115 167.150 177.895 ;
        RECT 167.615 177.345 169.450 178.025 ;
        RECT 167.615 177.115 169.305 177.345 ;
        RECT 169.460 177.115 170.830 177.895 ;
        RECT 170.840 177.115 172.210 177.895 ;
        RECT 172.220 177.115 173.590 177.895 ;
        RECT 173.600 177.115 174.970 177.895 ;
        RECT 174.990 177.200 175.420 177.985 ;
        RECT 175.440 177.345 177.275 178.025 ;
        RECT 175.585 177.115 177.275 177.345 ;
        RECT 178.200 177.115 179.570 177.895 ;
        RECT 179.580 177.115 180.950 177.895 ;
        RECT 180.960 177.115 182.330 177.895 ;
        RECT 182.340 177.795 183.270 178.025 ;
        RECT 182.340 177.115 186.240 177.795 ;
        RECT 186.480 177.115 187.850 177.895 ;
        RECT 187.870 177.200 188.300 177.985 ;
        RECT 188.320 177.345 190.155 178.025 ;
        RECT 190.620 177.345 192.455 178.025 ;
        RECT 188.465 177.115 190.155 177.345 ;
        RECT 190.765 177.115 192.455 177.345 ;
        RECT 192.920 177.795 193.850 178.025 ;
        RECT 192.920 177.115 196.820 177.795 ;
        RECT 197.980 177.115 199.350 177.895 ;
        RECT 199.360 177.115 200.730 177.895 ;
        RECT 200.750 177.200 201.180 177.985 ;
        RECT 201.660 177.115 203.030 177.895 ;
        RECT 203.960 177.795 205.980 178.025 ;
        RECT 209.055 178.010 210.405 178.045 ;
        RECT 220.045 178.010 221.395 178.045 ;
        RECT 209.055 177.965 211.345 178.010 ;
        RECT 209.055 177.795 212.285 177.965 ;
        RECT 203.960 177.365 213.610 177.795 ;
        RECT 203.960 177.115 209.055 177.365 ;
        RECT 210.415 177.330 213.610 177.365 ;
        RECT 211.355 177.285 213.610 177.330 ;
        RECT 211.850 177.115 213.610 177.285 ;
        RECT 213.630 177.200 214.060 177.985 ;
        RECT 219.105 177.965 221.395 178.010 ;
        RECT 214.080 177.115 215.450 177.895 ;
        RECT 215.460 177.115 216.830 177.895 ;
        RECT 218.165 177.795 221.395 177.965 ;
        RECT 224.470 178.025 225.390 178.045 ;
        RECT 224.470 177.795 226.490 178.025 ;
        RECT 216.840 177.365 226.490 177.795 ;
        RECT 216.840 177.330 220.035 177.365 ;
        RECT 216.840 177.285 219.095 177.330 ;
        RECT 216.840 177.115 218.600 177.285 ;
        RECT 221.395 177.115 226.490 177.365 ;
        RECT 226.510 177.200 226.940 177.985 ;
        RECT 226.960 177.115 228.330 177.895 ;
        RECT 228.340 177.115 229.710 177.895 ;
        RECT 229.720 177.115 231.090 177.895 ;
        RECT 231.100 177.115 232.470 177.895 ;
        RECT 232.480 177.115 233.850 177.895 ;
        RECT 234.780 177.115 236.150 177.925 ;
        RECT 162.240 176.925 162.410 177.115 ;
        RECT 163.620 176.925 163.790 177.115 ;
        RECT 165.455 176.955 165.575 177.065 ;
        RECT 165.920 176.925 166.090 177.115 ;
        RECT 169.135 176.925 169.305 177.115 ;
        RECT 169.600 176.925 169.770 177.115 ;
        RECT 170.980 176.925 171.150 177.115 ;
        RECT 172.360 176.925 172.530 177.115 ;
        RECT 173.740 176.925 173.910 177.115 ;
        RECT 175.585 176.925 175.755 177.115 ;
        RECT 177.875 176.955 177.995 177.065 ;
        RECT 178.340 176.925 178.510 177.115 ;
        RECT 179.720 176.925 179.890 177.115 ;
        RECT 181.100 176.925 181.270 177.115 ;
        RECT 182.755 176.925 182.925 177.115 ;
        RECT 186.620 176.925 186.790 177.115 ;
        RECT 188.465 176.925 188.635 177.115 ;
        RECT 190.765 176.925 190.935 177.115 ;
        RECT 193.335 176.925 193.505 177.115 ;
        RECT 197.210 176.960 197.370 177.070 ;
        RECT 198.120 176.925 198.290 177.115 ;
        RECT 199.500 176.925 199.670 177.115 ;
        RECT 201.335 176.955 201.455 177.065 ;
        RECT 201.800 176.925 201.970 177.115 ;
        RECT 203.190 176.960 203.350 177.070 ;
        RECT 213.300 176.925 213.470 177.115 ;
        RECT 214.220 176.925 214.390 177.115 ;
        RECT 215.600 176.925 215.770 177.115 ;
        RECT 216.980 176.925 217.150 177.115 ;
        RECT 228.020 176.925 228.190 177.115 ;
        RECT 229.400 176.925 229.570 177.115 ;
        RECT 230.780 176.925 230.950 177.115 ;
        RECT 232.160 176.925 232.330 177.115 ;
        RECT 233.540 176.925 233.710 177.115 ;
        RECT 234.010 176.960 234.170 177.070 ;
        RECT 235.840 176.925 236.010 177.115 ;
        RECT 162.240 106.320 162.410 106.510 ;
        RECT 165.000 106.320 165.170 106.510 ;
        RECT 166.840 106.320 167.010 106.510 ;
        RECT 168.680 106.320 168.850 106.510 ;
        RECT 170.520 106.320 170.690 106.510 ;
        RECT 171.255 106.320 171.425 106.510 ;
        RECT 175.855 106.320 176.025 106.510 ;
        RECT 179.730 106.365 179.890 106.475 ;
        RECT 180.640 106.320 180.810 106.510 ;
        RECT 182.480 106.320 182.650 106.510 ;
        RECT 184.320 106.320 184.490 106.510 ;
        RECT 186.160 106.320 186.330 106.510 ;
        RECT 188.455 106.370 188.575 106.480 ;
        RECT 189.195 106.320 189.365 106.510 ;
        RECT 193.055 106.370 193.175 106.480 ;
        RECT 193.520 106.320 193.690 106.510 ;
        RECT 195.360 106.320 195.530 106.510 ;
        RECT 197.200 106.320 197.370 106.510 ;
        RECT 199.040 106.320 199.210 106.510 ;
        RECT 201.340 106.320 201.510 106.510 ;
        RECT 202.720 106.320 202.890 106.510 ;
        RECT 205.940 106.320 206.110 106.510 ;
        RECT 206.675 106.320 206.845 106.510 ;
        RECT 210.540 106.320 210.710 106.510 ;
        RECT 213.300 106.320 213.470 106.510 ;
        RECT 214.220 106.320 214.390 106.510 ;
        RECT 216.980 106.320 217.150 106.510 ;
        RECT 217.440 106.320 217.610 106.510 ;
        RECT 219.555 106.320 219.725 106.510 ;
        RECT 223.420 106.320 223.590 106.510 ;
        RECT 226.180 106.320 226.350 106.510 ;
        RECT 230.320 106.320 230.490 106.510 ;
        RECT 230.775 106.370 230.895 106.480 ;
        RECT 232.620 106.320 232.790 106.510 ;
        RECT 233.075 106.370 233.195 106.480 ;
        RECT 234.920 106.320 235.090 106.510 ;
        RECT 235.375 106.370 235.495 106.480 ;
        RECT 237.220 106.320 237.390 106.510 ;
        RECT 239.060 106.320 239.230 106.510 ;
        RECT 239.975 106.370 240.095 106.480 ;
        RECT 240.715 106.320 240.885 106.510 ;
        RECT 244.580 106.320 244.750 106.510 ;
        RECT 251.480 106.320 251.650 106.510 ;
        RECT 251.935 106.370 252.055 106.480 ;
        RECT 252.870 106.365 253.030 106.475 ;
        RECT 257.000 106.320 257.170 106.510 ;
        RECT 257.460 106.320 257.630 106.510 ;
        RECT 260.680 106.320 260.850 106.510 ;
        RECT 262.520 106.320 262.690 106.510 ;
        RECT 264.360 106.320 264.530 106.510 ;
        RECT 264.815 106.370 264.935 106.480 ;
        RECT 267.120 106.320 267.290 106.510 ;
        RECT 268.960 106.320 269.130 106.510 ;
        RECT 269.420 106.320 269.590 106.510 ;
        RECT 274.480 106.320 274.650 106.510 ;
        RECT 274.940 106.320 275.110 106.510 ;
        RECT 276.780 106.320 276.950 106.510 ;
        RECT 280.000 106.320 280.170 106.510 ;
        RECT 281.840 106.320 282.010 106.510 ;
        RECT 283.680 106.320 283.850 106.510 ;
        RECT 285.520 106.320 285.690 106.510 ;
        RECT 287.360 106.320 287.530 106.510 ;
        RECT 289.200 106.320 289.370 106.510 ;
        RECT 289.660 106.320 289.830 106.510 ;
        RECT 292.880 106.320 293.050 106.510 ;
        RECT 293.340 106.320 293.510 106.510 ;
        RECT 294.720 106.320 294.890 106.510 ;
        RECT 304.380 106.320 304.550 106.510 ;
        RECT 306.220 106.320 306.390 106.510 ;
        RECT 308.060 106.320 308.230 106.510 ;
        RECT 310.820 106.320 310.990 106.510 ;
        RECT 162.100 105.510 163.470 106.320 ;
        RECT 163.480 105.640 165.310 106.320 ;
        RECT 165.320 105.640 167.150 106.320 ;
        RECT 167.160 105.640 168.990 106.320 ;
        RECT 169.000 105.640 170.830 106.320 ;
        RECT 170.840 105.640 174.740 106.320 ;
        RECT 163.480 105.410 164.825 105.640 ;
        RECT 165.320 105.410 166.665 105.640 ;
        RECT 167.160 105.410 168.505 105.640 ;
        RECT 169.000 105.410 170.345 105.640 ;
        RECT 170.840 105.410 171.770 105.640 ;
        RECT 174.990 105.450 175.420 106.235 ;
        RECT 175.440 105.640 179.340 106.320 ;
        RECT 180.500 105.640 182.330 106.320 ;
        RECT 182.340 105.640 184.170 106.320 ;
        RECT 184.180 105.640 186.010 106.320 ;
        RECT 186.020 105.640 187.850 106.320 ;
        RECT 175.440 105.410 176.370 105.640 ;
        RECT 180.985 105.410 182.330 105.640 ;
        RECT 182.825 105.410 184.170 105.640 ;
        RECT 184.665 105.410 186.010 105.640 ;
        RECT 186.505 105.410 187.850 105.640 ;
        RECT 187.870 105.450 188.300 106.235 ;
        RECT 188.780 105.640 192.680 106.320 ;
        RECT 193.380 105.640 195.210 106.320 ;
        RECT 195.220 105.640 197.050 106.320 ;
        RECT 197.060 105.640 198.890 106.320 ;
        RECT 198.900 105.640 200.730 106.320 ;
        RECT 188.780 105.410 189.710 105.640 ;
        RECT 193.865 105.410 195.210 105.640 ;
        RECT 195.705 105.410 197.050 105.640 ;
        RECT 197.545 105.410 198.890 105.640 ;
        RECT 199.385 105.410 200.730 105.640 ;
        RECT 200.750 105.450 201.180 106.235 ;
        RECT 201.200 105.510 202.570 106.320 ;
        RECT 202.580 105.640 204.410 106.320 ;
        RECT 203.065 105.410 204.410 105.640 ;
        RECT 204.420 105.640 206.250 106.320 ;
        RECT 206.260 105.640 210.160 106.320 ;
        RECT 204.420 105.410 205.765 105.640 ;
        RECT 206.260 105.410 207.190 105.640 ;
        RECT 210.400 105.510 211.770 106.320 ;
        RECT 211.780 105.640 213.610 106.320 ;
        RECT 211.780 105.410 213.125 105.640 ;
        RECT 213.630 105.450 214.060 106.235 ;
        RECT 214.080 105.510 215.450 106.320 ;
        RECT 215.460 105.640 217.290 106.320 ;
        RECT 217.300 105.640 219.130 106.320 ;
        RECT 215.460 105.410 216.805 105.640 ;
        RECT 217.785 105.410 219.130 105.640 ;
        RECT 219.140 105.640 223.040 106.320 ;
        RECT 219.140 105.410 220.070 105.640 ;
        RECT 223.280 105.510 224.650 106.320 ;
        RECT 224.660 105.640 226.490 106.320 ;
        RECT 224.660 105.410 226.005 105.640 ;
        RECT 226.510 105.450 226.940 106.235 ;
        RECT 227.055 105.640 230.520 106.320 ;
        RECT 231.100 105.640 232.930 106.320 ;
        RECT 233.400 105.640 235.230 106.320 ;
        RECT 235.700 105.640 237.530 106.320 ;
        RECT 237.540 105.640 239.370 106.320 ;
        RECT 227.055 105.410 227.975 105.640 ;
        RECT 231.100 105.410 232.445 105.640 ;
        RECT 233.400 105.410 234.745 105.640 ;
        RECT 235.700 105.410 237.045 105.640 ;
        RECT 237.540 105.410 238.885 105.640 ;
        RECT 239.390 105.450 239.820 106.235 ;
        RECT 240.300 105.640 244.200 106.320 ;
        RECT 244.550 105.640 248.015 106.320 ;
        RECT 240.300 105.410 241.230 105.640 ;
        RECT 247.095 105.410 248.015 105.640 ;
        RECT 248.215 105.640 251.680 106.320 ;
        RECT 248.215 105.410 249.135 105.640 ;
        RECT 252.270 105.450 252.700 106.235 ;
        RECT 253.735 105.640 257.200 106.320 ;
        RECT 257.320 105.640 259.150 106.320 ;
        RECT 253.735 105.410 254.655 105.640 ;
        RECT 257.805 105.410 259.150 105.640 ;
        RECT 259.160 105.640 260.990 106.320 ;
        RECT 261.000 105.640 262.830 106.320 ;
        RECT 262.840 105.640 264.670 106.320 ;
        RECT 259.160 105.410 260.505 105.640 ;
        RECT 261.000 105.410 262.345 105.640 ;
        RECT 262.840 105.410 264.185 105.640 ;
        RECT 265.150 105.450 265.580 106.235 ;
        RECT 265.600 105.640 267.430 106.320 ;
        RECT 267.440 105.640 269.270 106.320 ;
        RECT 269.390 105.640 272.855 106.320 ;
        RECT 265.600 105.410 266.945 105.640 ;
        RECT 267.440 105.410 268.785 105.640 ;
        RECT 271.935 105.410 272.855 105.640 ;
        RECT 272.960 105.640 274.790 106.320 ;
        RECT 274.800 105.640 276.630 106.320 ;
        RECT 272.960 105.410 274.305 105.640 ;
        RECT 275.285 105.410 276.630 105.640 ;
        RECT 276.640 105.510 278.010 106.320 ;
        RECT 278.030 105.450 278.460 106.235 ;
        RECT 278.480 105.640 280.310 106.320 ;
        RECT 280.320 105.640 282.150 106.320 ;
        RECT 282.160 105.640 283.990 106.320 ;
        RECT 284.000 105.640 285.830 106.320 ;
        RECT 285.840 105.640 287.670 106.320 ;
        RECT 287.680 105.640 289.510 106.320 ;
        RECT 278.480 105.410 279.825 105.640 ;
        RECT 280.320 105.410 281.665 105.640 ;
        RECT 282.160 105.410 283.505 105.640 ;
        RECT 284.000 105.410 285.345 105.640 ;
        RECT 285.840 105.410 287.185 105.640 ;
        RECT 287.680 105.410 289.025 105.640 ;
        RECT 289.520 105.510 290.890 106.320 ;
        RECT 290.910 105.450 291.340 106.235 ;
        RECT 291.360 105.640 293.190 106.320 ;
        RECT 291.360 105.410 292.705 105.640 ;
        RECT 293.200 105.510 294.570 106.320 ;
        RECT 294.580 105.640 303.770 106.320 ;
        RECT 299.090 105.420 300.020 105.640 ;
        RECT 302.850 105.410 303.770 105.640 ;
        RECT 303.790 105.450 304.220 106.235 ;
        RECT 304.240 105.640 306.070 106.320 ;
        RECT 306.080 105.640 307.910 106.320 ;
        RECT 307.920 105.640 309.750 106.320 ;
        RECT 304.725 105.410 306.070 105.640 ;
        RECT 306.565 105.410 307.910 105.640 ;
        RECT 308.405 105.410 309.750 105.640 ;
        RECT 309.760 105.510 311.130 106.320 ;
      LAYER nwell ;
        RECT 161.905 102.290 311.325 105.120 ;
      LAYER pwell ;
        RECT 162.100 101.090 163.470 101.900 ;
        RECT 163.940 101.770 165.285 102.000 ;
        RECT 170.290 101.770 171.220 101.990 ;
        RECT 174.050 101.770 174.970 102.000 ;
        RECT 163.940 101.090 165.770 101.770 ;
        RECT 165.780 101.090 174.970 101.770 ;
        RECT 174.990 101.175 175.420 101.960 ;
        RECT 175.440 101.090 176.810 101.900 ;
        RECT 181.330 101.770 182.260 101.990 ;
        RECT 185.090 101.770 186.010 102.000 ;
        RECT 190.530 101.770 191.460 101.990 ;
        RECT 194.290 101.770 195.210 102.000 ;
        RECT 176.820 101.090 186.010 101.770 ;
        RECT 186.020 101.090 195.210 101.770 ;
        RECT 195.220 101.770 196.150 102.000 ;
        RECT 195.220 101.090 199.120 101.770 ;
        RECT 199.360 101.090 200.730 101.900 ;
        RECT 200.750 101.175 201.180 101.960 ;
        RECT 201.685 101.770 203.030 102.000 ;
        RECT 207.550 101.770 208.480 101.990 ;
        RECT 211.310 101.770 212.230 102.000 ;
        RECT 201.200 101.090 203.030 101.770 ;
        RECT 203.040 101.090 212.230 101.770 ;
        RECT 212.240 101.770 213.170 102.000 ;
        RECT 221.810 101.770 222.740 101.990 ;
        RECT 225.570 101.770 226.490 102.000 ;
        RECT 212.240 101.090 216.140 101.770 ;
        RECT 217.300 101.090 226.490 101.770 ;
        RECT 226.510 101.175 226.940 101.960 ;
        RECT 226.960 101.770 227.890 102.000 ;
        RECT 231.100 101.770 232.445 102.000 ;
        RECT 226.960 101.090 230.860 101.770 ;
        RECT 231.100 101.090 232.930 101.770 ;
        RECT 232.940 101.090 236.610 101.900 ;
        RECT 241.130 101.770 242.060 101.990 ;
        RECT 244.890 101.770 245.810 102.000 ;
        RECT 236.620 101.090 245.810 101.770 ;
        RECT 245.820 101.770 246.750 102.000 ;
        RECT 249.960 101.770 251.305 102.000 ;
        RECT 245.820 101.090 249.720 101.770 ;
        RECT 249.960 101.090 251.790 101.770 ;
        RECT 252.270 101.175 252.700 101.960 ;
        RECT 257.230 101.770 258.160 101.990 ;
        RECT 260.990 101.770 261.910 102.000 ;
        RECT 266.430 101.770 267.360 101.990 ;
        RECT 270.190 101.770 271.110 102.000 ;
        RECT 274.320 101.770 275.250 102.000 ;
        RECT 252.720 101.090 261.910 101.770 ;
        RECT 261.920 101.090 271.110 101.770 ;
        RECT 271.350 101.090 275.250 101.770 ;
        RECT 275.260 101.770 276.605 102.000 ;
        RECT 275.260 101.090 277.090 101.770 ;
        RECT 278.030 101.175 278.460 101.960 ;
        RECT 278.480 101.770 279.400 102.000 ;
        RECT 282.230 101.770 283.160 101.990 ;
        RECT 293.110 101.770 294.040 101.990 ;
        RECT 296.870 101.770 297.790 102.000 ;
        RECT 278.480 101.090 287.670 101.770 ;
        RECT 288.600 101.090 297.790 101.770 ;
        RECT 297.800 101.770 298.730 102.000 ;
        RECT 302.425 101.770 303.770 102.000 ;
        RECT 297.800 101.090 301.700 101.770 ;
        RECT 301.940 101.090 303.770 101.770 ;
        RECT 303.790 101.175 304.220 101.960 ;
        RECT 304.240 101.770 305.170 102.000 ;
        RECT 304.240 101.090 308.140 101.770 ;
        RECT 308.380 101.090 309.750 101.900 ;
        RECT 309.760 101.090 311.130 101.900 ;
        RECT 162.240 100.880 162.410 101.090 ;
        RECT 163.615 100.930 163.735 101.040 ;
        RECT 165.000 100.880 165.170 101.070 ;
        RECT 165.460 100.880 165.630 101.090 ;
        RECT 165.920 100.900 166.090 101.090 ;
        RECT 167.300 100.880 167.470 101.070 ;
        RECT 175.580 100.900 175.750 101.090 ;
        RECT 176.775 100.880 176.945 101.070 ;
        RECT 176.960 100.900 177.130 101.090 ;
        RECT 182.020 100.880 182.190 101.070 ;
        RECT 182.475 100.930 182.595 101.040 ;
        RECT 184.320 100.880 184.490 101.070 ;
        RECT 184.775 100.930 184.895 101.040 ;
        RECT 186.160 100.900 186.330 101.090 ;
        RECT 186.620 100.880 186.790 101.070 ;
        RECT 187.090 100.925 187.250 101.035 ;
        RECT 188.460 100.880 188.630 101.070 ;
        RECT 195.635 100.900 195.805 101.090 ;
        RECT 197.660 100.880 197.830 101.070 ;
        RECT 199.500 100.900 199.670 101.090 ;
        RECT 201.340 100.880 201.510 101.090 ;
        RECT 203.180 100.900 203.350 101.090 ;
        RECT 211.460 100.880 211.630 101.070 ;
        RECT 212.655 100.900 212.825 101.090 ;
        RECT 213.300 100.880 213.470 101.070 ;
        RECT 214.230 100.925 214.390 101.035 ;
        RECT 216.520 100.880 216.690 101.070 ;
        RECT 216.975 100.930 217.095 101.040 ;
        RECT 217.440 100.880 217.610 101.090 ;
        RECT 226.640 100.880 226.810 101.070 ;
        RECT 227.375 100.900 227.545 101.090 ;
        RECT 228.025 100.880 228.195 101.070 ;
        RECT 231.700 100.880 231.870 101.070 ;
        RECT 232.620 100.900 232.790 101.090 ;
        RECT 233.080 100.900 233.250 101.090 ;
        RECT 236.760 100.900 236.930 101.090 ;
        RECT 237.220 100.880 237.390 101.070 ;
        RECT 239.055 100.930 239.175 101.040 ;
        RECT 239.980 100.880 240.150 101.070 ;
        RECT 246.235 100.900 246.405 101.090 ;
        RECT 249.180 100.880 249.350 101.070 ;
        RECT 251.480 100.900 251.650 101.090 ;
        RECT 251.935 100.930 252.055 101.040 ;
        RECT 252.675 100.880 252.845 101.070 ;
        RECT 252.860 100.900 253.030 101.090 ;
        RECT 257.920 100.880 258.090 101.070 ;
        RECT 261.785 100.880 261.955 101.070 ;
        RECT 262.060 100.900 262.230 101.090 ;
        RECT 263.900 100.880 264.070 101.070 ;
        RECT 264.370 100.925 264.530 101.035 ;
        RECT 274.480 100.880 274.650 101.070 ;
        RECT 274.665 100.900 274.835 101.090 ;
        RECT 274.940 100.880 275.110 101.070 ;
        RECT 276.780 100.900 276.950 101.090 ;
        RECT 277.250 100.935 277.410 101.045 ;
        RECT 287.360 100.900 287.530 101.090 ;
        RECT 287.545 100.880 287.715 101.070 ;
        RECT 287.830 100.935 287.990 101.045 ;
        RECT 288.280 100.880 288.450 101.070 ;
        RECT 288.740 100.900 288.910 101.090 ;
        RECT 290.130 100.925 290.290 101.035 ;
        RECT 291.500 100.880 291.670 101.070 ;
        RECT 293.335 100.930 293.455 101.040 ;
        RECT 293.800 100.880 293.970 101.070 ;
        RECT 298.215 100.900 298.385 101.090 ;
        RECT 302.080 100.900 302.250 101.090 ;
        RECT 304.380 100.880 304.550 101.070 ;
        RECT 304.655 100.900 304.825 101.090 ;
        RECT 304.840 100.880 305.010 101.070 ;
        RECT 306.675 100.930 306.795 101.040 ;
        RECT 307.140 100.880 307.310 101.070 ;
        RECT 308.520 100.900 308.690 101.090 ;
        RECT 308.990 100.925 309.150 101.035 ;
        RECT 310.820 100.880 310.990 101.090 ;
        RECT 162.100 100.070 163.470 100.880 ;
        RECT 163.480 100.200 165.310 100.880 ;
        RECT 165.320 100.200 167.150 100.880 ;
        RECT 167.160 100.200 176.350 100.880 ;
        RECT 163.480 99.970 164.825 100.200 ;
        RECT 165.805 99.970 167.150 100.200 ;
        RECT 171.670 99.980 172.600 100.200 ;
        RECT 175.430 99.970 176.350 100.200 ;
        RECT 176.360 100.200 180.260 100.880 ;
        RECT 180.500 100.200 182.330 100.880 ;
        RECT 182.800 100.200 184.630 100.880 ;
        RECT 185.100 100.200 186.930 100.880 ;
        RECT 176.360 99.970 177.290 100.200 ;
        RECT 180.500 99.970 181.845 100.200 ;
        RECT 182.800 99.970 184.145 100.200 ;
        RECT 185.100 99.970 186.445 100.200 ;
        RECT 187.870 100.010 188.300 100.795 ;
        RECT 188.320 100.200 197.510 100.880 ;
        RECT 192.830 99.980 193.760 100.200 ;
        RECT 196.590 99.970 197.510 100.200 ;
        RECT 197.520 100.070 201.190 100.880 ;
        RECT 201.200 100.070 202.570 100.880 ;
        RECT 202.580 100.200 211.770 100.880 ;
        RECT 211.780 100.200 213.610 100.880 ;
        RECT 202.580 99.970 203.500 100.200 ;
        RECT 206.330 99.980 207.260 100.200 ;
        RECT 211.780 99.970 213.125 100.200 ;
        RECT 213.630 100.010 214.060 100.795 ;
        RECT 215.000 100.200 216.830 100.880 ;
        RECT 217.300 100.200 226.490 100.880 ;
        RECT 215.000 99.970 216.345 100.200 ;
        RECT 221.810 99.980 222.740 100.200 ;
        RECT 225.570 99.970 226.490 100.200 ;
        RECT 226.500 100.070 227.870 100.880 ;
        RECT 227.880 99.970 231.535 100.880 ;
        RECT 231.560 100.070 237.070 100.880 ;
        RECT 237.080 100.070 238.910 100.880 ;
        RECT 239.390 100.010 239.820 100.795 ;
        RECT 239.840 100.200 249.030 100.880 ;
        RECT 244.350 99.980 245.280 100.200 ;
        RECT 248.110 99.970 249.030 100.200 ;
        RECT 249.040 99.970 252.250 100.880 ;
        RECT 252.260 100.200 256.160 100.880 ;
        RECT 256.400 100.200 258.230 100.880 ;
        RECT 258.470 100.200 262.370 100.880 ;
        RECT 252.260 99.970 253.190 100.200 ;
        RECT 256.400 99.970 257.745 100.200 ;
        RECT 261.440 99.970 262.370 100.200 ;
        RECT 262.380 100.200 264.210 100.880 ;
        RECT 262.380 99.970 263.725 100.200 ;
        RECT 265.150 100.010 265.580 100.795 ;
        RECT 265.600 100.200 274.790 100.880 ;
        RECT 274.800 100.200 283.990 100.880 ;
        RECT 284.230 100.200 288.130 100.880 ;
        RECT 288.140 100.200 289.970 100.880 ;
        RECT 265.600 99.970 266.520 100.200 ;
        RECT 269.350 99.980 270.280 100.200 ;
        RECT 279.310 99.980 280.240 100.200 ;
        RECT 283.070 99.970 283.990 100.200 ;
        RECT 287.200 99.970 288.130 100.200 ;
        RECT 288.625 99.970 289.970 100.200 ;
        RECT 290.910 100.010 291.340 100.795 ;
        RECT 291.360 100.200 293.190 100.880 ;
        RECT 293.660 100.200 302.850 100.880 ;
        RECT 291.845 99.970 293.190 100.200 ;
        RECT 298.170 99.980 299.100 100.200 ;
        RECT 301.930 99.970 302.850 100.200 ;
        RECT 302.860 100.200 304.690 100.880 ;
        RECT 304.700 100.200 306.530 100.880 ;
        RECT 307.000 100.200 308.830 100.880 ;
        RECT 302.860 99.970 304.205 100.200 ;
        RECT 305.185 99.970 306.530 100.200 ;
        RECT 307.485 99.970 308.830 100.200 ;
        RECT 309.760 100.070 311.130 100.880 ;
      LAYER nwell ;
        RECT 161.905 96.850 311.325 99.680 ;
      LAYER pwell ;
        RECT 162.100 95.650 163.470 96.460 ;
        RECT 163.480 96.330 164.825 96.560 ;
        RECT 170.290 96.330 171.220 96.550 ;
        RECT 174.050 96.330 174.970 96.560 ;
        RECT 163.480 95.650 165.310 96.330 ;
        RECT 165.780 95.650 174.970 96.330 ;
        RECT 174.990 95.735 175.420 96.520 ;
        RECT 175.440 96.330 176.370 96.560 ;
        RECT 175.440 95.650 179.340 96.330 ;
        RECT 179.580 95.650 181.410 96.460 ;
        RECT 181.420 95.650 184.170 96.560 ;
        RECT 188.690 96.330 189.620 96.550 ;
        RECT 192.450 96.330 193.370 96.560 ;
        RECT 184.180 95.650 193.370 96.330 ;
        RECT 193.380 96.330 194.310 96.560 ;
        RECT 193.380 95.650 197.280 96.330 ;
        RECT 197.530 95.650 200.270 96.330 ;
        RECT 200.750 95.735 201.180 96.520 ;
        RECT 201.200 95.650 202.570 96.460 ;
        RECT 202.590 95.650 205.320 96.560 ;
        RECT 205.340 95.650 208.550 96.560 ;
        RECT 211.215 96.330 212.135 96.560 ;
        RECT 208.670 95.650 212.135 96.330 ;
        RECT 212.240 95.650 217.750 96.460 ;
        RECT 217.760 95.650 220.510 96.460 ;
        RECT 220.520 95.650 223.270 96.560 ;
        RECT 223.280 95.650 226.490 96.560 ;
        RECT 226.510 95.735 226.940 96.520 ;
        RECT 226.975 95.650 230.630 96.560 ;
        RECT 230.640 95.650 236.150 96.460 ;
        RECT 236.160 95.650 241.670 96.460 ;
        RECT 241.680 95.650 243.050 96.460 ;
        RECT 243.060 95.650 246.270 96.560 ;
        RECT 246.280 95.650 249.935 96.560 ;
        RECT 249.960 95.650 251.790 96.460 ;
        RECT 252.270 95.735 252.700 96.520 ;
        RECT 252.735 95.650 256.390 96.560 ;
        RECT 257.320 95.650 260.520 96.560 ;
        RECT 260.540 95.650 266.050 96.460 ;
        RECT 266.060 95.650 271.570 96.460 ;
        RECT 271.580 95.650 273.410 96.460 ;
        RECT 277.080 96.330 278.010 96.560 ;
        RECT 274.110 95.650 278.010 96.330 ;
        RECT 278.030 95.735 278.460 96.520 ;
        RECT 283.450 96.330 284.380 96.550 ;
        RECT 287.210 96.330 288.130 96.560 ;
        RECT 288.625 96.330 289.970 96.560 ;
        RECT 278.940 95.650 288.130 96.330 ;
        RECT 288.140 95.650 289.970 96.330 ;
        RECT 289.980 96.330 290.910 96.560 ;
        RECT 299.090 96.330 300.020 96.550 ;
        RECT 302.850 96.330 303.770 96.560 ;
        RECT 289.980 95.650 293.880 96.330 ;
        RECT 294.580 95.650 303.770 96.330 ;
        RECT 303.790 95.735 304.220 96.520 ;
        RECT 304.240 96.330 305.170 96.560 ;
        RECT 304.240 95.650 308.140 96.330 ;
        RECT 308.380 95.650 309.750 96.460 ;
        RECT 309.760 95.650 311.130 96.460 ;
        RECT 162.240 95.440 162.410 95.650 ;
        RECT 165.000 95.440 165.170 95.650 ;
        RECT 165.460 95.600 165.630 95.630 ;
        RECT 165.455 95.490 165.630 95.600 ;
        RECT 165.460 95.440 165.630 95.490 ;
        RECT 165.920 95.460 166.090 95.650 ;
        RECT 169.140 95.440 169.310 95.630 ;
        RECT 175.855 95.460 176.025 95.650 ;
        RECT 178.800 95.440 178.970 95.630 ;
        RECT 179.720 95.460 179.890 95.650 ;
        RECT 181.560 95.460 181.730 95.650 ;
        RECT 184.320 95.440 184.490 95.650 ;
        RECT 188.735 95.440 188.905 95.630 ;
        RECT 192.600 95.440 192.770 95.630 ;
        RECT 193.795 95.460 193.965 95.650 ;
        RECT 195.360 95.440 195.530 95.630 ;
        RECT 199.960 95.460 200.130 95.650 ;
        RECT 200.415 95.490 200.535 95.600 ;
        RECT 200.880 95.440 201.050 95.630 ;
        RECT 201.340 95.460 201.510 95.650 ;
        RECT 202.720 95.460 202.890 95.650 ;
        RECT 206.400 95.440 206.570 95.630 ;
        RECT 208.240 95.460 208.410 95.650 ;
        RECT 208.700 95.460 208.870 95.650 ;
        RECT 209.160 95.440 209.330 95.630 ;
        RECT 212.380 95.440 212.550 95.650 ;
        RECT 214.220 95.440 214.390 95.630 ;
        RECT 217.900 95.460 218.070 95.650 ;
        RECT 219.740 95.440 219.910 95.630 ;
        RECT 220.660 95.460 220.830 95.650 ;
        RECT 223.420 95.460 223.590 95.650 ;
        RECT 227.100 95.440 227.270 95.630 ;
        RECT 227.560 95.440 227.730 95.630 ;
        RECT 230.315 95.460 230.485 95.650 ;
        RECT 230.780 95.440 230.950 95.650 ;
        RECT 236.300 95.440 236.470 95.650 ;
        RECT 239.055 95.490 239.175 95.600 ;
        RECT 239.980 95.440 240.150 95.630 ;
        RECT 241.820 95.460 241.990 95.650 ;
        RECT 244.575 95.440 244.745 95.630 ;
        RECT 245.040 95.440 245.210 95.630 ;
        RECT 245.960 95.460 246.130 95.650 ;
        RECT 246.425 95.460 246.595 95.650 ;
        RECT 250.100 95.460 250.270 95.650 ;
        RECT 251.475 95.440 251.645 95.630 ;
        RECT 251.940 95.600 252.110 95.630 ;
        RECT 251.935 95.490 252.110 95.600 ;
        RECT 251.940 95.440 252.110 95.490 ;
        RECT 256.075 95.460 256.245 95.650 ;
        RECT 256.550 95.495 256.710 95.605 ;
        RECT 257.470 95.485 257.630 95.595 ;
        RECT 258.385 95.440 258.555 95.630 ;
        RECT 260.225 95.460 260.395 95.650 ;
        RECT 260.680 95.460 260.850 95.650 ;
        RECT 262.060 95.440 262.230 95.630 ;
        RECT 265.740 95.440 265.910 95.630 ;
        RECT 266.200 95.460 266.370 95.650 ;
        RECT 271.260 95.440 271.430 95.630 ;
        RECT 271.720 95.460 271.890 95.650 ;
        RECT 273.555 95.490 273.675 95.600 ;
        RECT 276.775 95.490 276.895 95.600 ;
        RECT 277.240 95.440 277.410 95.630 ;
        RECT 277.425 95.460 277.595 95.650 ;
        RECT 278.615 95.490 278.735 95.600 ;
        RECT 279.080 95.460 279.250 95.650 ;
        RECT 280.275 95.440 280.445 95.630 ;
        RECT 286.440 95.440 286.610 95.630 ;
        RECT 286.900 95.440 287.070 95.630 ;
        RECT 288.280 95.460 288.450 95.650 ;
        RECT 290.395 95.460 290.565 95.650 ;
        RECT 290.575 95.490 290.695 95.600 ;
        RECT 291.510 95.485 291.670 95.595 ;
        RECT 294.255 95.490 294.375 95.600 ;
        RECT 294.720 95.460 294.890 95.650 ;
        RECT 295.825 95.440 295.995 95.630 ;
        RECT 296.560 95.440 296.730 95.630 ;
        RECT 304.655 95.460 304.825 95.650 ;
        RECT 305.755 95.490 305.875 95.600 ;
        RECT 306.220 95.440 306.390 95.630 ;
        RECT 308.060 95.440 308.230 95.630 ;
        RECT 308.520 95.460 308.690 95.650 ;
        RECT 310.820 95.440 310.990 95.650 ;
        RECT 162.100 94.630 163.470 95.440 ;
        RECT 163.480 94.760 165.310 95.440 ;
        RECT 163.480 94.530 164.825 94.760 ;
        RECT 165.320 94.630 168.990 95.440 ;
        RECT 169.000 94.760 178.610 95.440 ;
        RECT 173.510 94.540 174.440 94.760 ;
        RECT 177.270 94.530 178.610 94.760 ;
        RECT 178.660 94.630 184.170 95.440 ;
        RECT 184.180 94.630 187.850 95.440 ;
        RECT 187.870 94.570 188.300 95.355 ;
        RECT 188.320 94.760 192.220 95.440 ;
        RECT 188.320 94.530 189.250 94.760 ;
        RECT 192.460 94.530 195.210 95.440 ;
        RECT 195.220 94.630 200.730 95.440 ;
        RECT 200.740 94.630 206.250 95.440 ;
        RECT 206.270 94.530 209.000 95.440 ;
        RECT 209.020 94.530 212.230 95.440 ;
        RECT 212.240 94.630 213.610 95.440 ;
        RECT 213.630 94.570 214.060 95.355 ;
        RECT 214.080 94.630 219.590 95.440 ;
        RECT 219.600 94.630 223.270 95.440 ;
        RECT 224.200 94.530 227.410 95.440 ;
        RECT 227.420 94.530 230.630 95.440 ;
        RECT 230.640 94.630 236.150 95.440 ;
        RECT 236.160 94.630 238.910 95.440 ;
        RECT 239.390 94.570 239.820 95.355 ;
        RECT 239.840 94.630 241.210 95.440 ;
        RECT 241.235 94.530 244.890 95.440 ;
        RECT 244.900 94.530 248.110 95.440 ;
        RECT 248.135 94.530 251.790 95.440 ;
        RECT 251.800 94.630 257.310 95.440 ;
        RECT 258.240 94.530 261.895 95.440 ;
        RECT 261.920 94.530 265.130 95.440 ;
        RECT 265.150 94.570 265.580 95.355 ;
        RECT 265.600 94.630 271.110 95.440 ;
        RECT 271.120 94.630 276.630 95.440 ;
        RECT 277.100 94.530 279.850 95.440 ;
        RECT 279.860 94.760 283.760 95.440 ;
        RECT 279.860 94.530 280.790 94.760 ;
        RECT 284.000 94.530 286.750 95.440 ;
        RECT 286.760 94.630 290.430 95.440 ;
        RECT 290.910 94.570 291.340 95.355 ;
        RECT 292.510 94.760 296.410 95.440 ;
        RECT 296.420 94.760 305.610 95.440 ;
        RECT 306.080 94.760 307.910 95.440 ;
        RECT 307.920 94.760 309.750 95.440 ;
        RECT 295.480 94.530 296.410 94.760 ;
        RECT 300.930 94.540 301.860 94.760 ;
        RECT 304.690 94.530 305.610 94.760 ;
        RECT 306.565 94.530 307.910 94.760 ;
        RECT 308.405 94.530 309.750 94.760 ;
        RECT 309.760 94.630 311.130 95.440 ;
      LAYER nwell ;
        RECT 161.905 91.410 311.325 94.240 ;
      LAYER pwell ;
        RECT 162.100 90.210 163.470 91.020 ;
        RECT 163.480 90.210 168.990 91.020 ;
        RECT 169.000 90.210 170.830 91.020 ;
        RECT 173.955 90.890 174.875 91.120 ;
        RECT 171.410 90.210 174.875 90.890 ;
        RECT 174.990 90.295 175.420 91.080 ;
        RECT 175.440 90.890 176.370 91.120 ;
        RECT 179.675 90.890 180.595 91.120 ;
        RECT 175.440 90.210 179.340 90.890 ;
        RECT 179.675 90.210 183.140 90.890 ;
        RECT 183.260 90.210 188.770 91.020 ;
        RECT 188.780 90.210 192.450 91.020 ;
        RECT 193.970 90.890 194.900 91.120 ;
        RECT 193.065 90.210 194.900 90.890 ;
        RECT 195.415 90.210 198.890 91.120 ;
        RECT 198.900 90.210 200.730 91.020 ;
        RECT 200.750 90.295 201.180 91.080 ;
        RECT 201.200 90.210 203.030 91.020 ;
        RECT 203.985 90.890 205.330 91.120 ;
        RECT 203.500 90.210 205.330 90.890 ;
        RECT 205.340 90.210 207.170 91.020 ;
        RECT 207.190 90.210 209.920 91.120 ;
        RECT 210.090 90.210 213.745 91.120 ;
        RECT 214.080 90.210 219.590 91.020 ;
        RECT 219.600 90.210 225.110 91.020 ;
        RECT 225.120 90.210 226.490 91.020 ;
        RECT 226.510 90.295 226.940 91.080 ;
        RECT 226.975 90.210 230.630 91.120 ;
        RECT 230.640 90.210 233.850 91.120 ;
        RECT 233.860 90.210 239.370 91.020 ;
        RECT 239.380 90.210 241.210 91.020 ;
        RECT 241.220 90.210 244.890 91.120 ;
        RECT 244.915 90.210 248.570 91.120 ;
        RECT 248.580 90.210 252.250 91.020 ;
        RECT 252.270 90.295 252.700 91.080 ;
        RECT 252.720 90.210 258.230 91.020 ;
        RECT 258.240 90.210 260.070 91.020 ;
        RECT 260.540 90.210 263.750 91.120 ;
        RECT 263.760 90.210 266.970 91.120 ;
        RECT 268.315 90.920 269.270 91.120 ;
        RECT 266.990 90.240 269.270 90.920 ;
        RECT 162.240 90.000 162.410 90.210 ;
        RECT 163.620 90.000 163.790 90.210 ;
        RECT 169.140 90.020 169.310 90.210 ;
        RECT 170.975 90.050 171.095 90.160 ;
        RECT 171.440 90.020 171.610 90.210 ;
        RECT 175.855 90.020 176.025 90.210 ;
        RECT 177.880 90.000 178.050 90.190 ;
        RECT 178.615 90.000 178.785 90.190 ;
        RECT 182.480 90.000 182.650 90.190 ;
        RECT 182.940 90.020 183.110 90.210 ;
        RECT 183.400 90.020 183.570 90.210 ;
        RECT 188.920 90.020 189.090 90.210 ;
        RECT 193.065 90.190 193.230 90.210 ;
        RECT 190.760 90.020 190.930 90.190 ;
        RECT 190.760 90.000 190.900 90.020 ;
        RECT 191.220 90.000 191.390 90.190 ;
        RECT 192.595 90.050 192.715 90.160 ;
        RECT 193.060 90.020 193.230 90.190 ;
        RECT 196.740 90.000 196.910 90.190 ;
        RECT 198.575 90.020 198.745 90.210 ;
        RECT 199.040 90.020 199.210 90.210 ;
        RECT 201.340 90.020 201.510 90.210 ;
        RECT 202.260 90.020 202.430 90.190 ;
        RECT 203.175 90.050 203.295 90.160 ;
        RECT 203.640 90.020 203.810 90.210 ;
        RECT 205.480 90.020 205.650 90.210 ;
        RECT 202.265 90.000 202.430 90.020 ;
        RECT 206.860 90.000 207.030 90.190 ;
        RECT 209.620 90.020 209.790 90.210 ;
        RECT 210.090 90.190 210.250 90.210 ;
        RECT 210.080 90.020 210.250 90.190 ;
        RECT 210.535 90.000 210.705 90.190 ;
        RECT 211.000 90.000 211.170 90.190 ;
        RECT 214.220 90.000 214.390 90.210 ;
        RECT 218.370 90.000 218.540 90.190 ;
        RECT 218.820 90.000 218.990 90.190 ;
        RECT 219.740 90.020 219.910 90.210 ;
        RECT 224.340 90.000 224.510 90.190 ;
        RECT 225.260 90.020 225.430 90.210 ;
        RECT 228.020 90.000 228.190 90.190 ;
        RECT 230.315 90.020 230.485 90.210 ;
        RECT 162.100 89.190 163.470 90.000 ;
        RECT 163.480 89.190 168.990 90.000 ;
        RECT 169.000 89.320 178.190 90.000 ;
        RECT 178.200 89.320 182.100 90.000 ;
        RECT 169.000 89.090 169.920 89.320 ;
        RECT 172.750 89.100 173.680 89.320 ;
        RECT 178.200 89.090 179.130 89.320 ;
        RECT 182.340 89.190 187.850 90.000 ;
        RECT 187.870 89.130 188.300 89.915 ;
        RECT 188.330 89.180 190.900 90.000 ;
        RECT 191.080 89.190 196.590 90.000 ;
        RECT 196.600 89.190 202.110 90.000 ;
        RECT 202.265 89.320 204.100 90.000 ;
        RECT 188.330 89.090 189.920 89.180 ;
        RECT 203.170 89.090 204.100 89.320 ;
        RECT 204.430 89.090 207.160 90.000 ;
        RECT 207.375 89.090 210.850 90.000 ;
        RECT 210.860 89.190 213.610 90.000 ;
        RECT 213.630 89.130 214.060 89.915 ;
        RECT 214.080 89.190 215.450 90.000 ;
        RECT 215.460 89.090 218.670 90.000 ;
        RECT 218.680 89.190 224.190 90.000 ;
        RECT 224.200 89.190 227.870 90.000 ;
        RECT 227.880 89.190 229.250 90.000 ;
        RECT 229.260 89.970 230.215 90.000 ;
        RECT 231.245 89.970 231.415 90.190 ;
        RECT 231.700 90.000 231.870 90.190 ;
        RECT 233.540 90.020 233.710 90.210 ;
        RECT 234.000 90.020 234.170 90.210 ;
        RECT 237.220 90.000 237.390 90.190 ;
        RECT 239.055 90.050 239.175 90.160 ;
        RECT 239.520 90.020 239.690 90.210 ;
        RECT 239.980 90.000 240.150 90.190 ;
        RECT 241.365 90.020 241.535 90.210 ;
        RECT 242.730 90.000 242.900 90.190 ;
        RECT 245.960 90.000 246.130 90.190 ;
        RECT 248.255 90.020 248.425 90.210 ;
        RECT 248.720 90.020 248.890 90.210 ;
        RECT 251.480 90.000 251.650 90.190 ;
        RECT 252.860 90.020 253.030 90.210 ;
        RECT 257.000 90.000 257.170 90.190 ;
        RECT 258.380 90.020 258.550 90.210 ;
        RECT 260.225 90.160 260.395 90.190 ;
        RECT 259.755 90.050 259.875 90.160 ;
        RECT 260.215 90.050 260.395 90.160 ;
        RECT 260.225 90.000 260.395 90.050 ;
        RECT 260.680 90.020 260.850 90.210 ;
        RECT 263.900 90.000 264.070 90.210 ;
        RECT 267.115 90.020 267.285 90.240 ;
        RECT 268.315 90.210 269.270 90.240 ;
        RECT 269.280 90.210 274.790 91.020 ;
        RECT 274.800 90.210 277.550 91.020 ;
        RECT 278.030 90.295 278.460 91.080 ;
        RECT 278.480 90.210 282.150 91.120 ;
        RECT 282.160 90.210 284.910 91.120 ;
        RECT 284.920 90.210 288.590 91.020 ;
        RECT 288.600 90.210 289.970 91.020 ;
        RECT 289.980 90.890 290.910 91.120 ;
        RECT 299.090 90.890 300.020 91.110 ;
        RECT 302.850 90.890 303.770 91.120 ;
        RECT 289.980 90.210 293.880 90.890 ;
        RECT 294.580 90.210 303.770 90.890 ;
        RECT 303.790 90.295 304.220 91.080 ;
        RECT 304.240 90.210 307.910 91.020 ;
        RECT 308.405 90.890 309.750 91.120 ;
        RECT 307.920 90.210 309.750 90.890 ;
        RECT 309.760 90.210 311.130 91.020 ;
        RECT 269.420 90.020 269.590 90.210 ;
        RECT 270.340 90.000 270.510 90.190 ;
        RECT 270.800 90.000 270.970 90.190 ;
        RECT 274.490 90.045 274.650 90.155 ;
        RECT 274.940 90.020 275.110 90.210 ;
        RECT 229.260 89.290 231.540 89.970 ;
        RECT 229.260 89.090 230.215 89.290 ;
        RECT 231.560 89.190 237.070 90.000 ;
        RECT 237.080 89.190 238.910 90.000 ;
        RECT 239.390 89.130 239.820 89.915 ;
        RECT 239.840 89.190 242.590 90.000 ;
        RECT 242.600 89.090 245.810 90.000 ;
        RECT 245.820 89.190 251.330 90.000 ;
        RECT 251.340 89.190 256.850 90.000 ;
        RECT 256.860 89.190 259.610 90.000 ;
        RECT 260.080 89.090 263.735 90.000 ;
        RECT 263.760 89.190 265.130 90.000 ;
        RECT 265.150 89.130 265.580 89.915 ;
        RECT 265.835 89.320 270.650 90.000 ;
        RECT 270.660 89.190 274.330 90.000 ;
        RECT 275.405 89.970 275.575 90.190 ;
        RECT 277.695 90.050 277.815 90.160 ;
        RECT 278.625 90.020 278.795 90.210 ;
        RECT 282.760 90.000 282.930 90.190 ;
        RECT 283.220 90.000 283.390 90.190 ;
        RECT 284.600 90.020 284.770 90.210 ;
        RECT 285.060 90.020 285.230 90.210 ;
        RECT 288.740 90.020 288.910 90.210 ;
        RECT 290.395 90.190 290.565 90.210 ;
        RECT 290.305 90.020 290.565 90.190 ;
        RECT 290.305 90.000 290.475 90.020 ;
        RECT 291.500 90.000 291.670 90.190 ;
        RECT 294.255 90.050 294.375 90.160 ;
        RECT 294.720 90.020 294.890 90.210 ;
        RECT 295.180 90.000 295.350 90.190 ;
        RECT 304.380 90.020 304.550 90.210 ;
        RECT 304.840 90.000 305.010 90.190 ;
        RECT 307.600 90.000 307.770 90.190 ;
        RECT 308.060 90.020 308.230 90.210 ;
        RECT 309.435 90.050 309.555 90.160 ;
        RECT 310.820 90.000 310.990 90.210 ;
        RECT 277.065 89.970 278.010 90.000 ;
        RECT 275.260 89.290 278.010 89.970 ;
        RECT 278.255 89.320 283.070 90.000 ;
        RECT 277.065 89.090 278.010 89.290 ;
        RECT 283.080 89.190 286.750 90.000 ;
        RECT 286.990 89.320 290.890 90.000 ;
        RECT 289.960 89.090 290.890 89.320 ;
        RECT 290.910 89.130 291.340 89.915 ;
        RECT 291.360 89.190 295.030 90.000 ;
        RECT 295.040 89.320 304.650 90.000 ;
        RECT 304.700 89.320 307.440 90.000 ;
        RECT 299.550 89.100 300.480 89.320 ;
        RECT 303.310 89.090 304.650 89.320 ;
        RECT 307.460 89.190 309.290 90.000 ;
        RECT 309.760 89.190 311.130 90.000 ;
      LAYER nwell ;
        RECT 161.905 85.970 311.325 88.800 ;
      LAYER pwell ;
        RECT 162.100 84.770 163.470 85.580 ;
        RECT 163.480 84.770 165.310 85.580 ;
        RECT 165.780 85.450 166.700 85.680 ;
        RECT 169.530 85.450 170.460 85.670 ;
        RECT 165.780 84.770 174.970 85.450 ;
        RECT 174.990 84.855 175.420 85.640 ;
        RECT 175.440 85.450 176.370 85.680 ;
        RECT 179.580 85.450 180.510 85.680 ;
        RECT 185.570 85.590 187.160 85.680 ;
        RECT 188.330 85.590 189.920 85.680 ;
        RECT 175.440 84.770 179.340 85.450 ;
        RECT 179.580 84.770 183.480 85.450 ;
        RECT 183.720 84.770 185.550 85.580 ;
        RECT 185.570 84.770 188.140 85.590 ;
        RECT 188.330 84.770 190.900 85.590 ;
        RECT 191.080 84.770 192.910 85.580 ;
        RECT 193.690 85.450 194.620 85.680 ;
        RECT 193.690 84.770 195.525 85.450 ;
        RECT 195.875 84.770 199.350 85.680 ;
        RECT 199.360 84.770 200.730 85.580 ;
        RECT 200.750 84.855 201.180 85.640 ;
        RECT 203.170 85.450 204.100 85.680 ;
        RECT 202.265 84.770 204.100 85.450 ;
        RECT 205.535 84.770 209.010 85.680 ;
        RECT 209.020 84.770 210.390 85.580 ;
        RECT 211.450 85.450 212.380 85.680 ;
        RECT 210.545 84.770 212.380 85.450 ;
        RECT 212.700 84.770 218.210 85.580 ;
        RECT 218.220 84.770 223.730 85.580 ;
        RECT 223.740 84.770 226.490 85.580 ;
        RECT 226.510 84.855 226.940 85.640 ;
        RECT 226.960 84.770 232.470 85.580 ;
        RECT 232.480 84.770 237.990 85.580 ;
        RECT 238.000 84.770 241.670 85.580 ;
        RECT 242.140 85.450 243.485 85.680 ;
        RECT 242.140 84.770 243.970 85.450 ;
        RECT 244.060 84.770 246.270 85.680 ;
        RECT 249.940 85.450 250.870 85.680 ;
        RECT 247.200 84.770 250.870 85.450 ;
        RECT 250.880 84.770 252.250 85.580 ;
        RECT 252.270 84.855 252.700 85.640 ;
        RECT 252.720 84.770 258.230 85.580 ;
        RECT 258.240 84.770 263.750 85.580 ;
        RECT 264.220 84.770 267.380 85.680 ;
        RECT 267.440 84.770 272.950 85.580 ;
        RECT 272.960 84.770 276.630 85.580 ;
        RECT 276.640 84.770 278.010 85.580 ;
        RECT 278.030 84.855 278.460 85.640 ;
        RECT 278.480 84.770 280.570 85.580 ;
        RECT 281.710 84.770 284.440 85.680 ;
        RECT 284.460 84.770 288.130 85.580 ;
        RECT 293.110 85.450 294.040 85.670 ;
        RECT 296.870 85.450 297.790 85.680 ;
        RECT 288.600 84.770 297.790 85.450 ;
        RECT 297.800 85.450 298.730 85.680 ;
        RECT 297.800 84.770 301.700 85.450 ;
        RECT 301.940 84.770 303.770 85.580 ;
        RECT 303.790 84.855 304.220 85.640 ;
        RECT 304.240 85.450 305.170 85.680 ;
        RECT 304.240 84.770 308.140 85.450 ;
        RECT 308.380 84.770 309.750 85.550 ;
        RECT 309.760 84.770 311.130 85.580 ;
        RECT 162.240 84.560 162.410 84.770 ;
        RECT 163.620 84.560 163.790 84.770 ;
        RECT 165.455 84.610 165.575 84.720 ;
        RECT 169.140 84.560 169.310 84.750 ;
        RECT 174.660 84.580 174.830 84.770 ;
        RECT 175.855 84.580 176.025 84.770 ;
        RECT 179.720 84.560 179.890 84.750 ;
        RECT 179.995 84.580 180.165 84.770 ;
        RECT 180.180 84.560 180.350 84.750 ;
        RECT 182.935 84.610 183.055 84.720 ;
        RECT 183.400 84.560 183.570 84.750 ;
        RECT 183.860 84.580 184.030 84.770 ;
        RECT 188.000 84.750 188.140 84.770 ;
        RECT 190.760 84.750 190.900 84.770 ;
        RECT 186.160 84.560 186.330 84.750 ;
        RECT 188.000 84.580 188.170 84.750 ;
        RECT 190.760 84.580 190.930 84.750 ;
        RECT 190.760 84.560 190.900 84.580 ;
        RECT 191.220 84.560 191.390 84.770 ;
        RECT 195.360 84.750 195.525 84.770 ;
        RECT 193.055 84.610 193.175 84.720 ;
        RECT 195.360 84.580 195.530 84.750 ;
        RECT 196.740 84.560 196.910 84.750 ;
        RECT 199.035 84.580 199.205 84.770 ;
        RECT 199.500 84.580 199.670 84.770 ;
        RECT 202.265 84.750 202.430 84.770 ;
        RECT 201.350 84.615 201.510 84.725 ;
        RECT 202.260 84.560 202.430 84.750 ;
        RECT 204.570 84.615 204.730 84.725 ;
        RECT 205.950 84.605 206.110 84.715 ;
        RECT 206.860 84.560 207.030 84.750 ;
        RECT 208.695 84.580 208.865 84.770 ;
        RECT 209.160 84.580 209.330 84.770 ;
        RECT 210.545 84.750 210.710 84.770 ;
        RECT 209.615 84.610 209.735 84.720 ;
        RECT 210.540 84.580 210.710 84.750 ;
        RECT 212.840 84.580 213.010 84.770 ;
        RECT 213.295 84.560 213.465 84.750 ;
        RECT 214.225 84.560 214.395 84.750 ;
        RECT 217.900 84.560 218.070 84.750 ;
        RECT 218.360 84.580 218.530 84.770 ;
        RECT 223.420 84.560 223.590 84.750 ;
        RECT 223.880 84.580 224.050 84.770 ;
        RECT 227.100 84.560 227.270 84.770 ;
        RECT 230.320 84.560 230.490 84.750 ;
        RECT 232.620 84.580 232.790 84.770 ;
        RECT 235.840 84.560 236.010 84.750 ;
        RECT 238.140 84.580 238.310 84.770 ;
        RECT 239.990 84.605 240.150 84.715 ;
        RECT 241.815 84.610 241.935 84.720 ;
        RECT 242.275 84.560 242.445 84.750 ;
        RECT 243.660 84.580 243.830 84.770 ;
        RECT 245.955 84.560 246.125 84.770 ;
        RECT 246.430 84.615 246.590 84.725 ;
        RECT 247.340 84.580 247.510 84.770 ;
        RECT 162.100 83.750 163.470 84.560 ;
        RECT 163.480 83.750 168.990 84.560 ;
        RECT 169.000 83.750 170.830 84.560 ;
        RECT 170.840 83.880 180.030 84.560 ;
        RECT 170.840 83.650 171.760 83.880 ;
        RECT 174.590 83.660 175.520 83.880 ;
        RECT 180.040 83.750 182.790 84.560 ;
        RECT 183.260 83.650 186.010 84.560 ;
        RECT 186.020 83.750 187.850 84.560 ;
        RECT 187.870 83.690 188.300 84.475 ;
        RECT 188.330 83.740 190.900 84.560 ;
        RECT 191.080 83.750 196.590 84.560 ;
        RECT 196.600 83.750 202.110 84.560 ;
        RECT 202.120 83.750 205.790 84.560 ;
        RECT 206.720 83.750 208.810 84.560 ;
        RECT 188.330 83.650 189.920 83.740 ;
        RECT 210.135 83.650 213.610 84.560 ;
        RECT 213.630 83.690 214.060 84.475 ;
        RECT 214.080 83.650 217.555 84.560 ;
        RECT 217.760 83.750 223.270 84.560 ;
        RECT 223.280 83.750 226.950 84.560 ;
        RECT 226.960 83.650 230.170 84.560 ;
        RECT 230.180 83.750 235.690 84.560 ;
        RECT 235.700 83.750 239.370 84.560 ;
        RECT 239.390 83.690 239.820 84.475 ;
        RECT 240.820 83.650 242.590 84.560 ;
        RECT 242.615 83.650 246.270 84.560 ;
        RECT 246.280 84.530 247.650 84.560 ;
        RECT 249.640 84.530 249.810 84.750 ;
        RECT 250.100 84.560 250.270 84.750 ;
        RECT 251.020 84.580 251.190 84.770 ;
        RECT 252.860 84.580 253.030 84.770 ;
        RECT 253.320 84.560 253.490 84.750 ;
        RECT 253.780 84.560 253.950 84.750 ;
        RECT 257.460 84.560 257.630 84.750 ;
        RECT 258.380 84.580 258.550 84.770 ;
        RECT 258.840 84.560 259.010 84.750 ;
        RECT 246.280 83.850 249.950 84.530 ;
        RECT 249.960 83.880 251.790 84.560 ;
        RECT 251.800 83.880 253.630 84.560 ;
        RECT 246.280 83.650 247.665 83.850 ;
        RECT 250.445 83.650 251.790 83.880 ;
        RECT 253.640 83.750 257.310 84.560 ;
        RECT 257.320 83.750 258.690 84.560 ;
        RECT 258.700 83.650 261.910 84.560 ;
        RECT 262.065 84.530 262.235 84.750 ;
        RECT 263.895 84.610 264.015 84.720 ;
        RECT 264.815 84.610 264.935 84.720 ;
        RECT 267.120 84.580 267.290 84.770 ;
        RECT 267.580 84.580 267.750 84.770 ;
        RECT 267.580 84.560 267.730 84.580 ;
        RECT 268.040 84.560 268.210 84.750 ;
        RECT 273.100 84.580 273.270 84.770 ;
        RECT 273.560 84.560 273.730 84.750 ;
        RECT 276.780 84.580 276.950 84.770 ;
        RECT 278.620 84.580 278.790 84.770 ;
        RECT 279.080 84.560 279.250 84.750 ;
        RECT 281.375 84.610 281.495 84.720 ;
        RECT 281.840 84.580 282.010 84.770 ;
        RECT 284.600 84.560 284.770 84.770 ;
        RECT 287.355 84.610 287.475 84.720 ;
        RECT 287.820 84.560 287.990 84.750 ;
        RECT 288.275 84.610 288.395 84.720 ;
        RECT 288.740 84.580 288.910 84.770 ;
        RECT 290.575 84.610 290.695 84.720 ;
        RECT 291.500 84.560 291.670 84.750 ;
        RECT 294.255 84.610 294.375 84.720 ;
        RECT 294.720 84.560 294.890 84.750 ;
        RECT 298.215 84.580 298.385 84.770 ;
        RECT 302.080 84.580 302.250 84.770 ;
        RECT 304.195 84.560 304.365 84.750 ;
        RECT 304.655 84.580 304.825 84.770 ;
        RECT 308.060 84.560 308.230 84.750 ;
        RECT 309.440 84.580 309.610 84.770 ;
        RECT 310.820 84.560 310.990 84.770 ;
        RECT 263.725 84.530 264.670 84.560 ;
        RECT 261.920 83.850 264.670 84.530 ;
        RECT 263.725 83.650 264.670 83.850 ;
        RECT 265.150 83.690 265.580 84.475 ;
        RECT 265.800 83.740 267.730 84.560 ;
        RECT 267.900 83.750 273.410 84.560 ;
        RECT 273.420 83.750 278.930 84.560 ;
        RECT 278.940 83.750 284.450 84.560 ;
        RECT 284.460 83.750 287.210 84.560 ;
        RECT 287.680 83.750 289.770 84.560 ;
        RECT 265.800 83.650 266.750 83.740 ;
        RECT 290.910 83.690 291.340 84.475 ;
        RECT 291.360 83.750 294.110 84.560 ;
        RECT 294.580 83.880 303.770 84.560 ;
        RECT 299.090 83.660 300.020 83.880 ;
        RECT 302.850 83.650 303.770 83.880 ;
        RECT 303.780 83.880 307.680 84.560 ;
        RECT 303.780 83.650 304.710 83.880 ;
        RECT 307.920 83.750 309.750 84.560 ;
        RECT 309.760 83.750 311.130 84.560 ;
      LAYER nwell ;
        RECT 161.905 80.530 311.325 83.360 ;
      LAYER pwell ;
        RECT 162.100 79.330 163.470 80.140 ;
        RECT 163.480 79.330 165.310 80.140 ;
        RECT 165.780 80.010 166.700 80.240 ;
        RECT 169.530 80.010 170.460 80.230 ;
        RECT 165.780 79.330 174.970 80.010 ;
        RECT 174.990 79.415 175.420 80.200 ;
        RECT 175.440 79.330 179.110 80.140 ;
        RECT 179.120 79.330 180.490 80.140 ;
        RECT 180.500 80.010 181.430 80.240 ;
        RECT 180.500 79.330 184.400 80.010 ;
        RECT 184.640 79.330 190.150 80.140 ;
        RECT 190.160 79.330 191.990 80.140 ;
        RECT 193.800 80.040 195.180 80.240 ;
        RECT 192.475 79.360 195.180 80.040 ;
        RECT 162.240 79.120 162.410 79.330 ;
        RECT 163.620 79.120 163.790 79.330 ;
        RECT 165.455 79.170 165.575 79.280 ;
        RECT 169.140 79.120 169.310 79.310 ;
        RECT 173.095 79.120 173.265 79.310 ;
        RECT 174.660 79.140 174.830 79.330 ;
        RECT 175.580 79.140 175.750 79.330 ;
        RECT 176.960 79.120 177.130 79.310 ;
        RECT 179.260 79.140 179.430 79.330 ;
        RECT 180.915 79.140 181.085 79.330 ;
        RECT 184.780 79.140 184.950 79.330 ;
        RECT 186.620 79.120 186.790 79.310 ;
        RECT 188.460 79.120 188.630 79.310 ;
        RECT 190.300 79.140 190.470 79.330 ;
        RECT 191.215 79.170 191.335 79.280 ;
        RECT 191.680 79.140 191.850 79.310 ;
        RECT 192.135 79.170 192.255 79.280 ;
        RECT 192.600 79.140 192.770 79.360 ;
        RECT 193.800 79.330 195.180 79.360 ;
        RECT 195.220 79.330 197.970 80.240 ;
        RECT 197.980 79.330 200.730 80.140 ;
        RECT 200.750 79.415 201.180 80.200 ;
        RECT 201.200 79.330 203.030 80.010 ;
        RECT 203.960 79.330 210.470 80.240 ;
        RECT 211.240 79.330 217.750 80.240 ;
        RECT 217.760 79.330 223.270 80.140 ;
        RECT 225.080 80.040 226.490 80.240 ;
        RECT 223.755 79.360 226.490 80.040 ;
        RECT 226.510 79.415 226.940 80.200 ;
        RECT 197.660 79.140 197.830 79.330 ;
        RECT 198.120 79.120 198.290 79.330 ;
        RECT 201.340 79.140 201.510 79.330 ;
        RECT 201.795 79.120 201.965 79.310 ;
        RECT 202.270 79.165 202.430 79.275 ;
        RECT 162.100 78.310 163.470 79.120 ;
        RECT 163.480 78.310 168.990 79.120 ;
        RECT 169.000 78.310 172.670 79.120 ;
        RECT 172.680 78.440 176.580 79.120 ;
        RECT 176.820 78.440 186.430 79.120 ;
        RECT 172.680 78.210 173.610 78.440 ;
        RECT 181.330 78.220 182.260 78.440 ;
        RECT 185.090 78.210 186.430 78.440 ;
        RECT 186.480 78.310 187.850 79.120 ;
        RECT 187.870 78.250 188.300 79.035 ;
        RECT 188.320 78.310 190.410 79.120 ;
        RECT 192.005 78.440 193.370 79.120 ;
        RECT 193.615 78.440 198.430 79.120 ;
        RECT 198.635 78.210 202.110 79.120 ;
        RECT 203.180 79.090 203.350 79.310 ;
        RECT 204.105 79.140 204.275 79.330 ;
        RECT 206.860 79.120 207.030 79.310 ;
        RECT 211.920 79.120 212.090 79.310 ;
        RECT 214.230 79.165 214.390 79.275 ;
        RECT 215.415 79.120 215.585 79.310 ;
        RECT 217.435 79.140 217.605 79.330 ;
        RECT 217.900 79.140 218.070 79.330 ;
        RECT 219.280 79.140 219.450 79.310 ;
        RECT 219.285 79.120 219.450 79.140 ;
        RECT 221.580 79.120 221.750 79.310 ;
        RECT 223.415 79.170 223.535 79.280 ;
        RECT 223.880 79.120 224.050 79.360 ;
        RECT 225.095 79.330 226.490 79.360 ;
        RECT 226.960 79.330 228.330 80.140 ;
        RECT 228.355 79.330 232.010 80.240 ;
        RECT 232.030 79.330 234.760 80.240 ;
        RECT 234.780 79.330 238.450 80.140 ;
        RECT 238.920 79.330 242.130 80.240 ;
        RECT 242.155 79.330 245.810 80.240 ;
        RECT 245.820 79.330 249.030 80.240 ;
        RECT 249.240 80.150 250.190 80.240 ;
        RECT 249.240 79.330 251.170 80.150 ;
        RECT 252.270 79.415 252.700 80.200 ;
        RECT 252.720 79.330 256.390 80.140 ;
        RECT 256.400 79.330 260.055 80.240 ;
        RECT 260.080 79.330 263.735 80.240 ;
        RECT 263.760 79.330 266.970 80.240 ;
        RECT 268.785 80.040 269.730 80.240 ;
        RECT 276.410 80.150 278.000 80.240 ;
        RECT 266.980 79.360 269.730 80.040 ;
        RECT 205.340 79.090 206.710 79.120 ;
        RECT 203.040 78.410 206.710 79.090 ;
        RECT 206.720 78.440 211.535 79.120 ;
        RECT 205.325 78.210 206.710 78.410 ;
        RECT 211.780 78.310 213.610 79.120 ;
        RECT 213.630 78.250 214.060 79.035 ;
        RECT 215.000 78.440 218.900 79.120 ;
        RECT 219.285 78.440 221.120 79.120 ;
        RECT 215.000 78.210 215.930 78.440 ;
        RECT 220.190 78.210 221.120 78.440 ;
        RECT 221.440 78.310 223.270 79.120 ;
        RECT 223.740 78.210 226.490 79.120 ;
        RECT 226.640 79.090 226.810 79.310 ;
        RECT 227.100 79.140 227.270 79.330 ;
        RECT 230.320 79.120 230.490 79.310 ;
        RECT 231.695 79.140 231.865 79.330 ;
        RECT 232.160 79.140 232.330 79.330 ;
        RECT 234.920 79.140 235.090 79.330 ;
        RECT 235.840 79.120 236.010 79.310 ;
        RECT 238.595 79.170 238.715 79.280 ;
        RECT 239.060 79.140 239.230 79.330 ;
        RECT 239.980 79.120 240.150 79.310 ;
        RECT 242.735 79.170 242.855 79.280 ;
        RECT 228.800 79.090 230.170 79.120 ;
        RECT 226.500 78.410 230.170 79.090 ;
        RECT 228.785 78.210 230.170 78.410 ;
        RECT 230.180 78.310 235.690 79.120 ;
        RECT 235.700 78.310 239.370 79.120 ;
        RECT 239.390 78.250 239.820 79.035 ;
        RECT 239.840 78.310 242.590 79.120 ;
        RECT 243.205 79.090 243.375 79.310 ;
        RECT 245.495 79.140 245.665 79.330 ;
        RECT 245.960 79.120 246.130 79.310 ;
        RECT 248.720 79.140 248.890 79.330 ;
        RECT 251.020 79.310 251.170 79.330 ;
        RECT 251.020 79.140 251.190 79.310 ;
        RECT 251.480 79.120 251.650 79.310 ;
        RECT 252.860 79.140 253.030 79.330 ;
        RECT 256.545 79.140 256.715 79.330 ;
        RECT 256.995 79.170 257.115 79.280 ;
        RECT 257.460 79.120 257.630 79.310 ;
        RECT 260.225 79.140 260.395 79.330 ;
        RECT 260.680 79.120 260.850 79.310 ;
        RECT 263.900 79.120 264.070 79.330 ;
        RECT 265.740 79.140 265.910 79.310 ;
        RECT 267.125 79.140 267.295 79.360 ;
        RECT 268.785 79.330 269.730 79.360 ;
        RECT 269.740 79.330 275.250 80.140 ;
        RECT 275.430 79.330 278.000 80.150 ;
        RECT 278.030 79.415 278.460 80.200 ;
        RECT 278.480 79.330 280.310 80.140 ;
        RECT 280.320 80.010 281.250 80.240 ;
        RECT 280.320 79.330 284.220 80.010 ;
        RECT 284.460 79.330 287.210 80.140 ;
        RECT 287.680 79.330 292.495 80.010 ;
        RECT 292.740 79.330 294.110 80.140 ;
        RECT 298.630 80.010 299.560 80.230 ;
        RECT 302.390 80.010 303.310 80.240 ;
        RECT 294.120 79.330 303.310 80.010 ;
        RECT 303.790 79.415 304.220 80.200 ;
        RECT 304.240 79.330 309.750 80.140 ;
        RECT 309.760 79.330 311.130 80.140 ;
        RECT 265.760 79.120 265.910 79.140 ;
        RECT 268.040 79.120 268.210 79.310 ;
        RECT 269.880 79.140 270.050 79.330 ;
        RECT 275.430 79.310 275.570 79.330 ;
        RECT 273.560 79.120 273.730 79.310 ;
        RECT 275.400 79.140 275.570 79.310 ;
        RECT 276.315 79.170 276.435 79.280 ;
        RECT 276.780 79.120 276.950 79.310 ;
        RECT 278.620 79.140 278.790 79.330 ;
        RECT 280.735 79.140 280.905 79.330 ;
        RECT 284.600 79.140 284.770 79.330 ;
        RECT 285.980 79.120 286.150 79.310 ;
        RECT 287.355 79.170 287.475 79.280 ;
        RECT 287.820 79.140 287.990 79.330 ;
        RECT 291.505 79.120 291.675 79.310 ;
        RECT 292.880 79.140 293.050 79.330 ;
        RECT 294.260 79.140 294.430 79.330 ;
        RECT 302.540 79.120 302.710 79.310 ;
        RECT 303.455 79.170 303.575 79.280 ;
        RECT 304.380 79.140 304.550 79.330 ;
        RECT 308.060 79.120 308.230 79.310 ;
        RECT 310.820 79.120 310.990 79.330 ;
        RECT 244.865 79.090 245.810 79.120 ;
        RECT 243.060 78.410 245.810 79.090 ;
        RECT 244.865 78.210 245.810 78.410 ;
        RECT 245.820 78.310 251.330 79.120 ;
        RECT 251.340 78.310 256.850 79.120 ;
        RECT 257.320 78.210 260.530 79.120 ;
        RECT 260.540 78.210 263.750 79.120 ;
        RECT 263.760 78.310 265.130 79.120 ;
        RECT 265.150 78.250 265.580 79.035 ;
        RECT 265.760 78.300 267.690 79.120 ;
        RECT 267.900 78.310 273.410 79.120 ;
        RECT 273.420 78.310 276.170 79.120 ;
        RECT 276.640 78.440 285.830 79.120 ;
        RECT 285.840 78.440 290.655 79.120 ;
        RECT 266.740 78.210 267.690 78.300 ;
        RECT 281.150 78.220 282.080 78.440 ;
        RECT 284.910 78.210 285.830 78.440 ;
        RECT 290.910 78.250 291.340 79.035 ;
        RECT 291.360 78.210 302.370 79.120 ;
        RECT 302.400 78.310 307.910 79.120 ;
        RECT 307.920 78.310 309.750 79.120 ;
        RECT 309.760 78.310 311.130 79.120 ;
      LAYER nwell ;
        RECT 161.905 75.090 311.325 77.920 ;
      LAYER pwell ;
        RECT 162.100 73.890 163.470 74.700 ;
        RECT 163.480 73.890 165.310 74.700 ;
        RECT 170.290 74.570 171.220 74.790 ;
        RECT 174.050 74.570 174.970 74.800 ;
        RECT 165.780 73.890 174.970 74.570 ;
        RECT 174.990 73.975 175.420 74.760 ;
        RECT 175.440 73.890 179.110 74.700 ;
        RECT 183.630 74.570 184.560 74.790 ;
        RECT 187.390 74.570 188.310 74.800 ;
        RECT 179.120 73.890 188.310 74.570 ;
        RECT 188.320 73.890 191.520 74.800 ;
        RECT 191.540 74.570 192.460 74.800 ;
        RECT 195.290 74.570 196.220 74.790 ;
        RECT 191.540 73.890 200.730 74.570 ;
        RECT 200.750 73.975 201.180 74.760 ;
        RECT 201.200 74.570 202.130 74.800 ;
        RECT 201.200 73.890 205.100 74.570 ;
        RECT 205.350 73.890 208.090 74.570 ;
        RECT 208.100 73.890 209.930 74.700 ;
        RECT 213.600 74.570 214.530 74.800 ;
        RECT 219.050 74.570 219.980 74.790 ;
        RECT 222.810 74.570 223.730 74.800 ;
        RECT 210.630 73.890 214.530 74.570 ;
        RECT 214.540 73.890 223.730 74.570 ;
        RECT 223.740 74.570 225.085 74.800 ;
        RECT 223.740 73.890 225.570 74.570 ;
        RECT 226.510 73.975 226.940 74.760 ;
        RECT 226.960 73.890 232.470 74.700 ;
        RECT 232.480 73.890 236.150 74.700 ;
        RECT 236.160 74.600 237.115 74.800 ;
        RECT 236.160 73.920 238.440 74.600 ;
        RECT 236.160 73.890 237.115 73.920 ;
        RECT 162.240 73.680 162.410 73.890 ;
        RECT 163.620 73.680 163.790 73.890 ;
        RECT 165.455 73.730 165.575 73.840 ;
        RECT 165.920 73.700 166.090 73.890 ;
        RECT 167.310 73.725 167.470 73.835 ;
        RECT 175.580 73.700 175.750 73.890 ;
        RECT 177.420 73.680 177.590 73.870 ;
        RECT 178.155 73.680 178.325 73.870 ;
        RECT 179.260 73.700 179.430 73.890 ;
        RECT 182.030 73.725 182.190 73.835 ;
        RECT 183.215 73.680 183.385 73.870 ;
        RECT 187.090 73.725 187.250 73.835 ;
        RECT 188.460 73.680 188.630 73.870 ;
        RECT 191.225 73.700 191.395 73.890 ;
        RECT 193.520 73.680 193.690 73.870 ;
        RECT 196.735 73.730 196.855 73.840 ;
        RECT 197.200 73.680 197.370 73.870 ;
        RECT 200.420 73.700 200.590 73.890 ;
        RECT 201.615 73.700 201.785 73.890 ;
        RECT 207.780 73.700 207.950 73.890 ;
        RECT 208.240 73.700 208.410 73.890 ;
        RECT 209.165 73.680 209.335 73.870 ;
        RECT 209.620 73.680 209.790 73.870 ;
        RECT 210.075 73.730 210.195 73.840 ;
        RECT 213.295 73.730 213.415 73.840 ;
        RECT 213.945 73.700 214.115 73.890 ;
        RECT 214.220 73.680 214.390 73.870 ;
        RECT 214.680 73.700 214.850 73.890 ;
        RECT 223.420 73.680 223.590 73.870 ;
        RECT 225.260 73.700 225.430 73.890 ;
        RECT 225.730 73.735 225.890 73.845 ;
        RECT 227.100 73.700 227.270 73.890 ;
        RECT 228.950 73.725 229.110 73.835 ;
        RECT 229.860 73.680 230.030 73.870 ;
        RECT 232.620 73.700 232.790 73.890 ;
        RECT 233.080 73.680 233.250 73.870 ;
        RECT 235.845 73.680 236.015 73.870 ;
        RECT 238.145 73.700 238.315 73.920 ;
        RECT 238.460 73.890 243.970 74.700 ;
        RECT 243.980 73.890 249.490 74.700 ;
        RECT 249.500 73.890 252.250 74.700 ;
        RECT 252.270 73.975 252.700 74.760 ;
        RECT 252.720 73.890 256.390 74.700 ;
        RECT 256.400 73.890 257.770 74.700 ;
        RECT 257.780 73.890 261.435 74.800 ;
        RECT 261.460 73.890 264.670 74.800 ;
        RECT 264.680 73.890 270.190 74.700 ;
        RECT 270.200 73.890 273.870 74.700 ;
        RECT 277.080 74.570 278.010 74.800 ;
        RECT 274.110 73.890 278.010 74.570 ;
        RECT 278.030 73.975 278.460 74.760 ;
        RECT 283.450 74.570 284.380 74.790 ;
        RECT 287.210 74.570 288.130 74.800 ;
        RECT 278.940 73.890 288.130 74.570 ;
        RECT 288.140 73.890 289.970 74.700 ;
        RECT 293.640 74.570 294.570 74.800 ;
        RECT 290.670 73.890 294.570 74.570 ;
        RECT 294.580 74.570 295.500 74.800 ;
        RECT 298.330 74.570 299.260 74.790 ;
        RECT 294.580 73.890 303.770 74.570 ;
        RECT 303.790 73.975 304.220 74.760 ;
        RECT 304.240 73.890 309.750 74.700 ;
        RECT 309.760 73.890 311.130 74.700 ;
        RECT 238.600 73.700 238.770 73.890 ;
        RECT 239.980 73.680 240.150 73.870 ;
        RECT 244.120 73.700 244.290 73.890 ;
        RECT 244.575 73.680 244.745 73.870 ;
        RECT 245.040 73.680 245.210 73.870 ;
        RECT 249.640 73.700 249.810 73.890 ;
        RECT 250.560 73.680 250.730 73.870 ;
        RECT 252.860 73.700 253.030 73.890 ;
        RECT 256.080 73.680 256.250 73.870 ;
        RECT 256.540 73.700 256.710 73.890 ;
        RECT 257.925 73.840 258.095 73.890 ;
        RECT 257.915 73.730 258.095 73.840 ;
        RECT 257.925 73.700 258.095 73.730 ;
        RECT 258.380 73.680 258.550 73.870 ;
        RECT 261.600 73.700 261.770 73.890 ;
        RECT 264.360 73.680 264.530 73.870 ;
        RECT 264.820 73.840 264.990 73.890 ;
        RECT 264.815 73.730 264.990 73.840 ;
        RECT 264.820 73.700 264.990 73.730 ;
        RECT 265.740 73.680 265.910 73.870 ;
        RECT 270.340 73.700 270.510 73.890 ;
        RECT 271.260 73.680 271.430 73.870 ;
        RECT 274.015 73.730 274.135 73.840 ;
        RECT 274.475 73.680 274.645 73.870 ;
        RECT 277.425 73.700 277.595 73.890 ;
        RECT 278.615 73.730 278.735 73.840 ;
        RECT 279.080 73.700 279.250 73.890 ;
        RECT 286.440 73.680 286.610 73.870 ;
        RECT 287.175 73.680 287.345 73.870 ;
        RECT 288.280 73.700 288.450 73.890 ;
        RECT 290.115 73.730 290.235 73.840 ;
        RECT 291.500 73.680 291.670 73.870 ;
        RECT 293.985 73.700 294.155 73.890 ;
        RECT 297.020 73.680 297.190 73.870 ;
        RECT 303.460 73.700 303.630 73.890 ;
        RECT 304.380 73.700 304.550 73.890 ;
        RECT 306.675 73.730 306.795 73.840 ;
        RECT 307.140 73.680 307.310 73.870 ;
        RECT 308.990 73.725 309.150 73.835 ;
        RECT 310.820 73.680 310.990 73.890 ;
        RECT 162.100 72.870 163.470 73.680 ;
        RECT 163.480 72.870 167.150 73.680 ;
        RECT 168.120 73.000 177.730 73.680 ;
        RECT 177.740 73.000 181.640 73.680 ;
        RECT 182.800 73.000 186.700 73.680 ;
        RECT 168.120 72.770 169.460 73.000 ;
        RECT 172.290 72.780 173.220 73.000 ;
        RECT 177.740 72.770 178.670 73.000 ;
        RECT 182.800 72.770 183.730 73.000 ;
        RECT 187.870 72.810 188.300 73.595 ;
        RECT 188.320 73.000 193.135 73.680 ;
        RECT 193.430 72.770 196.590 73.680 ;
        RECT 197.060 73.000 206.250 73.680 ;
        RECT 201.570 72.780 202.500 73.000 ;
        RECT 205.330 72.770 206.250 73.000 ;
        RECT 206.260 72.770 209.460 73.680 ;
        RECT 209.480 72.870 213.150 73.680 ;
        RECT 213.630 72.810 214.060 73.595 ;
        RECT 214.080 73.000 223.270 73.680 ;
        RECT 218.590 72.780 219.520 73.000 ;
        RECT 222.350 72.770 223.270 73.000 ;
        RECT 223.280 72.870 228.790 73.680 ;
        RECT 229.720 72.770 232.930 73.680 ;
        RECT 232.940 72.870 235.690 73.680 ;
        RECT 235.700 72.770 239.355 73.680 ;
        RECT 239.390 72.810 239.820 73.595 ;
        RECT 239.840 72.870 241.210 73.680 ;
        RECT 241.235 72.770 244.890 73.680 ;
        RECT 244.900 72.870 250.410 73.680 ;
        RECT 250.420 72.870 255.930 73.680 ;
        RECT 255.940 72.870 257.770 73.680 ;
        RECT 258.240 72.770 261.450 73.680 ;
        RECT 261.460 72.770 264.670 73.680 ;
        RECT 265.150 72.810 265.580 73.595 ;
        RECT 265.600 72.870 271.110 73.680 ;
        RECT 271.120 72.870 273.870 73.680 ;
        RECT 274.350 72.770 277.550 73.680 ;
        RECT 277.560 73.000 286.750 73.680 ;
        RECT 286.760 73.000 290.660 73.680 ;
        RECT 277.560 72.770 278.480 73.000 ;
        RECT 281.310 72.780 282.240 73.000 ;
        RECT 286.760 72.770 287.690 73.000 ;
        RECT 290.910 72.810 291.340 73.595 ;
        RECT 291.360 72.870 296.870 73.680 ;
        RECT 296.880 73.000 306.490 73.680 ;
        RECT 307.000 73.000 308.830 73.680 ;
        RECT 301.390 72.780 302.320 73.000 ;
        RECT 305.150 72.770 306.490 73.000 ;
        RECT 307.485 72.770 308.830 73.000 ;
        RECT 309.760 72.870 311.130 73.680 ;
      LAYER nwell ;
        RECT 161.905 69.650 311.325 72.480 ;
      LAYER pwell ;
        RECT 162.100 68.450 163.470 69.260 ;
        RECT 163.480 68.450 168.990 69.260 ;
        RECT 169.000 68.450 170.830 69.260 ;
        RECT 170.840 69.130 171.770 69.360 ;
        RECT 170.840 68.450 174.740 69.130 ;
        RECT 174.990 68.535 175.420 69.320 ;
        RECT 175.440 69.130 176.370 69.360 ;
        RECT 175.440 68.450 179.340 69.130 ;
        RECT 179.580 68.450 183.250 69.260 ;
        RECT 183.260 68.680 187.850 69.360 ;
        RECT 184.220 68.450 187.850 68.680 ;
        RECT 188.095 68.450 192.910 69.130 ;
        RECT 193.840 68.680 198.430 69.360 ;
        RECT 194.800 68.450 198.430 68.680 ;
        RECT 198.440 68.450 200.270 69.260 ;
        RECT 200.750 68.535 201.180 69.320 ;
        RECT 201.200 69.130 202.130 69.360 ;
        RECT 201.200 68.450 205.100 69.130 ;
        RECT 205.340 68.450 210.850 69.260 ;
        RECT 211.975 68.450 215.450 69.360 ;
        RECT 215.460 68.450 220.970 69.260 ;
        RECT 220.980 68.450 226.490 69.260 ;
        RECT 226.510 68.535 226.940 69.320 ;
        RECT 226.960 68.450 232.470 69.260 ;
        RECT 233.400 69.130 234.535 69.360 ;
        RECT 233.400 68.450 236.610 69.130 ;
        RECT 236.620 68.450 240.290 69.260 ;
        RECT 241.230 69.130 244.230 69.360 ;
        RECT 241.230 69.040 245.810 69.130 ;
        RECT 241.220 68.680 245.810 69.040 ;
        RECT 241.220 68.490 242.150 68.680 ;
        RECT 241.230 68.450 242.150 68.490 ;
        RECT 244.240 68.450 245.810 68.680 ;
        RECT 245.820 68.450 249.475 69.360 ;
        RECT 249.500 68.450 252.250 69.260 ;
        RECT 252.270 68.535 252.700 69.320 ;
        RECT 252.720 68.450 256.390 69.260 ;
        RECT 256.400 68.450 257.770 69.260 ;
        RECT 257.780 68.450 261.435 69.360 ;
        RECT 261.460 68.450 265.115 69.360 ;
        RECT 266.475 69.160 267.430 69.360 ;
        RECT 265.150 68.480 267.430 69.160 ;
        RECT 162.240 68.240 162.410 68.450 ;
        RECT 163.620 68.240 163.790 68.450 ;
        RECT 166.375 68.290 166.495 68.400 ;
        RECT 169.140 68.260 169.310 68.450 ;
        RECT 171.255 68.260 171.425 68.450 ;
        RECT 175.580 68.240 175.750 68.430 ;
        RECT 175.855 68.260 176.025 68.450 ;
        RECT 176.050 68.285 176.210 68.395 ;
        RECT 176.960 68.240 177.130 68.430 ;
        RECT 179.720 68.260 179.890 68.450 ;
        RECT 186.620 68.240 186.790 68.430 ;
        RECT 187.535 68.260 187.705 68.450 ;
        RECT 191.225 68.240 191.395 68.430 ;
        RECT 192.600 68.260 192.770 68.450 ;
        RECT 193.060 68.240 193.230 68.430 ;
        RECT 193.520 68.240 193.690 68.430 ;
        RECT 196.275 68.290 196.395 68.400 ;
        RECT 196.745 68.240 196.915 68.430 ;
        RECT 198.115 68.260 198.285 68.450 ;
        RECT 198.580 68.260 198.750 68.450 ;
        RECT 200.420 68.400 200.590 68.430 ;
        RECT 200.415 68.290 200.590 68.400 ;
        RECT 200.420 68.240 200.590 68.290 ;
        RECT 201.615 68.260 201.785 68.450 ;
        RECT 202.260 68.240 202.430 68.430 ;
        RECT 205.480 68.260 205.650 68.450 ;
        RECT 210.080 68.240 210.250 68.430 ;
        RECT 211.010 68.295 211.170 68.405 ;
        RECT 213.295 68.240 213.465 68.430 ;
        RECT 214.225 68.240 214.395 68.430 ;
        RECT 215.135 68.260 215.305 68.450 ;
        RECT 215.600 68.260 215.770 68.450 ;
        RECT 217.900 68.240 218.070 68.430 ;
        RECT 221.120 68.240 221.290 68.450 ;
        RECT 226.185 68.260 226.355 68.430 ;
        RECT 226.635 68.290 226.755 68.400 ;
        RECT 227.100 68.260 227.270 68.450 ;
        RECT 228.940 68.260 229.110 68.430 ;
        RECT 226.185 68.240 226.320 68.260 ;
        RECT 228.940 68.240 229.090 68.260 ;
        RECT 229.400 68.240 229.570 68.430 ;
        RECT 232.630 68.295 232.790 68.405 ;
        RECT 234.920 68.240 235.090 68.430 ;
        RECT 236.300 68.260 236.470 68.450 ;
        RECT 236.760 68.260 236.930 68.450 ;
        RECT 238.610 68.285 238.770 68.395 ;
        RECT 240.450 68.295 240.610 68.405 ;
        RECT 245.500 68.260 245.670 68.450 ;
        RECT 245.965 68.260 246.135 68.450 ;
        RECT 248.720 68.240 248.890 68.430 ;
        RECT 249.180 68.240 249.350 68.430 ;
        RECT 249.640 68.260 249.810 68.450 ;
        RECT 252.860 68.260 253.030 68.450 ;
        RECT 254.700 68.240 254.870 68.430 ;
        RECT 256.540 68.260 256.710 68.450 ;
        RECT 257.925 68.260 258.095 68.450 ;
        RECT 258.380 68.260 258.550 68.430 ;
        RECT 261.605 68.260 261.775 68.450 ;
        RECT 258.400 68.240 258.550 68.260 ;
        RECT 162.100 67.430 163.470 68.240 ;
        RECT 163.480 67.430 166.230 68.240 ;
        RECT 166.700 67.560 175.890 68.240 ;
        RECT 176.820 67.560 186.430 68.240 ;
        RECT 166.700 67.330 167.620 67.560 ;
        RECT 170.450 67.340 171.380 67.560 ;
        RECT 181.330 67.340 182.260 67.560 ;
        RECT 185.090 67.330 186.430 67.560 ;
        RECT 186.480 67.430 187.850 68.240 ;
        RECT 187.870 67.370 188.300 68.155 ;
        RECT 188.320 67.330 191.520 68.240 ;
        RECT 191.540 67.560 193.370 68.240 ;
        RECT 193.380 67.430 196.130 68.240 ;
        RECT 196.600 67.330 200.075 68.240 ;
        RECT 200.280 67.560 202.110 68.240 ;
        RECT 200.765 67.330 202.110 67.560 ;
        RECT 202.120 67.430 207.630 68.240 ;
        RECT 207.640 67.330 210.390 68.240 ;
        RECT 210.690 67.330 213.610 68.240 ;
        RECT 213.630 67.370 214.060 68.155 ;
        RECT 214.080 67.330 217.555 68.240 ;
        RECT 217.760 67.330 220.970 68.240 ;
        RECT 220.980 67.430 222.810 68.240 ;
        RECT 222.820 67.330 226.320 68.240 ;
        RECT 227.160 67.420 229.090 68.240 ;
        RECT 229.260 67.430 234.770 68.240 ;
        RECT 234.780 67.430 238.450 68.240 ;
        RECT 227.160 67.330 228.110 67.420 ;
        RECT 239.390 67.370 239.820 68.155 ;
        RECT 239.925 67.560 249.030 68.240 ;
        RECT 249.040 67.430 254.550 68.240 ;
        RECT 254.560 67.430 258.230 68.240 ;
        RECT 258.400 67.420 260.330 68.240 ;
        RECT 259.380 67.330 260.330 67.420 ;
        RECT 260.540 68.210 261.485 68.240 ;
        RECT 262.975 68.210 263.145 68.430 ;
        RECT 263.440 68.240 263.610 68.430 ;
        RECT 265.275 68.260 265.445 68.480 ;
        RECT 266.475 68.450 267.430 68.480 ;
        RECT 267.440 68.450 269.270 69.260 ;
        RECT 269.450 68.680 273.800 69.360 ;
        RECT 269.450 68.450 273.220 68.680 ;
        RECT 273.880 68.450 275.250 69.260 ;
        RECT 275.260 68.450 278.010 69.360 ;
        RECT 278.030 68.535 278.460 69.320 ;
        RECT 282.990 69.130 283.920 69.350 ;
        RECT 286.750 69.130 287.670 69.360 ;
        RECT 278.480 68.450 287.670 69.130 ;
        RECT 287.680 68.450 291.350 69.260 ;
        RECT 295.870 69.130 296.800 69.350 ;
        RECT 299.630 69.130 300.550 69.360 ;
        RECT 291.360 68.450 300.550 69.130 ;
        RECT 301.030 68.450 303.770 69.130 ;
        RECT 303.790 68.535 304.220 69.320 ;
        RECT 304.240 69.130 305.170 69.360 ;
        RECT 304.240 68.450 308.140 69.130 ;
        RECT 308.380 68.450 309.750 69.260 ;
        RECT 309.760 68.450 311.130 69.260 ;
        RECT 265.740 68.240 265.910 68.430 ;
        RECT 267.580 68.260 267.750 68.450 ;
        RECT 269.450 68.430 269.590 68.450 ;
        RECT 269.420 68.240 269.590 68.430 ;
        RECT 270.805 68.240 270.975 68.430 ;
        RECT 273.100 68.240 273.270 68.430 ;
        RECT 274.020 68.260 274.190 68.450 ;
        RECT 277.700 68.260 277.870 68.450 ;
        RECT 278.620 68.260 278.790 68.450 ;
        RECT 279.815 68.240 279.985 68.430 ;
        RECT 285.980 68.240 286.150 68.430 ;
        RECT 286.440 68.240 286.610 68.430 ;
        RECT 287.820 68.260 287.990 68.450 ;
        RECT 290.130 68.285 290.290 68.395 ;
        RECT 291.500 68.260 291.670 68.450 ;
        RECT 291.775 68.240 291.945 68.430 ;
        RECT 295.640 68.240 295.810 68.430 ;
        RECT 298.395 68.290 298.515 68.400 ;
        RECT 298.860 68.240 299.030 68.430 ;
        RECT 300.695 68.290 300.815 68.400 ;
        RECT 303.460 68.260 303.630 68.450 ;
        RECT 304.655 68.260 304.825 68.450 ;
        RECT 308.520 68.260 308.690 68.450 ;
        RECT 309.440 68.240 309.610 68.430 ;
        RECT 310.820 68.240 310.990 68.450 ;
        RECT 260.540 67.530 263.290 68.210 ;
        RECT 260.540 67.330 261.485 67.530 ;
        RECT 263.300 67.430 265.130 68.240 ;
        RECT 265.150 67.370 265.580 68.155 ;
        RECT 265.600 67.430 269.270 68.240 ;
        RECT 269.280 67.430 270.650 68.240 ;
        RECT 270.660 67.330 272.870 68.240 ;
        RECT 272.960 67.430 278.470 68.240 ;
        RECT 279.400 67.560 283.300 68.240 ;
        RECT 279.400 67.330 280.330 67.560 ;
        RECT 283.540 67.330 286.290 68.240 ;
        RECT 286.300 67.430 289.970 68.240 ;
        RECT 290.910 67.370 291.340 68.155 ;
        RECT 291.360 67.560 295.260 68.240 ;
        RECT 291.360 67.330 292.290 67.560 ;
        RECT 295.500 67.430 298.250 68.240 ;
        RECT 298.720 67.560 308.330 68.240 ;
        RECT 303.230 67.340 304.160 67.560 ;
        RECT 306.990 67.330 308.330 67.560 ;
        RECT 308.380 67.460 309.750 68.240 ;
        RECT 309.760 67.430 311.130 68.240 ;
      LAYER nwell ;
        RECT 161.905 64.210 311.325 67.040 ;
      LAYER pwell ;
        RECT 162.100 63.010 163.470 63.820 ;
        RECT 163.480 63.010 165.310 63.820 ;
        RECT 165.360 63.690 166.700 63.920 ;
        RECT 169.530 63.690 170.460 63.910 ;
        RECT 165.360 63.010 174.970 63.690 ;
        RECT 174.990 63.095 175.420 63.880 ;
        RECT 175.440 63.690 176.370 63.920 ;
        RECT 180.500 63.690 181.430 63.920 ;
        RECT 175.440 63.010 179.340 63.690 ;
        RECT 180.500 63.010 184.400 63.690 ;
        RECT 185.620 63.010 187.390 63.920 ;
        RECT 187.400 63.010 191.070 63.820 ;
        RECT 191.080 63.010 192.450 63.820 ;
        RECT 193.795 63.720 194.750 63.920 ;
        RECT 192.470 63.040 194.750 63.720 ;
        RECT 162.240 62.800 162.410 63.010 ;
        RECT 163.620 62.820 163.790 63.010 ;
        RECT 165.000 62.800 165.170 62.990 ;
        RECT 165.460 62.800 165.630 62.990 ;
        RECT 174.660 62.820 174.830 63.010 ;
        RECT 175.855 62.820 176.025 63.010 ;
        RECT 178.340 62.800 178.510 62.990 ;
        RECT 179.730 62.855 179.890 62.965 ;
        RECT 180.915 62.820 181.085 63.010 ;
        RECT 181.100 62.820 181.270 62.990 ;
        RECT 181.100 62.800 181.240 62.820 ;
        RECT 181.560 62.800 181.730 62.990 ;
        RECT 184.790 62.855 184.950 62.965 ;
        RECT 187.075 62.820 187.245 63.010 ;
        RECT 187.540 62.820 187.710 63.010 ;
        RECT 191.220 62.990 191.390 63.010 ;
        RECT 192.595 62.990 192.765 63.040 ;
        RECT 193.795 63.010 194.750 63.040 ;
        RECT 194.830 63.240 198.885 63.920 ;
        RECT 194.830 63.010 198.750 63.240 ;
        RECT 198.900 63.010 200.730 63.820 ;
        RECT 200.750 63.095 201.180 63.880 ;
        RECT 201.200 63.010 204.675 63.920 ;
        RECT 204.880 63.010 208.550 63.820 ;
        RECT 208.755 63.010 212.230 63.920 ;
        RECT 212.435 63.010 215.910 63.920 ;
        RECT 216.115 63.010 219.590 63.920 ;
        RECT 219.800 63.830 220.750 63.920 ;
        RECT 219.800 63.010 221.730 63.830 ;
        RECT 221.900 63.010 225.570 63.820 ;
        RECT 226.510 63.095 226.940 63.880 ;
        RECT 226.960 63.010 232.470 63.820 ;
        RECT 232.480 63.010 237.990 63.820 ;
        RECT 238.000 63.010 240.750 63.820 ;
        RECT 240.760 63.010 244.880 63.920 ;
        RECT 244.900 63.010 246.730 63.690 ;
        RECT 246.740 63.010 252.250 63.820 ;
        RECT 252.270 63.095 252.700 63.880 ;
        RECT 252.720 63.010 258.230 63.820 ;
        RECT 258.240 63.010 263.750 63.820 ;
        RECT 263.760 63.010 269.270 63.820 ;
        RECT 271.540 63.720 272.950 63.920 ;
        RECT 270.215 63.040 272.950 63.720 ;
        RECT 191.215 62.820 191.390 62.990 ;
        RECT 192.590 62.820 192.765 62.990 ;
        RECT 187.540 62.800 187.680 62.820 ;
        RECT 191.215 62.800 191.385 62.820 ;
        RECT 192.590 62.800 192.760 62.820 ;
        RECT 193.065 62.800 193.235 62.990 ;
        RECT 196.275 62.850 196.395 62.960 ;
        RECT 196.740 62.800 196.910 62.990 ;
        RECT 198.580 62.820 198.750 63.010 ;
        RECT 199.040 62.820 199.210 63.010 ;
        RECT 200.880 62.800 201.050 62.990 ;
        RECT 201.345 62.820 201.515 63.010 ;
        RECT 205.020 62.820 205.190 63.010 ;
        RECT 206.400 62.800 206.570 62.990 ;
        RECT 208.235 62.850 208.355 62.960 ;
        RECT 208.700 62.800 208.870 62.990 ;
        RECT 211.915 62.820 212.085 63.010 ;
        RECT 212.850 62.845 213.010 62.955 ;
        RECT 214.220 62.800 214.390 62.990 ;
        RECT 215.595 62.820 215.765 63.010 ;
        RECT 218.360 62.800 218.530 62.990 ;
        RECT 219.275 62.820 219.445 63.010 ;
        RECT 221.580 62.990 221.730 63.010 ;
        RECT 220.200 62.800 220.370 62.990 ;
        RECT 221.580 62.820 221.750 62.990 ;
        RECT 222.040 62.820 222.210 63.010 ;
        RECT 223.415 62.850 223.535 62.960 ;
        RECT 225.730 62.855 225.890 62.965 ;
        RECT 227.100 62.800 227.270 63.010 ;
        RECT 227.560 62.800 227.730 62.990 ;
        RECT 230.595 62.800 230.765 62.990 ;
        RECT 232.620 62.820 232.790 63.010 ;
        RECT 234.735 62.800 234.905 62.990 ;
        RECT 238.140 62.820 238.310 63.010 ;
        RECT 238.610 62.845 238.770 62.955 ;
        RECT 240.900 62.820 241.070 63.010 ;
        RECT 242.740 62.820 242.910 63.010 ;
        RECT 243.200 62.800 243.370 62.990 ;
        RECT 245.040 62.820 245.210 63.010 ;
        RECT 246.880 62.800 247.050 63.010 ;
        RECT 247.350 62.800 247.520 62.990 ;
        RECT 251.020 62.800 251.190 62.990 ;
        RECT 251.755 62.800 251.925 62.990 ;
        RECT 252.860 62.820 253.030 63.010 ;
        RECT 255.620 62.800 255.790 62.990 ;
        RECT 162.100 61.990 163.470 62.800 ;
        RECT 163.480 62.120 165.310 62.800 ;
        RECT 163.480 61.890 164.825 62.120 ;
        RECT 165.320 61.990 168.990 62.800 ;
        RECT 169.040 62.120 178.650 62.800 ;
        RECT 169.040 61.890 170.380 62.120 ;
        RECT 173.210 61.900 174.140 62.120 ;
        RECT 178.670 61.980 181.240 62.800 ;
        RECT 181.420 61.990 185.090 62.800 ;
        RECT 185.110 61.980 187.680 62.800 ;
        RECT 178.670 61.890 180.260 61.980 ;
        RECT 185.110 61.890 186.700 61.980 ;
        RECT 187.870 61.930 188.300 62.715 ;
        RECT 188.320 61.890 191.530 62.800 ;
        RECT 191.540 62.020 192.910 62.800 ;
        RECT 192.920 62.120 196.130 62.800 ;
        RECT 194.765 61.890 196.130 62.120 ;
        RECT 196.600 61.890 200.660 62.800 ;
        RECT 200.740 61.990 206.250 62.800 ;
        RECT 206.260 61.990 208.090 62.800 ;
        RECT 208.560 61.890 212.620 62.800 ;
        RECT 213.630 61.930 214.060 62.715 ;
        RECT 214.080 61.890 218.140 62.800 ;
        RECT 218.220 61.990 220.050 62.800 ;
        RECT 220.140 61.890 223.140 62.800 ;
        RECT 223.835 62.120 227.300 62.800 ;
        RECT 223.835 61.890 224.755 62.120 ;
        RECT 227.420 61.990 230.170 62.800 ;
        RECT 230.180 62.120 234.080 62.800 ;
        RECT 234.320 62.120 238.220 62.800 ;
        RECT 230.180 61.890 231.110 62.120 ;
        RECT 234.320 61.890 235.250 62.120 ;
        RECT 239.390 61.930 239.820 62.715 ;
        RECT 239.935 62.120 243.400 62.800 ;
        RECT 243.520 62.120 247.190 62.800 ;
        RECT 239.935 61.890 240.855 62.120 ;
        RECT 243.520 61.890 244.450 62.120 ;
        RECT 247.200 62.020 248.570 62.800 ;
        RECT 248.580 61.890 251.330 62.800 ;
        RECT 251.340 62.120 255.240 62.800 ;
        RECT 251.340 61.890 252.270 62.120 ;
        RECT 255.480 61.990 257.310 62.800 ;
        RECT 257.460 62.770 257.630 62.990 ;
        RECT 258.380 62.820 258.550 63.010 ;
        RECT 263.900 62.800 264.070 63.010 ;
        RECT 264.370 62.845 264.530 62.955 ;
        RECT 265.740 62.800 265.910 62.990 ;
        RECT 269.430 62.855 269.590 62.965 ;
        RECT 270.340 62.820 270.510 63.040 ;
        RECT 271.555 63.010 272.950 63.040 ;
        RECT 272.960 63.010 276.630 63.820 ;
        RECT 276.640 63.010 278.010 63.820 ;
        RECT 278.030 63.095 278.460 63.880 ;
        RECT 278.480 63.010 281.230 63.820 ;
        RECT 281.700 63.690 282.630 63.920 ;
        RECT 285.840 63.690 286.770 63.920 ;
        RECT 281.700 63.010 285.600 63.690 ;
        RECT 285.840 63.010 289.740 63.690 ;
        RECT 289.980 63.010 293.650 63.820 ;
        RECT 298.630 63.690 299.560 63.910 ;
        RECT 302.390 63.690 303.730 63.920 ;
        RECT 294.120 63.010 303.730 63.690 ;
        RECT 303.790 63.095 304.220 63.880 ;
        RECT 304.240 63.010 309.750 63.820 ;
        RECT 309.760 63.010 311.130 63.820 ;
        RECT 271.260 62.800 271.430 62.990 ;
        RECT 273.100 62.820 273.270 63.010 ;
        RECT 276.780 62.820 276.950 63.010 ;
        RECT 278.620 62.820 278.790 63.010 ;
        RECT 280.000 62.800 280.170 62.990 ;
        RECT 280.460 62.800 280.630 62.990 ;
        RECT 281.375 62.850 281.495 62.960 ;
        RECT 282.115 62.820 282.285 63.010 ;
        RECT 286.255 62.820 286.425 63.010 ;
        RECT 289.660 62.800 289.830 62.990 ;
        RECT 290.120 62.820 290.290 63.010 ;
        RECT 291.500 62.800 291.670 62.990 ;
        RECT 294.260 62.960 294.430 63.010 ;
        RECT 293.795 62.850 293.915 62.960 ;
        RECT 294.255 62.850 294.430 62.960 ;
        RECT 294.260 62.820 294.430 62.850 ;
        RECT 298.125 62.800 298.295 62.990 ;
        RECT 299.135 62.800 299.305 62.990 ;
        RECT 303.275 62.800 303.445 62.990 ;
        RECT 304.380 62.820 304.550 63.010 ;
        RECT 307.140 62.800 307.310 62.990 ;
        RECT 310.820 62.800 310.990 63.010 ;
        RECT 259.620 62.770 260.990 62.800 ;
        RECT 257.320 62.090 260.990 62.770 ;
        RECT 259.605 61.890 260.990 62.090 ;
        RECT 261.000 62.120 264.210 62.800 ;
        RECT 261.000 61.890 262.135 62.120 ;
        RECT 265.150 61.930 265.580 62.715 ;
        RECT 265.600 61.990 271.110 62.800 ;
        RECT 271.120 61.990 276.630 62.800 ;
        RECT 277.560 61.890 280.310 62.800 ;
        RECT 280.320 62.120 289.510 62.800 ;
        RECT 284.830 61.900 285.760 62.120 ;
        RECT 288.590 61.890 289.510 62.120 ;
        RECT 289.520 61.990 290.890 62.800 ;
        RECT 290.910 61.930 291.340 62.715 ;
        RECT 291.360 61.990 294.110 62.800 ;
        RECT 294.810 62.120 298.710 62.800 ;
        RECT 297.780 61.890 298.710 62.120 ;
        RECT 298.720 62.120 302.620 62.800 ;
        RECT 302.860 62.120 306.760 62.800 ;
        RECT 298.720 61.890 299.650 62.120 ;
        RECT 302.860 61.890 303.790 62.120 ;
        RECT 307.000 61.990 309.750 62.800 ;
        RECT 309.760 61.990 311.130 62.800 ;
      LAYER nwell ;
        RECT 161.905 58.770 311.325 61.600 ;
      LAYER pwell ;
        RECT 162.100 57.570 163.470 58.380 ;
        RECT 163.480 57.570 168.990 58.380 ;
        RECT 169.000 57.570 170.830 58.380 ;
        RECT 170.840 58.250 171.770 58.480 ;
        RECT 170.840 57.570 174.740 58.250 ;
        RECT 174.990 57.655 175.420 58.440 ;
        RECT 175.440 58.250 176.785 58.480 ;
        RECT 177.750 58.390 179.340 58.480 ;
        RECT 175.440 57.570 177.270 58.250 ;
        RECT 177.750 57.570 180.320 58.390 ;
        RECT 180.500 57.570 181.870 58.380 ;
        RECT 182.015 58.250 185.525 58.480 ;
        RECT 182.015 57.570 186.010 58.250 ;
        RECT 186.040 57.570 191.530 58.480 ;
        RECT 191.540 57.570 195.575 58.480 ;
        RECT 196.820 58.390 197.770 58.480 ;
        RECT 195.840 57.570 197.770 58.390 ;
        RECT 197.980 57.570 200.730 58.380 ;
        RECT 200.750 57.655 201.180 58.440 ;
        RECT 201.280 57.570 204.280 58.480 ;
        RECT 204.420 57.570 209.930 58.380 ;
        RECT 209.940 57.570 212.690 58.380 ;
        RECT 213.330 57.570 216.830 58.480 ;
        RECT 216.920 57.570 219.920 58.480 ;
        RECT 220.060 58.250 220.990 58.480 ;
        RECT 224.510 58.250 225.440 58.480 ;
        RECT 220.060 57.570 223.960 58.250 ;
        RECT 224.510 57.570 226.345 58.250 ;
        RECT 226.510 57.655 226.940 58.440 ;
        RECT 229.615 58.250 230.535 58.480 ;
        RECT 227.070 57.570 230.535 58.250 ;
        RECT 230.640 57.570 232.470 58.380 ;
        RECT 236.990 58.250 237.920 58.470 ;
        RECT 240.750 58.250 241.670 58.480 ;
        RECT 244.420 58.250 245.350 58.480 ;
        RECT 232.480 57.570 241.670 58.250 ;
        RECT 241.680 57.570 245.350 58.250 ;
        RECT 245.360 57.570 246.730 58.380 ;
        RECT 246.740 57.570 248.110 58.350 ;
        RECT 251.320 58.250 252.250 58.480 ;
        RECT 248.350 57.570 252.250 58.250 ;
        RECT 252.270 57.655 252.700 58.440 ;
        RECT 257.230 58.250 258.160 58.470 ;
        RECT 260.990 58.250 261.910 58.480 ;
        RECT 252.720 57.570 261.910 58.250 ;
        RECT 261.920 57.570 267.430 58.380 ;
        RECT 268.430 57.800 272.780 58.480 ;
        RECT 269.010 57.570 272.780 57.800 ;
        RECT 272.960 57.570 276.630 58.380 ;
        RECT 276.640 57.570 278.010 58.380 ;
        RECT 278.030 57.655 278.460 58.440 ;
        RECT 281.680 58.250 282.610 58.480 ;
        RECT 288.050 58.250 288.980 58.470 ;
        RECT 291.810 58.250 293.150 58.480 ;
        RECT 278.710 57.570 282.610 58.250 ;
        RECT 283.540 57.570 293.150 58.250 ;
        RECT 293.200 57.570 294.570 58.380 ;
        RECT 294.580 58.250 295.500 58.480 ;
        RECT 298.330 58.250 299.260 58.470 ;
        RECT 294.580 57.570 303.770 58.250 ;
        RECT 303.790 57.655 304.220 58.440 ;
        RECT 304.240 57.570 309.750 58.380 ;
        RECT 309.760 57.570 311.130 58.380 ;
        RECT 162.240 57.360 162.410 57.570 ;
        RECT 163.620 57.360 163.790 57.570 ;
        RECT 166.380 57.360 166.550 57.550 ;
        RECT 169.140 57.380 169.310 57.570 ;
        RECT 171.255 57.380 171.425 57.570 ;
        RECT 175.855 57.360 176.025 57.550 ;
        RECT 176.960 57.380 177.130 57.570 ;
        RECT 180.180 57.550 180.320 57.570 ;
        RECT 177.415 57.410 177.535 57.520 ;
        RECT 180.180 57.380 180.350 57.550 ;
        RECT 180.640 57.380 180.810 57.570 ;
        RECT 182.020 57.380 182.190 57.550 ;
        RECT 182.490 57.405 182.650 57.515 ;
        RECT 182.020 57.360 182.160 57.380 ;
        RECT 183.405 57.360 183.575 57.550 ;
        RECT 185.695 57.380 185.865 57.570 ;
        RECT 187.075 57.360 187.245 57.550 ;
        RECT 187.535 57.410 187.655 57.520 ;
        RECT 191.215 57.380 191.385 57.570 ;
        RECT 191.685 57.550 191.855 57.570 ;
        RECT 195.840 57.550 195.990 57.570 ;
        RECT 191.680 57.380 191.855 57.550 ;
        RECT 191.680 57.360 191.850 57.380 ;
        RECT 192.140 57.360 192.310 57.550 ;
        RECT 195.360 57.360 195.530 57.550 ;
        RECT 195.820 57.380 195.990 57.550 ;
        RECT 198.120 57.380 198.290 57.570 ;
        RECT 201.340 57.380 201.510 57.570 ;
        RECT 204.560 57.380 204.730 57.570 ;
        RECT 206.400 57.380 206.570 57.550 ;
        RECT 206.400 57.360 206.565 57.380 ;
        RECT 206.860 57.360 207.030 57.550 ;
        RECT 210.080 57.380 210.250 57.570 ;
        RECT 213.330 57.550 213.465 57.570 ;
        RECT 210.550 57.405 210.710 57.515 ;
        RECT 211.460 57.380 211.630 57.550 ;
        RECT 212.835 57.410 212.955 57.520 ;
        RECT 213.295 57.380 213.465 57.550 ;
        RECT 211.465 57.360 211.630 57.380 ;
        RECT 214.220 57.360 214.390 57.550 ;
        RECT 216.980 57.380 217.150 57.570 ;
        RECT 218.820 57.360 218.990 57.550 ;
        RECT 219.280 57.360 219.450 57.550 ;
        RECT 220.475 57.380 220.645 57.570 ;
        RECT 226.180 57.550 226.345 57.570 ;
        RECT 226.180 57.380 226.350 57.550 ;
        RECT 227.100 57.380 227.270 57.570 ;
        RECT 228.480 57.360 228.650 57.550 ;
        RECT 230.780 57.380 230.950 57.570 ;
        RECT 232.620 57.380 232.790 57.570 ;
        RECT 237.680 57.360 237.850 57.550 ;
        RECT 241.820 57.380 241.990 57.570 ;
        RECT 244.120 57.380 244.290 57.550 ;
        RECT 245.500 57.380 245.670 57.570 ;
        RECT 246.890 57.550 247.060 57.570 ;
        RECT 246.420 57.380 246.590 57.550 ;
        RECT 246.880 57.380 247.060 57.550 ;
        RECT 250.570 57.405 250.730 57.515 ;
        RECT 241.820 57.360 241.985 57.380 ;
        RECT 244.120 57.360 244.285 57.380 ;
        RECT 246.420 57.360 246.585 57.380 ;
        RECT 246.880 57.360 247.050 57.380 ;
        RECT 251.480 57.360 251.650 57.550 ;
        RECT 251.665 57.380 251.835 57.570 ;
        RECT 252.860 57.380 253.030 57.570 ;
        RECT 262.060 57.380 262.230 57.570 ;
        RECT 272.640 57.550 272.780 57.570 ;
        RECT 262.980 57.360 263.150 57.550 ;
        RECT 263.440 57.360 263.610 57.550 ;
        RECT 267.590 57.415 267.750 57.525 ;
        RECT 268.960 57.360 269.130 57.550 ;
        RECT 269.420 57.360 269.590 57.550 ;
        RECT 272.640 57.380 272.810 57.550 ;
        RECT 273.100 57.380 273.270 57.570 ;
        RECT 276.780 57.380 276.950 57.570 ;
        RECT 282.025 57.380 282.195 57.570 ;
        RECT 282.770 57.415 282.930 57.525 ;
        RECT 283.680 57.360 283.850 57.570 ;
        RECT 284.140 57.360 284.310 57.550 ;
        RECT 290.120 57.360 290.290 57.550 ;
        RECT 290.575 57.410 290.695 57.520 ;
        RECT 291.500 57.360 291.670 57.550 ;
        RECT 293.340 57.380 293.510 57.570 ;
        RECT 296.560 57.360 296.730 57.550 ;
        RECT 299.315 57.410 299.435 57.520 ;
        RECT 299.780 57.360 299.950 57.550 ;
        RECT 303.460 57.380 303.630 57.570 ;
        RECT 304.380 57.380 304.550 57.570 ;
        RECT 309.435 57.410 309.555 57.520 ;
        RECT 310.820 57.360 310.990 57.570 ;
        RECT 162.100 56.550 163.470 57.360 ;
        RECT 163.480 56.550 166.230 57.360 ;
        RECT 166.240 56.680 175.430 57.360 ;
        RECT 170.750 56.460 171.680 56.680 ;
        RECT 174.510 56.450 175.430 56.680 ;
        RECT 175.440 56.680 179.340 57.360 ;
        RECT 175.440 56.450 176.370 56.680 ;
        RECT 179.590 56.540 182.160 57.360 ;
        RECT 179.590 56.450 181.180 56.540 ;
        RECT 183.260 56.450 185.030 57.360 ;
        RECT 185.555 57.130 187.245 57.360 ;
        RECT 185.555 56.450 187.390 57.130 ;
        RECT 187.870 56.490 188.300 57.275 ;
        RECT 188.320 56.680 191.990 57.360 ;
        RECT 192.000 56.680 195.210 57.360 ;
        RECT 195.220 56.680 204.410 57.360 ;
        RECT 188.320 56.450 189.250 56.680 ;
        RECT 194.075 56.450 195.210 56.680 ;
        RECT 199.730 56.460 200.660 56.680 ;
        RECT 203.490 56.450 204.410 56.680 ;
        RECT 204.730 56.680 206.565 57.360 ;
        RECT 204.730 56.450 205.660 56.680 ;
        RECT 206.720 56.550 210.390 57.360 ;
        RECT 211.465 56.680 213.300 57.360 ;
        RECT 212.370 56.450 213.300 56.680 ;
        RECT 213.630 56.490 214.060 57.275 ;
        RECT 214.080 56.550 215.450 57.360 ;
        RECT 215.555 56.680 219.020 57.360 ;
        RECT 219.140 56.680 228.330 57.360 ;
        RECT 228.340 56.680 237.530 57.360 ;
        RECT 215.555 56.450 216.475 56.680 ;
        RECT 223.650 56.460 224.580 56.680 ;
        RECT 227.410 56.450 228.330 56.680 ;
        RECT 232.850 56.460 233.780 56.680 ;
        RECT 236.610 56.450 237.530 56.680 ;
        RECT 237.540 56.550 239.370 57.360 ;
        RECT 239.390 56.490 239.820 57.275 ;
        RECT 240.150 56.680 241.985 57.360 ;
        RECT 242.450 56.680 244.285 57.360 ;
        RECT 244.750 56.680 246.585 57.360 ;
        RECT 240.150 56.450 241.080 56.680 ;
        RECT 242.450 56.450 243.380 56.680 ;
        RECT 244.750 56.450 245.680 56.680 ;
        RECT 246.740 56.550 250.410 57.360 ;
        RECT 251.340 56.680 260.530 57.360 ;
        RECT 255.850 56.460 256.780 56.680 ;
        RECT 259.610 56.450 260.530 56.680 ;
        RECT 261.200 56.550 263.290 57.360 ;
        RECT 263.300 56.550 265.130 57.360 ;
        RECT 265.150 56.490 265.580 57.275 ;
        RECT 265.695 56.680 269.160 57.360 ;
        RECT 265.695 56.450 266.615 56.680 ;
        RECT 269.280 56.550 274.790 57.360 ;
        RECT 274.800 56.680 283.990 57.360 ;
        RECT 274.800 56.450 275.720 56.680 ;
        RECT 278.550 56.460 279.480 56.680 ;
        RECT 284.000 56.550 285.370 57.360 ;
        RECT 285.615 56.680 290.430 57.360 ;
        RECT 290.910 56.490 291.340 57.275 ;
        RECT 291.360 56.680 296.175 57.360 ;
        RECT 296.420 56.550 299.170 57.360 ;
        RECT 299.640 56.680 308.920 57.360 ;
        RECT 301.000 56.460 301.920 56.680 ;
        RECT 306.585 56.560 308.920 56.680 ;
        RECT 308.000 56.450 308.920 56.560 ;
        RECT 309.760 56.550 311.130 57.360 ;
      LAYER nwell ;
        RECT 161.905 53.330 311.325 56.160 ;
      LAYER pwell ;
        RECT 162.100 52.130 163.470 52.940 ;
        RECT 163.480 52.130 165.310 52.940 ;
        RECT 170.290 52.810 171.220 53.030 ;
        RECT 174.050 52.810 174.970 53.040 ;
        RECT 165.780 52.130 174.970 52.810 ;
        RECT 174.990 52.215 175.420 53.000 ;
        RECT 175.440 52.130 178.180 52.810 ;
        RECT 178.200 52.130 183.710 52.940 ;
        RECT 186.255 52.810 187.390 53.040 ;
        RECT 184.180 52.130 187.390 52.810 ;
        RECT 187.400 52.840 188.330 53.040 ;
        RECT 189.660 52.840 190.610 53.040 ;
        RECT 187.400 52.360 190.610 52.840 ;
        RECT 187.545 52.160 190.610 52.360 ;
        RECT 162.240 51.920 162.410 52.130 ;
        RECT 163.620 51.920 163.790 52.130 ;
        RECT 165.455 51.970 165.575 52.080 ;
        RECT 165.920 51.940 166.090 52.130 ;
        RECT 166.380 51.920 166.550 52.110 ;
        RECT 175.580 51.920 175.750 52.130 ;
        RECT 178.340 51.920 178.510 52.130 ;
        RECT 182.030 51.965 182.190 52.075 ;
        RECT 183.855 51.920 184.025 52.110 ;
        RECT 184.320 51.940 184.490 52.130 ;
        RECT 187.545 52.110 187.715 52.160 ;
        RECT 189.675 52.130 190.610 52.160 ;
        RECT 190.910 52.130 193.830 53.040 ;
        RECT 195.900 52.950 196.850 53.040 ;
        RECT 194.920 52.130 196.850 52.950 ;
        RECT 197.060 52.130 199.250 53.040 ;
        RECT 199.360 52.130 200.730 52.940 ;
        RECT 200.750 52.215 201.180 53.000 ;
        RECT 201.200 52.130 202.570 52.940 ;
        RECT 203.630 52.810 204.560 53.040 ;
        RECT 202.725 52.130 204.560 52.810 ;
        RECT 204.880 52.130 208.550 52.940 ;
        RECT 209.610 52.810 210.540 53.040 ;
        RECT 215.370 52.810 216.300 53.030 ;
        RECT 219.130 52.810 220.050 53.040 ;
        RECT 208.705 52.130 210.540 52.810 ;
        RECT 210.860 52.130 220.050 52.810 ;
        RECT 220.060 52.130 221.430 52.940 ;
        RECT 221.675 52.130 226.490 52.810 ;
        RECT 226.510 52.215 226.940 53.000 ;
        RECT 233.070 52.810 234.000 53.040 ;
        RECT 226.960 52.130 231.775 52.810 ;
        RECT 232.165 52.130 234.000 52.810 ;
        RECT 235.565 52.130 239.220 53.040 ;
        RECT 239.380 52.130 240.750 52.940 ;
        RECT 240.855 52.810 241.775 53.040 ;
        RECT 240.855 52.130 244.320 52.810 ;
        RECT 244.440 52.130 247.600 53.040 ;
        RECT 250.315 52.810 251.235 53.040 ;
        RECT 247.770 52.130 251.235 52.810 ;
        RECT 252.270 52.215 252.700 53.000 ;
        RECT 253.030 52.810 253.960 53.040 ;
        RECT 261.000 52.810 261.920 53.040 ;
        RECT 264.750 52.810 265.680 53.030 ;
        RECT 270.295 52.810 271.215 53.040 ;
        RECT 253.030 52.130 254.865 52.810 ;
        RECT 255.020 52.130 259.835 52.810 ;
        RECT 261.000 52.130 270.190 52.810 ;
        RECT 270.295 52.130 273.760 52.810 ;
        RECT 273.880 52.130 277.550 52.940 ;
        RECT 278.030 52.215 278.460 53.000 ;
        RECT 278.480 52.130 281.230 52.940 ;
        RECT 281.240 52.810 282.170 53.040 ;
        RECT 281.240 52.130 285.140 52.810 ;
        RECT 285.380 52.130 296.390 53.040 ;
        RECT 296.420 52.130 300.090 52.940 ;
        RECT 301.020 52.130 303.760 52.810 ;
        RECT 303.790 52.215 304.220 53.000 ;
        RECT 304.700 52.130 306.070 52.910 ;
        RECT 306.175 52.810 307.095 53.040 ;
        RECT 306.175 52.130 309.640 52.810 ;
        RECT 309.760 52.130 311.130 52.940 ;
        RECT 187.540 51.940 187.715 52.110 ;
        RECT 187.540 51.920 187.710 51.940 ;
        RECT 188.460 51.920 188.630 52.110 ;
        RECT 189.835 51.970 189.955 52.080 ;
        RECT 190.300 51.920 190.470 52.110 ;
        RECT 193.515 51.940 193.685 52.130 ;
        RECT 194.920 52.110 195.070 52.130 ;
        RECT 193.990 51.975 194.150 52.085 ;
        RECT 194.900 51.940 195.070 52.110 ;
        RECT 195.360 51.920 195.530 52.110 ;
        RECT 197.205 51.940 197.375 52.130 ;
        RECT 199.500 51.940 199.670 52.130 ;
        RECT 201.340 51.940 201.510 52.130 ;
        RECT 202.725 52.110 202.890 52.130 ;
        RECT 202.720 51.940 202.890 52.110 ;
        RECT 204.560 51.920 204.730 52.110 ;
        RECT 205.020 51.940 205.190 52.130 ;
        RECT 208.705 52.110 208.870 52.130 ;
        RECT 208.700 51.940 208.870 52.110 ;
        RECT 211.000 51.940 211.170 52.130 ;
        RECT 214.220 51.920 214.390 52.110 ;
        RECT 217.900 51.920 218.070 52.110 ;
        RECT 220.200 51.940 220.370 52.130 ;
        RECT 222.965 51.920 223.135 52.110 ;
        RECT 226.180 51.940 226.350 52.130 ;
        RECT 227.100 51.940 227.270 52.130 ;
        RECT 232.165 52.110 232.330 52.130 ;
        RECT 239.060 52.110 239.220 52.130 ;
        RECT 232.160 51.940 232.330 52.110 ;
        RECT 234.000 51.920 234.170 52.110 ;
        RECT 234.470 51.975 234.630 52.085 ;
        RECT 239.060 51.920 239.230 52.110 ;
        RECT 239.520 51.940 239.690 52.130 ;
        RECT 239.980 51.920 240.150 52.110 ;
        RECT 244.120 51.940 244.290 52.130 ;
        RECT 245.040 51.920 245.210 52.110 ;
        RECT 245.500 51.920 245.670 52.110 ;
        RECT 247.340 51.940 247.510 52.130 ;
        RECT 247.800 51.940 247.970 52.130 ;
        RECT 254.700 52.110 254.865 52.130 ;
        RECT 250.560 51.940 250.730 52.110 ;
        RECT 251.030 51.965 251.190 52.075 ;
        RECT 251.490 51.975 251.650 52.085 ;
        RECT 254.700 51.940 254.870 52.110 ;
        RECT 255.160 51.940 255.330 52.130 ;
        RECT 255.620 51.940 255.790 52.110 ;
        RECT 250.560 51.920 250.720 51.940 ;
        RECT 255.620 51.920 255.780 51.940 ;
        RECT 256.080 51.920 256.250 52.110 ;
        RECT 260.230 51.975 260.390 52.085 ;
        RECT 264.360 51.920 264.530 52.110 ;
        RECT 264.815 51.970 264.935 52.080 ;
        RECT 266.660 51.920 266.830 52.110 ;
        RECT 267.130 51.965 267.290 52.075 ;
        RECT 268.040 51.920 268.210 52.110 ;
        RECT 269.880 51.940 270.050 52.130 ;
        RECT 273.560 51.940 273.730 52.130 ;
        RECT 274.020 51.940 274.190 52.130 ;
        RECT 277.240 51.920 277.410 52.110 ;
        RECT 277.695 51.970 277.815 52.080 ;
        RECT 278.620 51.940 278.790 52.130 ;
        RECT 279.080 51.920 279.250 52.110 ;
        RECT 281.655 51.940 281.825 52.130 ;
        RECT 285.525 51.940 285.695 52.130 ;
        RECT 288.280 51.920 288.450 52.110 ;
        RECT 291.500 51.920 291.670 52.110 ;
        RECT 296.560 51.940 296.730 52.130 ;
        RECT 297.020 51.920 297.190 52.110 ;
        RECT 300.250 51.975 300.410 52.085 ;
        RECT 301.160 51.940 301.330 52.130 ;
        RECT 304.375 51.970 304.495 52.080 ;
        RECT 305.760 51.940 305.930 52.130 ;
        RECT 308.980 51.920 309.150 52.110 ;
        RECT 309.440 52.080 309.610 52.130 ;
        RECT 309.435 51.970 309.610 52.080 ;
        RECT 309.440 51.940 309.610 51.970 ;
        RECT 310.820 51.920 310.990 52.130 ;
        RECT 162.100 51.110 163.470 51.920 ;
        RECT 163.480 51.110 166.230 51.920 ;
        RECT 166.240 51.240 175.430 51.920 ;
        RECT 175.440 51.240 178.180 51.920 ;
        RECT 170.750 51.020 171.680 51.240 ;
        RECT 174.510 51.010 175.430 51.240 ;
        RECT 178.200 51.110 181.870 51.920 ;
        RECT 182.820 51.010 184.170 51.920 ;
        RECT 184.180 51.240 187.850 51.920 ;
        RECT 184.180 51.010 185.110 51.240 ;
        RECT 187.870 51.050 188.300 51.835 ;
        RECT 188.330 51.010 189.680 51.920 ;
        RECT 190.160 51.240 194.975 51.920 ;
        RECT 195.220 51.240 204.410 51.920 ;
        RECT 204.420 51.240 213.610 51.920 ;
        RECT 199.730 51.020 200.660 51.240 ;
        RECT 203.490 51.010 204.410 51.240 ;
        RECT 208.930 51.020 209.860 51.240 ;
        RECT 212.690 51.010 213.610 51.240 ;
        RECT 213.630 51.050 214.060 51.835 ;
        RECT 214.080 51.110 217.750 51.920 ;
        RECT 217.760 51.240 222.575 51.920 ;
        RECT 222.820 51.010 233.830 51.920 ;
        RECT 233.860 51.110 235.690 51.920 ;
        RECT 235.795 51.240 239.260 51.920 ;
        RECT 235.795 51.010 236.715 51.240 ;
        RECT 239.390 51.050 239.820 51.835 ;
        RECT 239.840 51.110 241.670 51.920 ;
        RECT 241.775 51.240 245.240 51.920 ;
        RECT 241.775 51.010 242.695 51.240 ;
        RECT 245.360 51.110 246.730 51.920 ;
        RECT 247.065 51.010 250.720 51.920 ;
        RECT 252.125 51.010 255.780 51.920 ;
        RECT 255.940 51.240 260.755 51.920 ;
        RECT 261.095 51.240 264.560 51.920 ;
        RECT 261.095 51.010 262.015 51.240 ;
        RECT 265.150 51.050 265.580 51.835 ;
        RECT 265.610 51.010 266.960 51.920 ;
        RECT 267.900 51.240 277.090 51.920 ;
        RECT 272.410 51.020 273.340 51.240 ;
        RECT 276.170 51.010 277.090 51.240 ;
        RECT 277.100 51.110 278.930 51.920 ;
        RECT 278.940 51.240 288.130 51.920 ;
        RECT 283.450 51.020 284.380 51.240 ;
        RECT 287.210 51.010 288.130 51.240 ;
        RECT 288.140 51.110 290.230 51.920 ;
        RECT 290.910 51.050 291.340 51.835 ;
        RECT 291.360 51.110 296.870 51.920 ;
        RECT 296.880 51.110 299.630 51.920 ;
        RECT 299.645 51.240 309.290 51.920 ;
        RECT 299.645 51.120 302.345 51.240 ;
        RECT 299.645 51.010 301.415 51.120 ;
        RECT 307.010 51.020 307.930 51.240 ;
        RECT 309.760 51.110 311.130 51.920 ;
      LAYER nwell ;
        RECT 161.905 47.890 311.325 50.720 ;
      LAYER pwell ;
        RECT 162.100 46.690 163.470 47.500 ;
        RECT 163.480 46.690 168.990 47.500 ;
        RECT 169.000 46.690 170.830 47.500 ;
        RECT 170.840 47.370 171.770 47.600 ;
        RECT 170.840 46.690 174.740 47.370 ;
        RECT 174.990 46.775 175.420 47.560 ;
        RECT 175.440 46.690 176.810 47.500 ;
        RECT 176.820 47.370 177.750 47.600 ;
        RECT 183.615 47.370 184.535 47.600 ;
        RECT 176.820 46.690 180.720 47.370 ;
        RECT 181.070 46.690 184.535 47.370 ;
        RECT 184.640 46.690 190.150 47.500 ;
        RECT 190.160 46.690 192.910 47.500 ;
        RECT 193.385 46.690 194.750 47.370 ;
        RECT 194.995 46.690 199.810 47.370 ;
        RECT 200.750 46.775 201.180 47.560 ;
        RECT 201.200 46.690 204.870 47.500 ;
        RECT 204.880 47.370 205.800 47.600 ;
        RECT 208.630 47.370 209.560 47.590 ;
        RECT 218.590 47.370 219.520 47.590 ;
        RECT 222.350 47.370 223.270 47.600 ;
        RECT 204.880 46.690 214.070 47.370 ;
        RECT 214.080 46.690 223.270 47.370 ;
        RECT 223.280 46.690 226.030 47.500 ;
        RECT 226.510 46.775 226.940 47.560 ;
        RECT 226.960 46.690 229.710 47.500 ;
        RECT 234.690 47.370 235.620 47.590 ;
        RECT 238.450 47.370 239.370 47.600 ;
        RECT 230.180 46.690 239.370 47.370 ;
        RECT 239.380 46.690 241.210 47.500 ;
        RECT 245.730 47.370 246.660 47.590 ;
        RECT 249.490 47.370 250.410 47.600 ;
        RECT 241.220 46.690 250.410 47.370 ;
        RECT 250.420 46.690 252.250 47.500 ;
        RECT 252.270 46.775 252.700 47.560 ;
        RECT 252.720 46.690 254.550 47.500 ;
        RECT 259.070 47.370 260.000 47.590 ;
        RECT 262.830 47.370 263.750 47.600 ;
        RECT 254.560 46.690 263.750 47.370 ;
        RECT 263.855 47.370 264.775 47.600 ;
        RECT 263.855 46.690 267.320 47.370 ;
        RECT 267.440 46.690 271.095 47.600 ;
        RECT 271.120 46.690 273.870 47.500 ;
        RECT 274.435 47.370 275.355 47.600 ;
        RECT 274.435 46.690 277.900 47.370 ;
        RECT 278.030 46.775 278.460 47.560 ;
        RECT 278.480 47.370 279.400 47.600 ;
        RECT 282.230 47.370 283.160 47.590 ;
        RECT 292.190 47.370 293.120 47.590 ;
        RECT 295.950 47.370 296.870 47.600 ;
        RECT 300.455 47.370 301.375 47.600 ;
        RECT 278.480 46.690 287.670 47.370 ;
        RECT 287.680 46.690 296.870 47.370 ;
        RECT 297.910 46.690 301.375 47.370 ;
        RECT 301.480 46.690 303.310 47.500 ;
        RECT 303.790 46.775 304.220 47.560 ;
        RECT 304.240 46.690 309.750 47.500 ;
        RECT 309.760 46.690 311.130 47.500 ;
        RECT 162.240 46.480 162.410 46.690 ;
        RECT 163.620 46.480 163.790 46.690 ;
        RECT 169.140 46.480 169.310 46.690 ;
        RECT 171.255 46.500 171.425 46.690 ;
        RECT 171.900 46.480 172.070 46.670 ;
        RECT 175.580 46.500 175.750 46.690 ;
        RECT 177.235 46.500 177.405 46.690 ;
        RECT 181.100 46.500 181.270 46.690 ;
        RECT 181.835 46.480 182.005 46.670 ;
        RECT 184.780 46.500 184.950 46.690 ;
        RECT 185.700 46.480 185.870 46.670 ;
        RECT 187.535 46.530 187.655 46.640 ;
        RECT 188.470 46.525 188.630 46.635 ;
        RECT 189.380 46.480 189.550 46.670 ;
        RECT 190.300 46.500 190.470 46.690 ;
        RECT 193.060 46.500 193.230 46.670 ;
        RECT 199.050 46.525 199.210 46.635 ;
        RECT 199.500 46.500 199.670 46.690 ;
        RECT 199.960 46.480 200.130 46.670 ;
        RECT 201.340 46.500 201.510 46.690 ;
        RECT 203.915 46.480 204.085 46.670 ;
        RECT 207.780 46.480 207.950 46.670 ;
        RECT 213.025 46.480 213.195 46.670 ;
        RECT 213.760 46.500 213.930 46.690 ;
        RECT 214.220 46.480 214.390 46.690 ;
        RECT 216.055 46.530 216.175 46.640 ;
        RECT 216.520 46.480 216.690 46.670 ;
        RECT 223.420 46.500 223.590 46.690 ;
        RECT 225.715 46.530 225.835 46.640 ;
        RECT 226.175 46.530 226.295 46.640 ;
        RECT 227.100 46.500 227.270 46.690 ;
        RECT 229.860 46.640 230.030 46.670 ;
        RECT 229.855 46.530 230.030 46.640 ;
        RECT 229.860 46.500 230.030 46.530 ;
        RECT 229.860 46.480 230.020 46.500 ;
        RECT 230.320 46.480 230.490 46.690 ;
        RECT 239.520 46.500 239.690 46.690 ;
        RECT 239.980 46.500 240.150 46.670 ;
        RECT 241.360 46.500 241.530 46.690 ;
        RECT 239.990 46.480 240.150 46.500 ;
        RECT 247.340 46.480 247.510 46.670 ;
        RECT 247.795 46.530 247.915 46.640 ;
        RECT 248.260 46.480 248.430 46.670 ;
        RECT 250.560 46.500 250.730 46.690 ;
        RECT 252.860 46.500 253.030 46.690 ;
        RECT 254.700 46.500 254.870 46.690 ;
        RECT 260.680 46.480 260.850 46.670 ;
        RECT 263.900 46.480 264.070 46.670 ;
        RECT 264.370 46.525 264.530 46.635 ;
        RECT 265.740 46.480 265.910 46.670 ;
        RECT 267.120 46.500 267.290 46.690 ;
        RECT 267.585 46.500 267.755 46.690 ;
        RECT 269.875 46.480 270.045 46.670 ;
        RECT 271.260 46.500 271.430 46.690 ;
        RECT 272.175 46.480 272.345 46.670 ;
        RECT 272.640 46.480 272.810 46.670 ;
        RECT 274.015 46.530 274.135 46.640 ;
        RECT 277.700 46.500 277.870 46.690 ;
        RECT 278.155 46.530 278.275 46.640 ;
        RECT 282.025 46.480 282.195 46.670 ;
        RECT 282.760 46.480 282.930 46.670 ;
        RECT 286.440 46.480 286.610 46.670 ;
        RECT 287.360 46.500 287.530 46.690 ;
        RECT 287.820 46.500 287.990 46.690 ;
        RECT 290.130 46.525 290.290 46.635 ;
        RECT 297.030 46.535 297.190 46.645 ;
        RECT 297.940 46.500 298.110 46.690 ;
        RECT 300.240 46.480 300.410 46.670 ;
        RECT 300.700 46.480 300.870 46.670 ;
        RECT 301.620 46.500 301.790 46.690 ;
        RECT 303.455 46.530 303.575 46.640 ;
        RECT 304.380 46.500 304.550 46.690 ;
        RECT 306.220 46.480 306.390 46.670 ;
        RECT 310.820 46.480 310.990 46.690 ;
        RECT 162.100 45.670 163.470 46.480 ;
        RECT 163.480 45.670 168.990 46.480 ;
        RECT 169.000 45.670 171.750 46.480 ;
        RECT 171.760 45.800 181.370 46.480 ;
        RECT 176.270 45.580 177.200 45.800 ;
        RECT 180.030 45.570 181.370 45.800 ;
        RECT 181.420 45.800 185.320 46.480 ;
        RECT 181.420 45.570 182.350 45.800 ;
        RECT 185.560 45.670 187.390 46.480 ;
        RECT 187.870 45.610 188.300 46.395 ;
        RECT 189.240 45.800 198.850 46.480 ;
        RECT 199.930 45.800 203.395 46.480 ;
        RECT 193.750 45.580 194.680 45.800 ;
        RECT 197.510 45.570 198.850 45.800 ;
        RECT 202.475 45.570 203.395 45.800 ;
        RECT 203.500 45.800 207.400 46.480 ;
        RECT 203.500 45.570 204.430 45.800 ;
        RECT 207.640 45.670 209.470 46.480 ;
        RECT 209.710 45.800 213.610 46.480 ;
        RECT 212.680 45.570 213.610 45.800 ;
        RECT 213.630 45.610 214.060 46.395 ;
        RECT 214.080 45.670 215.910 46.480 ;
        RECT 216.380 45.800 225.570 46.480 ;
        RECT 220.890 45.580 221.820 45.800 ;
        RECT 224.650 45.570 225.570 45.800 ;
        RECT 226.365 45.570 230.020 46.480 ;
        RECT 230.180 45.800 239.370 46.480 ;
        RECT 234.690 45.580 235.620 45.800 ;
        RECT 238.450 45.570 239.370 45.800 ;
        RECT 239.390 45.610 239.820 46.395 ;
        RECT 239.990 45.570 243.645 46.480 ;
        RECT 244.075 45.800 247.540 46.480 ;
        RECT 248.120 45.800 257.310 46.480 ;
        RECT 244.075 45.570 244.995 45.800 ;
        RECT 252.630 45.580 253.560 45.800 ;
        RECT 256.390 45.570 257.310 45.800 ;
        RECT 257.415 45.800 260.880 46.480 ;
        RECT 257.415 45.570 258.335 45.800 ;
        RECT 261.000 45.570 264.210 46.480 ;
        RECT 265.150 45.610 265.580 46.395 ;
        RECT 265.600 45.800 267.890 46.480 ;
        RECT 266.970 45.570 267.890 45.800 ;
        RECT 267.915 45.800 270.190 46.480 ;
        RECT 267.915 45.570 269.285 45.800 ;
        RECT 270.300 45.570 272.490 46.480 ;
        RECT 272.500 45.670 278.010 46.480 ;
        RECT 278.710 45.800 282.610 46.480 ;
        RECT 282.730 45.800 286.195 46.480 ;
        RECT 281.680 45.570 282.610 45.800 ;
        RECT 285.275 45.570 286.195 45.800 ;
        RECT 286.300 45.670 289.970 46.480 ;
        RECT 290.910 45.610 291.340 46.395 ;
        RECT 291.360 45.800 300.550 46.480 ;
        RECT 291.360 45.570 292.280 45.800 ;
        RECT 295.110 45.580 296.040 45.800 ;
        RECT 300.560 45.670 306.070 46.480 ;
        RECT 306.080 45.670 309.750 46.480 ;
        RECT 309.760 45.670 311.130 46.480 ;
      LAYER nwell ;
        RECT 161.905 42.450 311.325 45.280 ;
      LAYER pwell ;
        RECT 162.100 41.250 163.470 42.060 ;
        RECT 163.480 41.250 165.310 42.060 ;
        RECT 170.290 41.930 171.220 42.150 ;
        RECT 174.050 41.930 174.970 42.160 ;
        RECT 165.780 41.250 174.970 41.930 ;
        RECT 174.990 41.335 175.420 42.120 ;
        RECT 179.950 41.930 180.880 42.150 ;
        RECT 183.710 41.930 184.630 42.160 ;
        RECT 189.150 41.930 190.080 42.150 ;
        RECT 192.910 41.930 194.250 42.160 ;
        RECT 175.440 41.250 184.630 41.930 ;
        RECT 184.640 41.250 194.250 41.930 ;
        RECT 194.300 41.930 195.230 42.160 ;
        RECT 194.300 41.250 198.200 41.930 ;
        RECT 198.440 41.250 200.270 42.060 ;
        RECT 200.750 41.335 201.180 42.120 ;
        RECT 205.710 41.930 206.640 42.150 ;
        RECT 209.470 41.930 210.390 42.160 ;
        RECT 212.245 41.930 213.610 42.160 ;
        RECT 218.130 41.930 219.060 42.150 ;
        RECT 221.890 41.930 222.810 42.160 ;
        RECT 225.475 41.930 226.395 42.160 ;
        RECT 201.200 41.250 210.390 41.930 ;
        RECT 210.400 41.250 213.610 41.930 ;
        RECT 213.620 41.250 222.810 41.930 ;
        RECT 222.930 41.250 226.395 41.930 ;
        RECT 226.510 41.335 226.940 42.120 ;
        RECT 234.690 41.930 235.620 42.150 ;
        RECT 238.450 41.930 239.370 42.160 ;
        RECT 226.970 41.250 229.710 41.930 ;
        RECT 230.180 41.250 239.370 41.930 ;
        RECT 239.705 41.250 243.360 42.160 ;
        RECT 243.615 41.930 244.535 42.160 ;
        RECT 243.615 41.250 247.080 41.930 ;
        RECT 247.200 41.250 248.570 42.060 ;
        RECT 251.235 41.930 252.155 42.160 ;
        RECT 248.690 41.250 252.155 41.930 ;
        RECT 252.270 41.335 252.700 42.120 ;
        RECT 252.720 41.250 255.460 41.930 ;
        RECT 255.480 41.250 257.310 42.060 ;
        RECT 258.090 41.930 259.020 42.160 ;
        RECT 261.130 41.930 262.060 42.160 ;
        RECT 258.090 41.250 259.925 41.930 ;
        RECT 162.240 41.040 162.410 41.250 ;
        RECT 163.620 41.200 163.790 41.250 ;
        RECT 163.615 41.090 163.790 41.200 ;
        RECT 163.620 41.060 163.790 41.090 ;
        RECT 164.080 41.040 164.250 41.230 ;
        RECT 165.455 41.090 165.575 41.200 ;
        RECT 165.920 41.060 166.090 41.250 ;
        RECT 175.580 41.060 175.750 41.250 ;
        RECT 176.500 41.040 176.670 41.230 ;
        RECT 177.235 41.040 177.405 41.230 ;
        RECT 181.100 41.040 181.270 41.230 ;
        RECT 183.855 41.090 183.975 41.200 ;
        RECT 184.780 41.060 184.950 41.250 ;
        RECT 187.540 41.040 187.710 41.230 ;
        RECT 188.735 41.040 188.905 41.230 ;
        RECT 193.980 41.040 194.150 41.230 ;
        RECT 194.440 41.040 194.610 41.230 ;
        RECT 194.715 41.060 194.885 41.250 ;
        RECT 195.820 41.040 195.990 41.230 ;
        RECT 198.580 41.060 198.750 41.250 ;
        RECT 200.415 41.090 200.535 41.200 ;
        RECT 201.340 41.060 201.510 41.250 ;
        RECT 208.240 41.040 208.410 41.230 ;
        RECT 208.700 41.040 208.870 41.230 ;
        RECT 210.545 41.060 210.715 41.250 ;
        RECT 213.300 41.040 213.470 41.230 ;
        RECT 213.760 41.060 213.930 41.250 ;
        RECT 222.960 41.040 223.130 41.250 ;
        RECT 223.420 41.040 223.590 41.230 ;
        RECT 228.665 41.040 228.835 41.230 ;
        RECT 229.400 41.060 229.570 41.250 ;
        RECT 229.675 41.040 229.845 41.230 ;
        RECT 229.855 41.090 229.975 41.200 ;
        RECT 230.320 41.060 230.490 41.250 ;
        RECT 243.200 41.230 243.360 41.250 ;
        RECT 233.535 41.090 233.655 41.200 ;
        RECT 234.275 41.040 234.445 41.230 ;
        RECT 238.140 41.040 238.310 41.230 ;
        RECT 241.820 41.060 241.990 41.230 ;
        RECT 241.820 41.040 241.985 41.060 ;
        RECT 242.555 41.040 242.725 41.230 ;
        RECT 243.200 41.060 243.370 41.230 ;
        RECT 246.695 41.040 246.865 41.230 ;
        RECT 246.880 41.060 247.050 41.250 ;
        RECT 247.340 41.060 247.510 41.250 ;
        RECT 248.720 41.060 248.890 41.250 ;
        RECT 252.860 41.060 253.030 41.250 ;
        RECT 253.780 41.040 253.950 41.230 ;
        RECT 254.240 41.040 254.410 41.230 ;
        RECT 255.620 41.060 255.790 41.250 ;
        RECT 259.760 41.230 259.925 41.250 ;
        RECT 260.225 41.250 262.060 41.930 ;
        RECT 262.380 41.250 264.210 42.060 ;
        RECT 264.230 41.250 265.580 42.160 ;
        RECT 265.600 41.250 266.970 42.060 ;
        RECT 271.490 41.930 272.420 42.150 ;
        RECT 275.250 41.930 276.170 42.160 ;
        RECT 266.980 41.250 276.170 41.930 ;
        RECT 276.180 41.250 278.010 42.160 ;
        RECT 278.030 41.335 278.460 42.120 ;
        RECT 278.480 41.250 280.295 42.160 ;
        RECT 280.875 41.930 281.795 42.160 ;
        RECT 280.875 41.250 284.340 41.930 ;
        RECT 284.470 41.250 285.820 42.160 ;
        RECT 285.935 41.930 286.855 42.160 ;
        RECT 285.935 41.250 289.400 41.930 ;
        RECT 289.520 41.250 295.030 42.060 ;
        RECT 295.040 41.250 300.550 42.060 ;
        RECT 300.560 41.250 303.310 42.060 ;
        RECT 303.790 41.335 304.220 42.120 ;
        RECT 304.240 41.250 306.070 42.060 ;
        RECT 306.565 41.930 307.910 42.160 ;
        RECT 306.080 41.250 307.910 41.930 ;
        RECT 307.920 41.250 309.750 42.060 ;
        RECT 309.760 41.250 311.130 42.060 ;
        RECT 260.225 41.230 260.390 41.250 ;
        RECT 256.075 41.090 256.195 41.200 ;
        RECT 257.455 41.040 257.625 41.230 ;
        RECT 257.925 41.040 258.095 41.230 ;
        RECT 259.760 41.060 259.930 41.230 ;
        RECT 260.220 41.060 260.390 41.230 ;
        RECT 262.060 41.040 262.230 41.230 ;
        RECT 262.520 41.060 262.690 41.250 ;
        RECT 264.360 41.060 264.530 41.250 ;
        RECT 264.815 41.090 264.935 41.200 ;
        RECT 265.740 41.060 265.910 41.250 ;
        RECT 267.120 41.060 267.290 41.250 ;
        RECT 268.960 41.040 269.130 41.230 ;
        RECT 269.430 41.085 269.590 41.195 ;
        RECT 271.715 41.040 271.885 41.230 ;
        RECT 277.695 41.060 277.865 41.250 ;
        RECT 280.000 41.060 280.170 41.250 ;
        RECT 280.455 41.090 280.575 41.200 ;
        RECT 280.920 41.040 281.090 41.230 ;
        RECT 284.140 41.060 284.310 41.250 ;
        RECT 284.600 41.060 284.770 41.250 ;
        RECT 289.200 41.060 289.370 41.250 ;
        RECT 289.660 41.060 289.830 41.250 ;
        RECT 290.120 41.040 290.290 41.230 ;
        RECT 290.575 41.090 290.695 41.200 ;
        RECT 291.500 41.040 291.670 41.230 ;
        RECT 295.180 41.060 295.350 41.250 ;
        RECT 297.030 41.085 297.190 41.195 ;
        RECT 297.940 41.040 298.110 41.230 ;
        RECT 300.700 41.060 300.870 41.250 ;
        RECT 303.455 41.090 303.575 41.200 ;
        RECT 304.380 41.060 304.550 41.250 ;
        RECT 306.220 41.060 306.390 41.250 ;
        RECT 307.140 41.040 307.310 41.230 ;
        RECT 308.060 41.060 308.230 41.250 ;
        RECT 308.990 41.085 309.150 41.195 ;
        RECT 310.820 41.040 310.990 41.250 ;
        RECT 162.100 40.230 163.470 41.040 ;
        RECT 164.050 40.360 167.515 41.040 ;
        RECT 166.595 40.130 167.515 40.360 ;
        RECT 167.620 40.360 176.810 41.040 ;
        RECT 176.820 40.360 180.720 41.040 ;
        RECT 167.620 40.130 168.540 40.360 ;
        RECT 171.370 40.140 172.300 40.360 ;
        RECT 176.820 40.130 177.750 40.360 ;
        RECT 180.960 40.230 183.710 41.040 ;
        RECT 184.275 40.360 187.740 41.040 ;
        RECT 184.275 40.130 185.195 40.360 ;
        RECT 187.870 40.170 188.300 40.955 ;
        RECT 188.320 40.360 192.220 41.040 ;
        RECT 192.460 40.360 194.290 41.040 ;
        RECT 188.320 40.130 189.250 40.360 ;
        RECT 194.300 40.230 195.670 41.040 ;
        RECT 195.680 40.360 204.870 41.040 ;
        RECT 200.190 40.140 201.120 40.360 ;
        RECT 203.950 40.130 204.870 40.360 ;
        RECT 204.975 40.360 208.440 41.040 ;
        RECT 204.975 40.130 205.895 40.360 ;
        RECT 208.560 40.230 209.930 41.040 ;
        RECT 210.035 40.360 213.500 41.040 ;
        RECT 210.035 40.130 210.955 40.360 ;
        RECT 213.630 40.170 214.060 40.955 ;
        RECT 214.080 40.360 223.270 41.040 ;
        RECT 214.080 40.130 215.000 40.360 ;
        RECT 217.830 40.140 218.760 40.360 ;
        RECT 223.280 40.230 225.110 41.040 ;
        RECT 225.350 40.360 229.250 41.040 ;
        RECT 228.320 40.130 229.250 40.360 ;
        RECT 229.260 40.360 233.160 41.040 ;
        RECT 233.860 40.360 237.760 41.040 ;
        RECT 229.260 40.130 230.190 40.360 ;
        RECT 233.860 40.130 234.790 40.360 ;
        RECT 238.000 40.230 239.370 41.040 ;
        RECT 239.390 40.170 239.820 40.955 ;
        RECT 240.150 40.360 241.985 41.040 ;
        RECT 242.140 40.360 246.040 41.040 ;
        RECT 246.280 40.360 250.180 41.040 ;
        RECT 250.515 40.360 253.980 41.040 ;
        RECT 240.150 40.130 241.080 40.360 ;
        RECT 242.140 40.130 243.070 40.360 ;
        RECT 246.280 40.130 247.210 40.360 ;
        RECT 250.515 40.130 251.435 40.360 ;
        RECT 254.100 40.230 255.930 41.040 ;
        RECT 256.420 40.130 257.770 41.040 ;
        RECT 257.780 40.130 261.670 41.040 ;
        RECT 261.920 40.130 264.670 41.040 ;
        RECT 265.150 40.170 265.580 40.955 ;
        RECT 265.695 40.360 269.160 41.040 ;
        RECT 265.695 40.130 266.615 40.360 ;
        RECT 270.260 40.130 272.030 41.040 ;
        RECT 272.040 40.360 281.230 41.040 ;
        RECT 281.240 40.360 290.430 41.040 ;
        RECT 272.040 40.130 272.960 40.360 ;
        RECT 275.790 40.140 276.720 40.360 ;
        RECT 281.240 40.130 282.160 40.360 ;
        RECT 284.990 40.140 285.920 40.360 ;
        RECT 290.910 40.170 291.340 40.955 ;
        RECT 291.360 40.230 296.870 41.040 ;
        RECT 297.800 40.360 306.990 41.040 ;
        RECT 307.000 40.360 308.830 41.040 ;
        RECT 302.310 40.140 303.240 40.360 ;
        RECT 306.070 40.130 306.990 40.360 ;
        RECT 307.485 40.130 308.830 40.360 ;
        RECT 309.760 40.230 311.130 41.040 ;
      LAYER nwell ;
        RECT 161.905 37.010 311.325 39.840 ;
      LAYER pwell ;
        RECT 162.100 35.810 163.470 36.620 ;
        RECT 163.480 35.810 167.150 36.620 ;
        RECT 170.275 36.490 171.195 36.720 ;
        RECT 173.955 36.490 174.875 36.720 ;
        RECT 167.730 35.810 171.195 36.490 ;
        RECT 171.410 35.810 174.875 36.490 ;
        RECT 174.990 35.895 175.420 36.680 ;
        RECT 175.440 36.490 176.370 36.720 ;
        RECT 175.440 35.810 179.340 36.490 ;
        RECT 179.580 35.810 181.410 36.620 ;
        RECT 184.535 36.490 185.455 36.720 ;
        RECT 181.990 35.810 185.455 36.490 ;
        RECT 185.560 36.490 186.480 36.720 ;
        RECT 189.310 36.490 190.240 36.710 ;
        RECT 197.415 36.490 198.335 36.720 ;
        RECT 185.560 35.810 194.750 36.490 ;
        RECT 194.870 35.810 198.335 36.490 ;
        RECT 198.440 35.810 200.270 36.620 ;
        RECT 200.750 35.895 201.180 36.680 ;
        RECT 201.200 35.810 203.030 36.620 ;
        RECT 203.500 36.490 204.430 36.720 ;
        RECT 207.735 36.490 208.655 36.720 ;
        RECT 217.740 36.490 218.670 36.720 ;
        RECT 221.795 36.490 222.715 36.720 ;
        RECT 225.475 36.490 226.395 36.720 ;
        RECT 203.500 35.810 207.400 36.490 ;
        RECT 207.735 35.810 211.200 36.490 ;
        RECT 211.330 35.810 214.070 36.490 ;
        RECT 214.770 35.810 218.670 36.490 ;
        RECT 219.250 35.810 222.715 36.490 ;
        RECT 222.930 35.810 226.395 36.490 ;
        RECT 226.510 35.895 226.940 36.680 ;
        RECT 226.960 35.810 229.710 36.620 ;
        RECT 234.690 36.490 235.620 36.710 ;
        RECT 238.450 36.490 239.790 36.720 ;
        RECT 245.270 36.490 246.200 36.710 ;
        RECT 249.030 36.490 249.950 36.720 ;
        RECT 230.180 35.810 239.790 36.490 ;
        RECT 240.760 35.810 249.950 36.490 ;
        RECT 249.960 35.810 251.790 36.620 ;
        RECT 252.270 35.895 252.700 36.680 ;
        RECT 252.720 35.810 254.550 36.620 ;
        RECT 255.020 36.490 255.940 36.720 ;
        RECT 258.770 36.490 259.700 36.710 ;
        RECT 266.980 36.490 267.900 36.720 ;
        RECT 255.020 35.810 264.210 36.490 ;
        RECT 264.220 35.810 266.960 36.490 ;
        RECT 266.980 35.810 269.270 36.490 ;
        RECT 269.280 35.810 272.950 36.620 ;
        RECT 274.015 36.490 277.525 36.720 ;
        RECT 274.015 35.810 278.010 36.490 ;
        RECT 278.030 35.895 278.460 36.680 ;
        RECT 278.575 36.490 279.495 36.720 ;
        RECT 282.160 36.520 283.110 36.720 ;
        RECT 284.440 36.520 285.370 36.720 ;
        RECT 278.575 35.810 282.040 36.490 ;
        RECT 282.160 36.040 285.370 36.520 ;
        RECT 282.160 35.840 285.225 36.040 ;
        RECT 282.160 35.810 283.095 35.840 ;
        RECT 162.240 35.600 162.410 35.810 ;
        RECT 163.620 35.600 163.790 35.810 ;
        RECT 165.455 35.650 165.575 35.760 ;
        RECT 167.295 35.650 167.415 35.760 ;
        RECT 167.760 35.620 167.930 35.810 ;
        RECT 171.440 35.620 171.610 35.810 ;
        RECT 174.660 35.600 174.830 35.790 ;
        RECT 175.395 35.600 175.565 35.790 ;
        RECT 175.855 35.620 176.025 35.810 ;
        RECT 179.255 35.650 179.375 35.760 ;
        RECT 179.720 35.620 179.890 35.810 ;
        RECT 181.555 35.650 181.675 35.760 ;
        RECT 182.020 35.620 182.190 35.810 ;
        RECT 183.125 35.600 183.295 35.790 ;
        RECT 187.265 35.600 187.435 35.790 ;
        RECT 194.440 35.620 194.610 35.810 ;
        RECT 194.900 35.620 195.070 35.810 ;
        RECT 197.200 35.600 197.370 35.790 ;
        RECT 197.660 35.600 197.830 35.790 ;
        RECT 198.580 35.620 198.750 35.810 ;
        RECT 200.420 35.760 200.590 35.790 ;
        RECT 200.415 35.650 200.590 35.760 ;
        RECT 200.420 35.600 200.590 35.650 ;
        RECT 201.340 35.620 201.510 35.810 ;
        RECT 203.175 35.650 203.295 35.760 ;
        RECT 203.915 35.620 204.085 35.810 ;
        RECT 209.615 35.650 209.735 35.760 ;
        RECT 210.080 35.600 210.250 35.790 ;
        RECT 211.000 35.620 211.170 35.810 ;
        RECT 213.760 35.620 213.930 35.810 ;
        RECT 214.215 35.650 214.335 35.760 ;
        RECT 214.495 35.600 214.665 35.790 ;
        RECT 218.085 35.620 218.255 35.810 ;
        RECT 218.815 35.650 218.935 35.760 ;
        RECT 219.280 35.620 219.450 35.810 ;
        RECT 222.960 35.620 223.130 35.810 ;
        RECT 227.100 35.600 227.270 35.810 ;
        RECT 227.560 35.600 227.730 35.790 ;
        RECT 229.400 35.600 229.570 35.790 ;
        RECT 229.855 35.650 229.975 35.760 ;
        RECT 230.320 35.620 230.490 35.810 ;
        RECT 239.990 35.760 240.150 35.765 ;
        RECT 238.610 35.645 238.770 35.755 ;
        RECT 239.975 35.655 240.150 35.760 ;
        RECT 239.975 35.650 240.095 35.655 ;
        RECT 240.440 35.600 240.610 35.790 ;
        RECT 240.900 35.620 241.070 35.810 ;
        RECT 249.640 35.600 249.810 35.790 ;
        RECT 250.100 35.620 250.270 35.810 ;
        RECT 251.935 35.650 252.055 35.760 ;
        RECT 252.860 35.620 253.030 35.810 ;
        RECT 254.695 35.650 254.815 35.760 ;
        RECT 255.155 35.650 255.275 35.760 ;
        RECT 255.620 35.600 255.790 35.790 ;
        RECT 263.900 35.620 264.070 35.810 ;
        RECT 264.360 35.620 264.530 35.810 ;
        RECT 264.815 35.650 264.935 35.760 ;
        RECT 267.580 35.620 267.750 35.790 ;
        RECT 267.580 35.600 267.730 35.620 ;
        RECT 268.040 35.600 268.210 35.790 ;
        RECT 268.960 35.620 269.130 35.810 ;
        RECT 269.420 35.620 269.590 35.810 ;
        RECT 273.110 35.655 273.270 35.765 ;
        RECT 273.560 35.600 273.730 35.790 ;
        RECT 277.695 35.620 277.865 35.810 ;
        RECT 279.080 35.600 279.250 35.790 ;
        RECT 281.840 35.620 282.010 35.810 ;
        RECT 284.600 35.600 284.770 35.790 ;
        RECT 285.055 35.620 285.225 35.840 ;
        RECT 285.380 35.810 290.890 36.620 ;
        RECT 290.900 35.810 296.410 36.620 ;
        RECT 296.420 35.810 301.930 36.620 ;
        RECT 301.940 35.810 303.770 36.620 ;
        RECT 303.790 35.895 304.220 36.680 ;
        RECT 304.700 35.810 306.070 36.590 ;
        RECT 308.735 36.490 309.655 36.720 ;
        RECT 306.190 35.810 309.655 36.490 ;
        RECT 309.760 35.810 311.130 36.620 ;
        RECT 285.520 35.620 285.690 35.810 ;
        RECT 290.130 35.645 290.290 35.755 ;
        RECT 291.040 35.620 291.210 35.810 ;
        RECT 291.500 35.600 291.670 35.790 ;
        RECT 296.560 35.620 296.730 35.810 ;
        RECT 297.020 35.600 297.190 35.790 ;
        RECT 302.080 35.620 302.250 35.810 ;
        RECT 304.375 35.650 304.495 35.760 ;
        RECT 304.840 35.620 305.010 35.810 ;
        RECT 306.220 35.620 306.390 35.810 ;
        RECT 308.520 35.600 308.690 35.790 ;
        RECT 308.990 35.645 309.150 35.755 ;
        RECT 310.820 35.600 310.990 35.810 ;
        RECT 162.100 34.790 163.470 35.600 ;
        RECT 163.480 34.790 165.310 35.600 ;
        RECT 165.780 34.920 174.970 35.600 ;
        RECT 174.980 34.920 178.880 35.600 ;
        RECT 179.810 34.920 183.710 35.600 ;
        RECT 183.950 34.920 187.850 35.600 ;
        RECT 165.780 34.690 166.700 34.920 ;
        RECT 169.530 34.700 170.460 34.920 ;
        RECT 174.980 34.690 175.910 34.920 ;
        RECT 182.780 34.690 183.710 34.920 ;
        RECT 186.920 34.690 187.850 34.920 ;
        RECT 187.870 34.730 188.300 35.515 ;
        RECT 188.320 34.920 197.510 35.600 ;
        RECT 188.320 34.690 189.240 34.920 ;
        RECT 192.070 34.700 193.000 34.920 ;
        RECT 197.520 34.790 200.270 35.600 ;
        RECT 200.280 34.920 209.470 35.600 ;
        RECT 210.050 34.920 213.515 35.600 ;
        RECT 204.790 34.700 205.720 34.920 ;
        RECT 208.550 34.690 209.470 34.920 ;
        RECT 212.595 34.690 213.515 34.920 ;
        RECT 213.630 34.730 214.060 35.515 ;
        RECT 214.080 34.920 217.980 35.600 ;
        RECT 218.220 34.920 227.410 35.600 ;
        RECT 214.080 34.690 215.010 34.920 ;
        RECT 218.220 34.690 219.140 34.920 ;
        RECT 221.970 34.700 222.900 34.920 ;
        RECT 227.420 34.790 229.250 35.600 ;
        RECT 229.260 34.920 238.450 35.600 ;
        RECT 233.770 34.700 234.700 34.920 ;
        RECT 237.530 34.690 238.450 34.920 ;
        RECT 239.390 34.730 239.820 35.515 ;
        RECT 240.300 34.920 249.490 35.600 ;
        RECT 244.810 34.700 245.740 34.920 ;
        RECT 248.570 34.690 249.490 34.920 ;
        RECT 249.500 34.790 255.010 35.600 ;
        RECT 255.480 34.920 264.670 35.600 ;
        RECT 259.990 34.700 260.920 34.920 ;
        RECT 263.750 34.690 264.670 34.920 ;
        RECT 265.150 34.730 265.580 35.515 ;
        RECT 265.800 34.780 267.730 35.600 ;
        RECT 267.900 34.790 273.410 35.600 ;
        RECT 273.420 34.790 278.930 35.600 ;
        RECT 278.940 34.790 284.450 35.600 ;
        RECT 284.460 34.790 289.970 35.600 ;
        RECT 265.800 34.690 266.750 34.780 ;
        RECT 290.910 34.730 291.340 35.515 ;
        RECT 291.360 34.790 296.870 35.600 ;
        RECT 296.880 34.790 299.630 35.600 ;
        RECT 299.640 34.920 308.830 35.600 ;
        RECT 299.640 34.690 300.560 34.920 ;
        RECT 303.390 34.700 304.320 34.920 ;
        RECT 309.760 34.790 311.130 35.600 ;
      LAYER nwell ;
        RECT 161.905 31.570 311.325 34.400 ;
      LAYER pwell ;
        RECT 162.100 30.370 163.470 31.180 ;
        RECT 163.480 30.370 165.310 31.180 ;
        RECT 170.290 31.050 171.220 31.270 ;
        RECT 174.050 31.050 174.970 31.280 ;
        RECT 165.780 30.370 174.970 31.050 ;
        RECT 174.990 30.455 175.420 31.240 ;
        RECT 175.440 31.050 176.370 31.280 ;
        RECT 175.440 30.370 179.340 31.050 ;
        RECT 179.580 30.370 181.410 31.180 ;
        RECT 181.880 31.050 182.800 31.280 ;
        RECT 185.630 31.050 186.560 31.270 ;
        RECT 191.080 31.050 192.010 31.280 ;
        RECT 181.880 30.370 191.070 31.050 ;
        RECT 191.080 30.370 194.980 31.050 ;
        RECT 195.220 30.370 197.970 31.180 ;
        RECT 197.990 30.370 200.730 31.050 ;
        RECT 200.750 30.455 201.180 31.240 ;
        RECT 201.200 31.050 202.130 31.280 ;
        RECT 206.260 31.050 207.180 31.280 ;
        RECT 210.010 31.050 210.940 31.270 ;
        RECT 201.200 30.370 205.100 31.050 ;
        RECT 206.260 30.370 215.450 31.050 ;
        RECT 215.460 30.370 217.290 31.180 ;
        RECT 219.955 31.050 220.875 31.280 ;
        RECT 217.410 30.370 220.875 31.050 ;
        RECT 220.980 30.370 222.350 31.180 ;
        RECT 222.360 31.050 223.290 31.280 ;
        RECT 222.360 30.370 226.260 31.050 ;
        RECT 226.510 30.455 226.940 31.240 ;
        RECT 231.470 31.050 232.400 31.270 ;
        RECT 235.230 31.050 236.150 31.280 ;
        RECT 226.960 30.370 236.150 31.050 ;
        RECT 236.255 31.050 237.175 31.280 ;
        RECT 236.255 30.370 239.720 31.050 ;
        RECT 239.850 30.370 242.590 31.050 ;
        RECT 242.600 30.370 244.430 31.050 ;
        RECT 244.440 30.370 249.950 31.180 ;
        RECT 249.960 30.370 251.790 31.180 ;
        RECT 252.270 30.455 252.700 31.240 ;
        RECT 252.720 30.370 258.230 31.180 ;
        RECT 258.240 30.370 260.070 31.180 ;
        RECT 260.100 30.370 261.450 31.280 ;
        RECT 261.460 30.370 266.970 31.180 ;
        RECT 266.980 30.370 272.490 31.180 ;
        RECT 272.500 30.370 278.010 31.180 ;
        RECT 278.030 30.455 278.460 31.240 ;
        RECT 278.480 30.370 283.990 31.180 ;
        RECT 284.000 30.370 289.510 31.180 ;
        RECT 289.520 30.370 295.030 31.180 ;
        RECT 295.040 30.370 300.550 31.180 ;
        RECT 300.560 30.370 303.310 31.180 ;
        RECT 303.790 30.455 304.220 31.240 ;
        RECT 304.240 30.370 309.750 31.180 ;
        RECT 309.760 30.370 311.130 31.180 ;
        RECT 162.240 30.160 162.410 30.370 ;
        RECT 163.620 30.180 163.790 30.370 ;
        RECT 165.000 30.160 165.170 30.350 ;
        RECT 165.460 30.320 165.630 30.350 ;
        RECT 165.455 30.210 165.630 30.320 ;
        RECT 165.460 30.160 165.630 30.210 ;
        RECT 165.920 30.180 166.090 30.370 ;
        RECT 170.980 30.160 171.150 30.350 ;
        RECT 174.655 30.210 174.775 30.320 ;
        RECT 175.120 30.160 175.290 30.350 ;
        RECT 175.855 30.180 176.025 30.370 ;
        RECT 179.720 30.180 179.890 30.370 ;
        RECT 181.555 30.210 181.675 30.320 ;
        RECT 187.540 30.160 187.710 30.350 ;
        RECT 188.460 30.160 188.630 30.350 ;
        RECT 190.760 30.180 190.930 30.370 ;
        RECT 191.495 30.180 191.665 30.370 ;
        RECT 193.980 30.160 194.150 30.350 ;
        RECT 195.360 30.180 195.530 30.370 ;
        RECT 200.420 30.180 200.590 30.370 ;
        RECT 201.615 30.180 201.785 30.370 ;
        RECT 204.560 30.160 204.730 30.350 ;
        RECT 205.490 30.215 205.650 30.325 ;
        RECT 208.240 30.160 208.410 30.350 ;
        RECT 208.700 30.160 208.870 30.350 ;
        RECT 212.380 30.160 212.550 30.350 ;
        RECT 214.220 30.160 214.390 30.350 ;
        RECT 215.140 30.180 215.310 30.370 ;
        RECT 215.600 30.180 215.770 30.370 ;
        RECT 217.440 30.180 217.610 30.370 ;
        RECT 219.740 30.160 219.910 30.350 ;
        RECT 221.120 30.180 221.290 30.370 ;
        RECT 222.775 30.180 222.945 30.370 ;
        RECT 225.260 30.160 225.430 30.350 ;
        RECT 227.100 30.180 227.270 30.370 ;
        RECT 230.790 30.205 230.950 30.315 ;
        RECT 234.920 30.160 235.090 30.350 ;
        RECT 235.380 30.160 235.550 30.350 ;
        RECT 239.055 30.210 239.175 30.320 ;
        RECT 239.520 30.180 239.690 30.370 ;
        RECT 239.980 30.160 240.150 30.350 ;
        RECT 242.280 30.180 242.450 30.370 ;
        RECT 244.120 30.180 244.290 30.370 ;
        RECT 244.580 30.180 244.750 30.370 ;
        RECT 245.500 30.160 245.670 30.350 ;
        RECT 250.100 30.180 250.270 30.370 ;
        RECT 251.020 30.160 251.190 30.350 ;
        RECT 251.935 30.210 252.055 30.320 ;
        RECT 252.860 30.180 253.030 30.370 ;
        RECT 256.540 30.160 256.710 30.350 ;
        RECT 258.380 30.180 258.550 30.370 ;
        RECT 260.215 30.180 260.385 30.370 ;
        RECT 261.600 30.180 261.770 30.370 ;
        RECT 262.060 30.160 262.230 30.350 ;
        RECT 264.815 30.210 264.935 30.320 ;
        RECT 265.740 30.160 265.910 30.350 ;
        RECT 267.120 30.180 267.290 30.370 ;
        RECT 271.260 30.160 271.430 30.350 ;
        RECT 272.640 30.180 272.810 30.370 ;
        RECT 276.780 30.160 276.950 30.350 ;
        RECT 278.620 30.180 278.790 30.370 ;
        RECT 282.300 30.160 282.470 30.350 ;
        RECT 284.140 30.180 284.310 30.370 ;
        RECT 287.820 30.160 287.990 30.350 ;
        RECT 289.660 30.180 289.830 30.370 ;
        RECT 290.575 30.210 290.695 30.320 ;
        RECT 291.500 30.160 291.670 30.350 ;
        RECT 295.180 30.180 295.350 30.370 ;
        RECT 297.020 30.160 297.190 30.350 ;
        RECT 300.700 30.180 300.870 30.370 ;
        RECT 302.540 30.160 302.710 30.350 ;
        RECT 303.455 30.210 303.575 30.320 ;
        RECT 304.380 30.180 304.550 30.370 ;
        RECT 308.060 30.160 308.230 30.350 ;
        RECT 310.820 30.160 310.990 30.370 ;
        RECT 162.100 29.350 163.470 30.160 ;
        RECT 163.480 29.480 165.310 30.160 ;
        RECT 163.480 29.250 164.825 29.480 ;
        RECT 165.320 29.350 170.830 30.160 ;
        RECT 170.840 29.350 174.510 30.160 ;
        RECT 175.090 29.480 178.555 30.160 ;
        RECT 177.635 29.250 178.555 29.480 ;
        RECT 178.660 29.480 187.850 30.160 ;
        RECT 178.660 29.250 179.580 29.480 ;
        RECT 182.410 29.260 183.340 29.480 ;
        RECT 187.870 29.290 188.300 30.075 ;
        RECT 188.320 29.350 193.830 30.160 ;
        RECT 193.840 29.350 195.670 30.160 ;
        RECT 195.680 29.480 204.870 30.160 ;
        RECT 204.975 29.480 208.440 30.160 ;
        RECT 195.680 29.250 196.600 29.480 ;
        RECT 199.430 29.260 200.360 29.480 ;
        RECT 204.975 29.250 205.895 29.480 ;
        RECT 208.560 29.350 212.230 30.160 ;
        RECT 212.240 29.350 213.610 30.160 ;
        RECT 213.630 29.290 214.060 30.075 ;
        RECT 214.080 29.350 219.590 30.160 ;
        RECT 219.600 29.350 225.110 30.160 ;
        RECT 225.120 29.350 230.630 30.160 ;
        RECT 231.655 29.480 235.120 30.160 ;
        RECT 231.655 29.250 232.575 29.480 ;
        RECT 235.240 29.350 238.910 30.160 ;
        RECT 239.390 29.290 239.820 30.075 ;
        RECT 239.840 29.350 245.350 30.160 ;
        RECT 245.360 29.350 250.870 30.160 ;
        RECT 250.880 29.350 256.390 30.160 ;
        RECT 256.400 29.350 261.910 30.160 ;
        RECT 261.920 29.350 264.670 30.160 ;
        RECT 265.150 29.290 265.580 30.075 ;
        RECT 265.600 29.350 271.110 30.160 ;
        RECT 271.120 29.350 276.630 30.160 ;
        RECT 276.640 29.350 282.150 30.160 ;
        RECT 282.160 29.350 287.670 30.160 ;
        RECT 287.680 29.350 290.430 30.160 ;
        RECT 290.910 29.290 291.340 30.075 ;
        RECT 291.360 29.350 296.870 30.160 ;
        RECT 296.880 29.350 302.390 30.160 ;
        RECT 302.400 29.350 307.910 30.160 ;
        RECT 307.920 29.350 309.750 30.160 ;
        RECT 309.760 29.350 311.130 30.160 ;
      LAYER nwell ;
        RECT 161.905 26.130 311.325 28.960 ;
      LAYER pwell ;
        RECT 162.100 24.930 163.470 25.740 ;
        RECT 163.480 24.930 168.990 25.740 ;
        RECT 169.000 24.930 174.510 25.740 ;
        RECT 174.990 25.015 175.420 25.800 ;
        RECT 175.440 24.930 178.190 25.740 ;
        RECT 178.295 25.610 179.215 25.840 ;
        RECT 178.295 24.930 181.760 25.610 ;
        RECT 181.880 24.930 183.250 25.740 ;
        RECT 185.915 25.610 186.835 25.840 ;
        RECT 183.370 24.930 186.835 25.610 ;
        RECT 186.940 24.930 192.450 25.740 ;
        RECT 192.460 24.930 197.970 25.740 ;
        RECT 197.980 24.930 200.730 25.740 ;
        RECT 200.750 25.015 201.180 25.800 ;
        RECT 201.200 24.930 206.710 25.740 ;
        RECT 206.720 24.930 212.230 25.740 ;
        RECT 212.240 24.930 217.750 25.740 ;
        RECT 217.760 24.930 223.270 25.740 ;
        RECT 223.280 24.930 226.030 25.740 ;
        RECT 226.510 25.015 226.940 25.800 ;
        RECT 226.960 24.930 232.470 25.740 ;
        RECT 232.480 24.930 237.990 25.740 ;
        RECT 238.000 24.930 243.510 25.740 ;
        RECT 243.520 24.930 249.030 25.740 ;
        RECT 249.040 24.930 251.790 25.740 ;
        RECT 252.270 25.015 252.700 25.800 ;
        RECT 252.720 24.930 258.230 25.740 ;
        RECT 258.240 24.930 263.750 25.740 ;
        RECT 263.760 24.930 269.270 25.740 ;
        RECT 269.280 24.930 274.790 25.740 ;
        RECT 274.800 24.930 277.550 25.740 ;
        RECT 278.030 25.015 278.460 25.800 ;
        RECT 278.480 24.930 283.990 25.740 ;
        RECT 284.000 24.930 289.510 25.740 ;
        RECT 289.520 24.930 295.030 25.740 ;
        RECT 295.040 24.930 300.550 25.740 ;
        RECT 300.560 24.930 303.310 25.740 ;
        RECT 303.790 25.015 304.220 25.800 ;
        RECT 304.240 24.930 309.750 25.740 ;
        RECT 309.760 24.930 311.130 25.740 ;
        RECT 162.240 24.720 162.410 24.930 ;
        RECT 163.620 24.720 163.790 24.930 ;
        RECT 169.140 24.720 169.310 24.930 ;
        RECT 174.660 24.880 174.830 24.910 ;
        RECT 174.655 24.770 174.830 24.880 ;
        RECT 174.660 24.720 174.830 24.770 ;
        RECT 175.580 24.740 175.750 24.930 ;
        RECT 180.180 24.720 180.350 24.910 ;
        RECT 181.560 24.740 181.730 24.930 ;
        RECT 182.020 24.740 182.190 24.930 ;
        RECT 183.400 24.740 183.570 24.930 ;
        RECT 185.700 24.720 185.870 24.910 ;
        RECT 187.080 24.740 187.250 24.930 ;
        RECT 187.535 24.770 187.655 24.880 ;
        RECT 188.460 24.720 188.630 24.910 ;
        RECT 192.600 24.740 192.770 24.930 ;
        RECT 193.980 24.720 194.150 24.910 ;
        RECT 198.120 24.740 198.290 24.930 ;
        RECT 199.500 24.720 199.670 24.910 ;
        RECT 201.340 24.740 201.510 24.930 ;
        RECT 205.020 24.720 205.190 24.910 ;
        RECT 206.860 24.740 207.030 24.930 ;
        RECT 210.540 24.720 210.710 24.910 ;
        RECT 212.380 24.740 212.550 24.930 ;
        RECT 213.295 24.770 213.415 24.880 ;
        RECT 214.220 24.720 214.390 24.910 ;
        RECT 217.900 24.740 218.070 24.930 ;
        RECT 219.740 24.720 219.910 24.910 ;
        RECT 223.420 24.740 223.590 24.930 ;
        RECT 225.260 24.720 225.430 24.910 ;
        RECT 226.175 24.770 226.295 24.880 ;
        RECT 227.100 24.740 227.270 24.930 ;
        RECT 230.780 24.720 230.950 24.910 ;
        RECT 232.620 24.740 232.790 24.930 ;
        RECT 236.300 24.720 236.470 24.910 ;
        RECT 238.140 24.740 238.310 24.930 ;
        RECT 239.055 24.770 239.175 24.880 ;
        RECT 239.980 24.720 240.150 24.910 ;
        RECT 243.660 24.740 243.830 24.930 ;
        RECT 245.500 24.720 245.670 24.910 ;
        RECT 249.180 24.740 249.350 24.930 ;
        RECT 251.020 24.720 251.190 24.910 ;
        RECT 251.935 24.770 252.055 24.880 ;
        RECT 252.860 24.740 253.030 24.930 ;
        RECT 256.540 24.720 256.710 24.910 ;
        RECT 258.380 24.740 258.550 24.930 ;
        RECT 262.060 24.720 262.230 24.910 ;
        RECT 263.900 24.740 264.070 24.930 ;
        RECT 264.815 24.770 264.935 24.880 ;
        RECT 265.740 24.720 265.910 24.910 ;
        RECT 269.420 24.740 269.590 24.930 ;
        RECT 271.260 24.720 271.430 24.910 ;
        RECT 274.940 24.740 275.110 24.930 ;
        RECT 276.780 24.720 276.950 24.910 ;
        RECT 277.695 24.770 277.815 24.880 ;
        RECT 278.620 24.740 278.790 24.930 ;
        RECT 282.300 24.720 282.470 24.910 ;
        RECT 284.140 24.740 284.310 24.930 ;
        RECT 287.820 24.720 287.990 24.910 ;
        RECT 289.660 24.740 289.830 24.930 ;
        RECT 290.575 24.770 290.695 24.880 ;
        RECT 291.500 24.720 291.670 24.910 ;
        RECT 295.180 24.740 295.350 24.930 ;
        RECT 297.020 24.720 297.190 24.910 ;
        RECT 300.700 24.740 300.870 24.930 ;
        RECT 302.540 24.720 302.710 24.910 ;
        RECT 303.455 24.770 303.575 24.880 ;
        RECT 304.380 24.740 304.550 24.930 ;
        RECT 308.060 24.720 308.230 24.910 ;
        RECT 310.820 24.720 310.990 24.930 ;
        RECT 162.100 23.910 163.470 24.720 ;
        RECT 163.480 23.910 168.990 24.720 ;
        RECT 169.000 23.910 174.510 24.720 ;
        RECT 174.520 23.910 180.030 24.720 ;
        RECT 180.040 23.910 185.550 24.720 ;
        RECT 185.560 23.910 187.390 24.720 ;
        RECT 187.870 23.850 188.300 24.635 ;
        RECT 188.320 23.910 193.830 24.720 ;
        RECT 193.840 23.910 199.350 24.720 ;
        RECT 199.360 23.910 204.870 24.720 ;
        RECT 204.880 23.910 210.390 24.720 ;
        RECT 210.400 23.910 213.150 24.720 ;
        RECT 213.630 23.850 214.060 24.635 ;
        RECT 214.080 23.910 219.590 24.720 ;
        RECT 219.600 23.910 225.110 24.720 ;
        RECT 225.120 23.910 230.630 24.720 ;
        RECT 230.640 23.910 236.150 24.720 ;
        RECT 236.160 23.910 238.910 24.720 ;
        RECT 239.390 23.850 239.820 24.635 ;
        RECT 239.840 23.910 245.350 24.720 ;
        RECT 245.360 23.910 250.870 24.720 ;
        RECT 250.880 23.910 256.390 24.720 ;
        RECT 256.400 23.910 261.910 24.720 ;
        RECT 261.920 23.910 264.670 24.720 ;
        RECT 265.150 23.850 265.580 24.635 ;
        RECT 265.600 23.910 271.110 24.720 ;
        RECT 271.120 23.910 276.630 24.720 ;
        RECT 276.640 23.910 282.150 24.720 ;
        RECT 282.160 23.910 287.670 24.720 ;
        RECT 287.680 23.910 290.430 24.720 ;
        RECT 290.910 23.850 291.340 24.635 ;
        RECT 291.360 23.910 296.870 24.720 ;
        RECT 296.880 23.910 302.390 24.720 ;
        RECT 302.400 23.910 307.910 24.720 ;
        RECT 307.920 23.910 309.750 24.720 ;
        RECT 309.760 23.910 311.130 24.720 ;
      LAYER nwell ;
        RECT 161.905 20.690 311.325 23.520 ;
      LAYER pwell ;
        RECT 162.100 19.490 163.470 20.300 ;
        RECT 163.480 19.490 168.990 20.300 ;
        RECT 169.000 19.490 174.510 20.300 ;
        RECT 174.990 19.575 175.420 20.360 ;
        RECT 175.440 19.490 180.950 20.300 ;
        RECT 180.960 19.490 186.470 20.300 ;
        RECT 186.480 19.490 191.990 20.300 ;
        RECT 192.000 19.490 197.510 20.300 ;
        RECT 197.520 19.490 200.270 20.300 ;
        RECT 200.750 19.575 201.180 20.360 ;
        RECT 201.200 19.490 206.710 20.300 ;
        RECT 206.720 19.490 212.230 20.300 ;
        RECT 212.240 19.490 217.750 20.300 ;
        RECT 217.760 19.490 223.270 20.300 ;
        RECT 223.280 19.490 226.030 20.300 ;
        RECT 226.510 19.575 226.940 20.360 ;
        RECT 226.960 19.490 232.470 20.300 ;
        RECT 232.480 19.490 237.990 20.300 ;
        RECT 238.000 19.490 243.510 20.300 ;
        RECT 243.520 19.490 249.030 20.300 ;
        RECT 249.040 19.490 251.790 20.300 ;
        RECT 252.270 19.575 252.700 20.360 ;
        RECT 252.720 19.490 258.230 20.300 ;
        RECT 258.240 19.490 263.750 20.300 ;
        RECT 263.760 19.490 269.270 20.300 ;
        RECT 269.280 19.490 274.790 20.300 ;
        RECT 274.800 19.490 277.550 20.300 ;
        RECT 278.030 19.575 278.460 20.360 ;
        RECT 278.480 19.490 283.990 20.300 ;
        RECT 284.000 19.490 289.510 20.300 ;
        RECT 289.520 19.490 295.030 20.300 ;
        RECT 295.040 19.490 300.550 20.300 ;
        RECT 300.560 19.490 303.310 20.300 ;
        RECT 303.790 19.575 304.220 20.360 ;
        RECT 304.240 19.490 309.750 20.300 ;
        RECT 309.760 19.490 311.130 20.300 ;
        RECT 162.240 19.280 162.410 19.490 ;
        RECT 163.620 19.280 163.790 19.490 ;
        RECT 169.140 19.280 169.310 19.490 ;
        RECT 174.660 19.440 174.830 19.470 ;
        RECT 174.655 19.330 174.830 19.440 ;
        RECT 174.660 19.280 174.830 19.330 ;
        RECT 175.580 19.300 175.750 19.490 ;
        RECT 180.180 19.280 180.350 19.470 ;
        RECT 181.100 19.300 181.270 19.490 ;
        RECT 185.700 19.280 185.870 19.470 ;
        RECT 186.620 19.300 186.790 19.490 ;
        RECT 187.535 19.330 187.655 19.440 ;
        RECT 188.460 19.280 188.630 19.470 ;
        RECT 192.140 19.300 192.310 19.490 ;
        RECT 193.980 19.280 194.150 19.470 ;
        RECT 197.660 19.300 197.830 19.490 ;
        RECT 199.500 19.280 199.670 19.470 ;
        RECT 200.415 19.330 200.535 19.440 ;
        RECT 201.340 19.300 201.510 19.490 ;
        RECT 205.020 19.280 205.190 19.470 ;
        RECT 206.860 19.300 207.030 19.490 ;
        RECT 210.540 19.280 210.710 19.470 ;
        RECT 212.380 19.300 212.550 19.490 ;
        RECT 213.295 19.330 213.415 19.440 ;
        RECT 214.220 19.280 214.390 19.470 ;
        RECT 217.900 19.300 218.070 19.490 ;
        RECT 219.740 19.280 219.910 19.470 ;
        RECT 223.420 19.300 223.590 19.490 ;
        RECT 225.260 19.280 225.430 19.470 ;
        RECT 226.175 19.330 226.295 19.440 ;
        RECT 227.100 19.300 227.270 19.490 ;
        RECT 230.780 19.280 230.950 19.470 ;
        RECT 232.620 19.300 232.790 19.490 ;
        RECT 236.300 19.280 236.470 19.470 ;
        RECT 238.140 19.300 238.310 19.490 ;
        RECT 239.055 19.330 239.175 19.440 ;
        RECT 239.980 19.280 240.150 19.470 ;
        RECT 243.660 19.300 243.830 19.490 ;
        RECT 245.500 19.280 245.670 19.470 ;
        RECT 249.180 19.300 249.350 19.490 ;
        RECT 251.020 19.280 251.190 19.470 ;
        RECT 251.935 19.330 252.055 19.440 ;
        RECT 252.860 19.300 253.030 19.490 ;
        RECT 256.540 19.280 256.710 19.470 ;
        RECT 258.380 19.300 258.550 19.490 ;
        RECT 262.060 19.280 262.230 19.470 ;
        RECT 263.900 19.300 264.070 19.490 ;
        RECT 264.815 19.330 264.935 19.440 ;
        RECT 265.740 19.280 265.910 19.470 ;
        RECT 269.420 19.300 269.590 19.490 ;
        RECT 271.260 19.280 271.430 19.470 ;
        RECT 274.940 19.300 275.110 19.490 ;
        RECT 276.780 19.280 276.950 19.470 ;
        RECT 277.695 19.330 277.815 19.440 ;
        RECT 278.620 19.300 278.790 19.490 ;
        RECT 282.300 19.280 282.470 19.470 ;
        RECT 284.140 19.300 284.310 19.490 ;
        RECT 287.820 19.280 287.990 19.470 ;
        RECT 289.660 19.300 289.830 19.490 ;
        RECT 290.575 19.330 290.695 19.440 ;
        RECT 291.500 19.280 291.670 19.470 ;
        RECT 295.180 19.300 295.350 19.490 ;
        RECT 297.020 19.280 297.190 19.470 ;
        RECT 300.700 19.300 300.870 19.490 ;
        RECT 302.540 19.280 302.710 19.470 ;
        RECT 303.455 19.330 303.575 19.440 ;
        RECT 304.380 19.300 304.550 19.490 ;
        RECT 308.060 19.280 308.230 19.470 ;
        RECT 310.820 19.280 310.990 19.490 ;
        RECT 162.100 18.470 163.470 19.280 ;
        RECT 163.480 18.470 168.990 19.280 ;
        RECT 169.000 18.470 174.510 19.280 ;
        RECT 174.520 18.470 180.030 19.280 ;
        RECT 180.040 18.470 185.550 19.280 ;
        RECT 185.560 18.470 187.390 19.280 ;
        RECT 187.870 18.410 188.300 19.195 ;
        RECT 188.320 18.470 193.830 19.280 ;
        RECT 193.840 18.470 199.350 19.280 ;
        RECT 199.360 18.470 204.870 19.280 ;
        RECT 204.880 18.470 210.390 19.280 ;
        RECT 210.400 18.470 213.150 19.280 ;
        RECT 213.630 18.410 214.060 19.195 ;
        RECT 214.080 18.470 219.590 19.280 ;
        RECT 219.600 18.470 225.110 19.280 ;
        RECT 225.120 18.470 230.630 19.280 ;
        RECT 230.640 18.470 236.150 19.280 ;
        RECT 236.160 18.470 238.910 19.280 ;
        RECT 239.390 18.410 239.820 19.195 ;
        RECT 239.840 18.470 245.350 19.280 ;
        RECT 245.360 18.470 250.870 19.280 ;
        RECT 250.880 18.470 256.390 19.280 ;
        RECT 256.400 18.470 261.910 19.280 ;
        RECT 261.920 18.470 264.670 19.280 ;
        RECT 265.150 18.410 265.580 19.195 ;
        RECT 265.600 18.470 271.110 19.280 ;
        RECT 271.120 18.470 276.630 19.280 ;
        RECT 276.640 18.470 282.150 19.280 ;
        RECT 282.160 18.470 287.670 19.280 ;
        RECT 287.680 18.470 290.430 19.280 ;
        RECT 290.910 18.410 291.340 19.195 ;
        RECT 291.360 18.470 296.870 19.280 ;
        RECT 296.880 18.470 302.390 19.280 ;
        RECT 302.400 18.470 307.910 19.280 ;
        RECT 307.920 18.470 309.750 19.280 ;
        RECT 309.760 18.470 311.130 19.280 ;
      LAYER nwell ;
        RECT 161.905 15.250 311.325 18.080 ;
      LAYER pwell ;
        RECT 162.100 14.050 163.470 14.860 ;
        RECT 163.480 14.050 168.990 14.860 ;
        RECT 169.000 14.050 174.510 14.860 ;
        RECT 174.990 14.135 175.420 14.920 ;
        RECT 175.440 14.050 180.950 14.860 ;
        RECT 180.960 14.050 186.470 14.860 ;
        RECT 186.480 14.050 187.850 14.860 ;
        RECT 187.870 14.135 188.300 14.920 ;
        RECT 188.320 14.050 193.830 14.860 ;
        RECT 193.840 14.050 199.350 14.860 ;
        RECT 199.360 14.050 200.730 14.860 ;
        RECT 200.750 14.135 201.180 14.920 ;
        RECT 201.200 14.050 206.710 14.860 ;
        RECT 206.720 14.050 212.230 14.860 ;
        RECT 212.240 14.050 213.610 14.860 ;
        RECT 213.630 14.135 214.060 14.920 ;
        RECT 214.080 14.050 219.590 14.860 ;
        RECT 219.600 14.050 225.110 14.860 ;
        RECT 225.120 14.050 226.490 14.860 ;
        RECT 226.510 14.135 226.940 14.920 ;
        RECT 226.960 14.050 232.470 14.860 ;
        RECT 232.480 14.050 237.990 14.860 ;
        RECT 238.000 14.050 239.370 14.860 ;
        RECT 239.390 14.135 239.820 14.920 ;
        RECT 239.840 14.050 245.350 14.860 ;
        RECT 245.360 14.050 250.870 14.860 ;
        RECT 250.880 14.050 252.250 14.860 ;
        RECT 252.270 14.135 252.700 14.920 ;
        RECT 252.720 14.050 258.230 14.860 ;
        RECT 258.240 14.050 263.750 14.860 ;
        RECT 263.760 14.050 265.130 14.860 ;
        RECT 265.150 14.135 265.580 14.920 ;
        RECT 265.600 14.050 271.110 14.860 ;
        RECT 271.120 14.050 276.630 14.860 ;
        RECT 276.640 14.050 278.010 14.860 ;
        RECT 278.030 14.135 278.460 14.920 ;
        RECT 278.480 14.050 283.990 14.860 ;
        RECT 284.000 14.050 289.510 14.860 ;
        RECT 289.520 14.050 290.890 14.860 ;
        RECT 290.910 14.135 291.340 14.920 ;
        RECT 291.360 14.050 296.870 14.860 ;
        RECT 296.880 14.050 302.390 14.860 ;
        RECT 302.400 14.050 303.770 14.860 ;
        RECT 303.790 14.135 304.220 14.920 ;
        RECT 304.240 14.050 309.750 14.860 ;
        RECT 309.760 14.050 311.130 14.860 ;
        RECT 162.240 13.860 162.410 14.050 ;
        RECT 163.620 13.860 163.790 14.050 ;
        RECT 169.140 13.860 169.310 14.050 ;
        RECT 174.655 13.890 174.775 14.000 ;
        RECT 175.580 13.860 175.750 14.050 ;
        RECT 181.100 13.860 181.270 14.050 ;
        RECT 186.620 13.860 186.790 14.050 ;
        RECT 188.460 13.860 188.630 14.050 ;
        RECT 193.980 13.860 194.150 14.050 ;
        RECT 199.500 13.860 199.670 14.050 ;
        RECT 201.340 13.860 201.510 14.050 ;
        RECT 206.860 13.860 207.030 14.050 ;
        RECT 212.380 13.860 212.550 14.050 ;
        RECT 214.220 13.860 214.390 14.050 ;
        RECT 219.740 13.860 219.910 14.050 ;
        RECT 225.260 13.860 225.430 14.050 ;
        RECT 227.100 13.860 227.270 14.050 ;
        RECT 232.620 13.860 232.790 14.050 ;
        RECT 238.140 13.860 238.310 14.050 ;
        RECT 239.980 13.860 240.150 14.050 ;
        RECT 245.500 13.860 245.670 14.050 ;
        RECT 251.020 13.860 251.190 14.050 ;
        RECT 252.860 13.860 253.030 14.050 ;
        RECT 258.380 13.860 258.550 14.050 ;
        RECT 263.900 13.860 264.070 14.050 ;
        RECT 265.740 13.860 265.910 14.050 ;
        RECT 271.260 13.860 271.430 14.050 ;
        RECT 276.780 13.860 276.950 14.050 ;
        RECT 278.620 13.860 278.790 14.050 ;
        RECT 284.140 13.860 284.310 14.050 ;
        RECT 289.660 13.860 289.830 14.050 ;
        RECT 291.500 13.860 291.670 14.050 ;
        RECT 297.020 13.860 297.190 14.050 ;
        RECT 302.540 13.860 302.710 14.050 ;
        RECT 304.380 13.860 304.550 14.050 ;
        RECT 310.820 13.860 310.990 14.050 ;
      LAYER nwell ;
        RECT 3.250 3.250 156.750 5.750 ;
      LAYER li1 ;
        RECT 4.300 222.030 102.625 222.430 ;
        RECT 4.300 4.700 4.700 222.030 ;
        RECT 62.895 216.545 99.045 217.075 ;
        RECT 62.895 213.695 63.425 216.545 ;
        RECT 63.925 215.855 80.385 216.025 ;
        RECT 63.925 214.385 64.155 215.855 ;
        RECT 80.155 214.385 80.385 215.855 ;
        RECT 63.925 214.215 80.385 214.385 ;
        RECT 80.885 213.695 81.055 216.545 ;
        RECT 81.555 215.855 98.015 216.025 ;
        RECT 81.555 214.385 81.785 215.855 ;
        RECT 97.785 214.385 98.015 215.855 ;
        RECT 81.555 214.215 98.015 214.385 ;
        RECT 98.515 213.695 99.045 216.545 ;
        RECT 62.895 213.525 99.045 213.695 ;
        RECT 9.325 211.690 45.335 211.860 ;
        RECT 9.325 201.840 9.495 211.690 ;
        RECT 10.225 211.000 18.225 211.170 ;
        RECT 18.515 211.000 26.515 211.170 ;
        RECT 9.995 202.745 10.165 210.785 ;
        RECT 18.285 202.745 18.455 210.785 ;
        RECT 26.575 202.745 26.745 210.785 ;
        RECT 10.225 202.360 18.225 202.530 ;
        RECT 18.515 202.360 26.515 202.530 ;
        RECT 27.245 201.840 27.415 211.690 ;
        RECT 28.145 211.000 36.145 211.170 ;
        RECT 36.435 211.000 44.435 211.170 ;
        RECT 27.915 202.745 28.085 210.785 ;
        RECT 36.205 202.745 36.375 210.785 ;
        RECT 44.495 202.745 44.665 210.785 ;
        RECT 28.145 202.360 36.145 202.530 ;
        RECT 36.435 202.360 44.435 202.530 ;
        RECT 45.165 201.840 45.335 211.690 ;
        RECT 62.895 210.675 63.425 213.525 ;
        RECT 64.155 212.835 80.155 213.005 ;
        RECT 63.925 211.580 64.095 212.620 ;
        RECT 80.215 211.580 80.385 212.620 ;
        RECT 64.155 211.195 80.155 211.365 ;
        RECT 80.885 210.675 81.055 213.525 ;
        RECT 81.785 212.835 97.785 213.005 ;
        RECT 81.555 211.580 81.725 212.620 ;
        RECT 97.845 211.580 98.015 212.620 ;
        RECT 81.785 211.195 97.785 211.365 ;
        RECT 98.515 210.675 99.045 213.525 ;
        RECT 62.895 210.505 99.045 210.675 ;
        RECT 9.325 201.670 45.335 201.840 ;
        RECT 9.325 191.820 9.495 201.670 ;
        RECT 10.225 200.980 18.225 201.150 ;
        RECT 18.515 200.980 26.515 201.150 ;
        RECT 9.995 192.725 10.165 200.765 ;
        RECT 18.285 192.725 18.455 200.765 ;
        RECT 26.575 192.725 26.745 200.765 ;
        RECT 10.225 192.340 18.225 192.510 ;
        RECT 18.515 192.340 26.515 192.510 ;
        RECT 27.245 191.820 27.415 201.670 ;
        RECT 28.145 200.980 36.145 201.150 ;
        RECT 36.435 200.980 44.435 201.150 ;
        RECT 27.915 192.725 28.085 200.765 ;
        RECT 36.205 192.725 36.375 200.765 ;
        RECT 44.495 192.725 44.665 200.765 ;
        RECT 28.145 192.340 36.145 192.510 ;
        RECT 36.435 192.340 44.435 192.510 ;
        RECT 45.165 191.820 45.335 201.670 ;
        RECT 9.325 191.650 45.335 191.820 ;
        RECT 49.250 210.180 56.310 210.350 ;
        RECT 9.325 190.700 15.415 190.870 ;
        RECT 9.325 180.850 9.495 190.700 ;
        RECT 10.225 190.010 12.225 190.180 ;
        RECT 12.515 190.010 14.515 190.180 ;
        RECT 9.995 181.755 10.165 189.795 ;
        RECT 12.285 181.755 12.455 189.795 ;
        RECT 14.575 181.755 14.745 189.795 ;
        RECT 10.225 181.370 12.225 181.540 ;
        RECT 12.515 181.370 14.515 181.540 ;
        RECT 15.245 180.850 15.415 190.700 ;
        RECT 9.325 180.680 15.415 180.850 ;
        RECT 16.345 190.700 45.335 190.870 ;
        RECT 16.345 180.850 16.515 190.700 ;
        RECT 17.245 190.010 19.245 190.180 ;
        RECT 19.535 190.010 21.535 190.180 ;
        RECT 21.825 190.010 23.825 190.180 ;
        RECT 24.115 190.010 26.115 190.180 ;
        RECT 26.405 190.010 28.405 190.180 ;
        RECT 28.695 190.010 30.695 190.180 ;
        RECT 30.985 190.010 32.985 190.180 ;
        RECT 33.275 190.010 35.275 190.180 ;
        RECT 35.565 190.010 37.565 190.180 ;
        RECT 37.855 190.010 39.855 190.180 ;
        RECT 40.145 190.010 42.145 190.180 ;
        RECT 42.435 190.010 44.435 190.180 ;
        RECT 17.015 181.755 17.185 189.795 ;
        RECT 19.305 181.755 19.475 189.795 ;
        RECT 21.595 181.755 21.765 189.795 ;
        RECT 23.885 181.755 24.055 189.795 ;
        RECT 26.175 181.755 26.345 189.795 ;
        RECT 28.465 181.755 28.635 189.795 ;
        RECT 30.755 181.755 30.925 189.795 ;
        RECT 33.045 181.755 33.215 189.795 ;
        RECT 35.335 181.755 35.505 189.795 ;
        RECT 37.625 181.755 37.795 189.795 ;
        RECT 39.915 181.755 40.085 189.795 ;
        RECT 42.205 181.755 42.375 189.795 ;
        RECT 44.495 181.755 44.665 189.795 ;
        RECT 17.245 181.370 19.245 181.540 ;
        RECT 19.535 181.370 21.535 181.540 ;
        RECT 21.825 181.370 23.825 181.540 ;
        RECT 24.115 181.370 26.115 181.540 ;
        RECT 26.405 181.370 28.405 181.540 ;
        RECT 28.695 181.370 30.695 181.540 ;
        RECT 30.985 181.370 32.985 181.540 ;
        RECT 33.275 181.370 35.275 181.540 ;
        RECT 35.565 181.370 37.565 181.540 ;
        RECT 37.855 181.370 39.855 181.540 ;
        RECT 40.145 181.370 42.145 181.540 ;
        RECT 42.435 181.370 44.435 181.540 ;
        RECT 45.165 180.850 45.335 190.700 ;
        RECT 49.250 187.850 49.420 210.180 ;
        RECT 50.095 207.435 50.785 209.595 ;
        RECT 51.265 207.435 51.955 209.595 ;
        RECT 52.435 207.435 53.125 209.595 ;
        RECT 53.605 207.435 54.295 209.595 ;
        RECT 54.775 207.435 55.465 209.595 ;
        RECT 50.095 188.435 50.785 190.595 ;
        RECT 51.265 188.435 51.955 190.595 ;
        RECT 52.435 188.435 53.125 190.595 ;
        RECT 53.605 188.435 54.295 190.595 ;
        RECT 54.775 188.435 55.465 190.595 ;
        RECT 56.140 187.850 56.310 210.180 ;
        RECT 49.250 187.680 56.310 187.850 ;
        RECT 62.895 207.655 63.425 210.505 ;
        RECT 64.155 209.815 80.155 209.985 ;
        RECT 63.925 208.560 64.095 209.600 ;
        RECT 80.215 208.560 80.385 209.600 ;
        RECT 64.155 208.175 80.155 208.345 ;
        RECT 80.885 207.655 81.055 210.505 ;
        RECT 81.785 209.815 97.785 209.985 ;
        RECT 81.555 208.560 81.725 209.600 ;
        RECT 97.845 208.560 98.015 209.600 ;
        RECT 81.785 208.175 97.785 208.345 ;
        RECT 98.515 207.655 99.045 210.505 ;
        RECT 62.895 207.485 99.045 207.655 ;
        RECT 62.895 204.635 63.425 207.485 ;
        RECT 64.155 206.795 80.155 206.965 ;
        RECT 63.925 205.540 64.095 206.580 ;
        RECT 80.215 205.540 80.385 206.580 ;
        RECT 64.155 205.155 80.155 205.325 ;
        RECT 80.885 204.635 81.055 207.485 ;
        RECT 81.785 206.795 97.785 206.965 ;
        RECT 81.555 205.540 81.725 206.580 ;
        RECT 97.845 205.540 98.015 206.580 ;
        RECT 81.785 205.155 97.785 205.325 ;
        RECT 98.515 204.635 99.045 207.485 ;
        RECT 62.895 204.465 99.045 204.635 ;
        RECT 62.895 201.615 63.425 204.465 ;
        RECT 64.155 203.775 80.155 203.945 ;
        RECT 63.925 202.520 64.095 203.560 ;
        RECT 80.215 202.520 80.385 203.560 ;
        RECT 64.155 202.135 80.155 202.305 ;
        RECT 80.885 201.615 81.055 204.465 ;
        RECT 81.785 203.775 97.785 203.945 ;
        RECT 81.555 202.520 81.725 203.560 ;
        RECT 97.845 202.520 98.015 203.560 ;
        RECT 81.785 202.135 97.785 202.305 ;
        RECT 98.515 201.615 99.045 204.465 ;
        RECT 62.895 201.445 99.045 201.615 ;
        RECT 62.895 198.595 63.425 201.445 ;
        RECT 64.155 200.755 80.155 200.925 ;
        RECT 63.925 199.500 64.095 200.540 ;
        RECT 80.215 199.500 80.385 200.540 ;
        RECT 64.155 199.115 80.155 199.285 ;
        RECT 80.885 198.595 81.055 201.445 ;
        RECT 81.785 200.755 97.785 200.925 ;
        RECT 81.555 199.500 81.725 200.540 ;
        RECT 97.845 199.500 98.015 200.540 ;
        RECT 81.785 199.115 97.785 199.285 ;
        RECT 98.515 198.595 99.045 201.445 ;
        RECT 62.895 198.425 99.045 198.595 ;
        RECT 62.895 195.575 63.425 198.425 ;
        RECT 64.155 197.735 80.155 197.905 ;
        RECT 63.925 196.480 64.095 197.520 ;
        RECT 80.215 196.480 80.385 197.520 ;
        RECT 64.155 196.095 80.155 196.265 ;
        RECT 80.885 195.575 81.055 198.425 ;
        RECT 81.785 197.735 97.785 197.905 ;
        RECT 81.555 196.480 81.725 197.520 ;
        RECT 97.845 196.480 98.015 197.520 ;
        RECT 81.785 196.095 97.785 196.265 ;
        RECT 98.515 195.575 99.045 198.425 ;
        RECT 62.895 195.405 99.045 195.575 ;
        RECT 62.895 192.555 63.425 195.405 ;
        RECT 64.155 194.715 80.155 194.885 ;
        RECT 63.925 193.460 64.095 194.500 ;
        RECT 80.215 193.460 80.385 194.500 ;
        RECT 64.155 193.075 80.155 193.245 ;
        RECT 80.885 192.555 81.055 195.405 ;
        RECT 81.785 194.715 97.785 194.885 ;
        RECT 81.555 193.460 81.725 194.500 ;
        RECT 97.845 193.460 98.015 194.500 ;
        RECT 81.785 193.075 97.785 193.245 ;
        RECT 98.515 192.555 99.045 195.405 ;
        RECT 62.895 192.385 99.045 192.555 ;
        RECT 62.895 189.535 63.425 192.385 ;
        RECT 64.155 191.695 80.155 191.865 ;
        RECT 63.925 190.440 64.095 191.480 ;
        RECT 80.215 190.440 80.385 191.480 ;
        RECT 64.155 190.055 80.155 190.225 ;
        RECT 80.885 189.535 81.055 192.385 ;
        RECT 81.785 191.695 97.785 191.865 ;
        RECT 81.555 190.440 81.725 191.480 ;
        RECT 97.845 190.440 98.015 191.480 ;
        RECT 81.785 190.055 97.785 190.225 ;
        RECT 98.515 189.535 99.045 192.385 ;
        RECT 62.895 189.365 99.045 189.535 ;
        RECT 16.345 180.680 45.335 180.850 ;
        RECT 62.895 186.515 63.425 189.365 ;
        RECT 64.155 188.675 80.155 188.845 ;
        RECT 63.925 187.420 64.095 188.460 ;
        RECT 80.215 187.420 80.385 188.460 ;
        RECT 64.155 187.035 80.155 187.205 ;
        RECT 80.885 186.515 81.055 189.365 ;
        RECT 81.785 188.675 97.785 188.845 ;
        RECT 81.555 187.420 81.725 188.460 ;
        RECT 97.845 187.420 98.015 188.460 ;
        RECT 81.785 187.035 97.785 187.205 ;
        RECT 98.515 186.515 99.045 189.365 ;
        RECT 62.895 186.345 99.045 186.515 ;
        RECT 62.895 183.495 63.425 186.345 ;
        RECT 64.155 185.655 80.155 185.825 ;
        RECT 63.925 184.400 64.095 185.440 ;
        RECT 80.215 184.400 80.385 185.440 ;
        RECT 64.155 184.015 80.155 184.185 ;
        RECT 80.885 183.495 81.055 186.345 ;
        RECT 81.785 185.655 97.785 185.825 ;
        RECT 81.555 184.400 81.725 185.440 ;
        RECT 97.845 184.400 98.015 185.440 ;
        RECT 81.785 184.015 97.785 184.185 ;
        RECT 98.515 183.495 99.045 186.345 ;
        RECT 62.895 183.325 99.045 183.495 ;
        RECT 62.895 180.475 63.425 183.325 ;
        RECT 64.155 182.635 80.155 182.805 ;
        RECT 63.925 181.380 64.095 182.420 ;
        RECT 80.215 181.380 80.385 182.420 ;
        RECT 64.155 180.995 80.155 181.165 ;
        RECT 80.885 180.475 81.055 183.325 ;
        RECT 81.785 182.635 97.785 182.805 ;
        RECT 81.555 181.380 81.725 182.420 ;
        RECT 97.845 181.380 98.015 182.420 ;
        RECT 81.785 180.995 97.785 181.165 ;
        RECT 98.515 180.475 99.045 183.325 ;
        RECT 102.225 181.020 102.625 222.030 ;
        RECT 108.630 220.425 153.130 220.595 ;
        RECT 108.630 216.575 108.800 220.425 ;
        RECT 109.585 219.735 110.585 219.905 ;
        RECT 110.875 219.735 111.875 219.905 ;
        RECT 109.355 217.480 109.525 219.520 ;
        RECT 110.645 217.480 110.815 219.520 ;
        RECT 111.935 217.480 112.105 219.520 ;
        RECT 109.585 217.095 110.585 217.265 ;
        RECT 110.875 217.095 111.875 217.265 ;
        RECT 112.660 216.575 112.830 220.425 ;
        RECT 113.615 219.735 114.615 219.905 ;
        RECT 114.905 219.735 115.905 219.905 ;
        RECT 113.385 217.480 113.555 219.520 ;
        RECT 114.675 217.480 114.845 219.520 ;
        RECT 115.965 217.480 116.135 219.520 ;
        RECT 113.615 217.095 114.615 217.265 ;
        RECT 114.905 217.095 115.905 217.265 ;
        RECT 116.690 216.575 116.860 220.425 ;
        RECT 117.645 219.735 118.645 219.905 ;
        RECT 118.935 219.735 119.935 219.905 ;
        RECT 117.415 217.480 117.585 219.520 ;
        RECT 118.705 217.480 118.875 219.520 ;
        RECT 119.995 217.480 120.165 219.520 ;
        RECT 117.645 217.095 118.645 217.265 ;
        RECT 118.935 217.095 119.935 217.265 ;
        RECT 120.720 216.575 120.890 220.425 ;
        RECT 121.675 219.735 122.675 219.905 ;
        RECT 122.965 219.735 123.965 219.905 ;
        RECT 121.445 217.480 121.615 219.520 ;
        RECT 122.735 217.480 122.905 219.520 ;
        RECT 124.025 217.480 124.195 219.520 ;
        RECT 121.675 217.095 122.675 217.265 ;
        RECT 122.965 217.095 123.965 217.265 ;
        RECT 124.750 216.575 124.920 220.425 ;
        RECT 125.705 219.735 126.705 219.905 ;
        RECT 126.995 219.735 127.995 219.905 ;
        RECT 125.475 217.480 125.645 219.520 ;
        RECT 126.765 217.480 126.935 219.520 ;
        RECT 128.055 217.480 128.225 219.520 ;
        RECT 125.705 217.095 126.705 217.265 ;
        RECT 126.995 217.095 127.995 217.265 ;
        RECT 128.780 216.575 128.950 220.425 ;
        RECT 129.735 219.735 130.735 219.905 ;
        RECT 131.025 219.735 132.025 219.905 ;
        RECT 129.505 217.480 129.675 219.520 ;
        RECT 130.795 217.480 130.965 219.520 ;
        RECT 132.085 217.480 132.255 219.520 ;
        RECT 129.735 217.095 130.735 217.265 ;
        RECT 131.025 217.095 132.025 217.265 ;
        RECT 132.810 216.575 132.980 220.425 ;
        RECT 133.765 219.735 134.765 219.905 ;
        RECT 135.055 219.735 136.055 219.905 ;
        RECT 133.535 217.480 133.705 219.520 ;
        RECT 134.825 217.480 134.995 219.520 ;
        RECT 136.115 217.480 136.285 219.520 ;
        RECT 133.765 217.095 134.765 217.265 ;
        RECT 135.055 217.095 136.055 217.265 ;
        RECT 136.840 216.575 137.010 220.425 ;
        RECT 137.795 219.735 138.795 219.905 ;
        RECT 139.085 219.735 140.085 219.905 ;
        RECT 137.565 217.480 137.735 219.520 ;
        RECT 138.855 217.480 139.025 219.520 ;
        RECT 140.145 217.480 140.315 219.520 ;
        RECT 137.795 217.095 138.795 217.265 ;
        RECT 139.085 217.095 140.085 217.265 ;
        RECT 140.870 216.575 141.040 220.425 ;
        RECT 141.825 219.735 142.825 219.905 ;
        RECT 143.115 219.735 144.115 219.905 ;
        RECT 141.595 217.480 141.765 219.520 ;
        RECT 142.885 217.480 143.055 219.520 ;
        RECT 144.175 217.480 144.345 219.520 ;
        RECT 141.825 217.095 142.825 217.265 ;
        RECT 143.115 217.095 144.115 217.265 ;
        RECT 144.900 216.575 145.070 220.425 ;
        RECT 145.855 219.735 146.855 219.905 ;
        RECT 147.145 219.735 148.145 219.905 ;
        RECT 145.625 217.480 145.795 219.520 ;
        RECT 146.915 217.480 147.085 219.520 ;
        RECT 148.205 217.480 148.375 219.520 ;
        RECT 145.855 217.095 146.855 217.265 ;
        RECT 147.145 217.095 148.145 217.265 ;
        RECT 148.930 216.575 149.100 220.425 ;
        RECT 149.885 219.735 150.885 219.905 ;
        RECT 151.175 219.735 152.175 219.905 ;
        RECT 149.655 217.480 149.825 219.520 ;
        RECT 150.945 217.480 151.115 219.520 ;
        RECT 152.235 217.480 152.405 219.520 ;
        RECT 149.885 217.095 150.885 217.265 ;
        RECT 151.175 217.095 152.175 217.265 ;
        RECT 152.960 216.575 153.130 220.425 ;
        RECT 108.630 216.405 153.130 216.575 ;
        RECT 108.630 213.455 153.130 213.625 ;
        RECT 108.630 203.605 108.800 213.455 ;
        RECT 109.585 212.765 110.585 212.935 ;
        RECT 110.875 212.765 111.875 212.935 ;
        RECT 109.355 204.510 109.525 212.550 ;
        RECT 110.645 204.510 110.815 212.550 ;
        RECT 111.935 204.510 112.105 212.550 ;
        RECT 109.585 204.125 110.585 204.295 ;
        RECT 110.875 204.125 111.875 204.295 ;
        RECT 112.660 203.605 112.830 213.455 ;
        RECT 113.615 212.765 114.615 212.935 ;
        RECT 114.905 212.765 115.905 212.935 ;
        RECT 113.385 204.510 113.555 212.550 ;
        RECT 114.675 204.510 114.845 212.550 ;
        RECT 115.965 204.510 116.135 212.550 ;
        RECT 113.615 204.125 114.615 204.295 ;
        RECT 114.905 204.125 115.905 204.295 ;
        RECT 116.690 203.605 116.860 213.455 ;
        RECT 117.645 212.765 118.645 212.935 ;
        RECT 118.935 212.765 119.935 212.935 ;
        RECT 117.415 204.510 117.585 212.550 ;
        RECT 118.705 204.510 118.875 212.550 ;
        RECT 119.995 204.510 120.165 212.550 ;
        RECT 117.645 204.125 118.645 204.295 ;
        RECT 118.935 204.125 119.935 204.295 ;
        RECT 120.720 203.605 120.890 213.455 ;
        RECT 121.675 212.765 122.675 212.935 ;
        RECT 122.965 212.765 123.965 212.935 ;
        RECT 121.445 204.510 121.615 212.550 ;
        RECT 122.735 204.510 122.905 212.550 ;
        RECT 124.025 204.510 124.195 212.550 ;
        RECT 121.675 204.125 122.675 204.295 ;
        RECT 122.965 204.125 123.965 204.295 ;
        RECT 124.750 203.605 124.920 213.455 ;
        RECT 125.705 212.765 126.705 212.935 ;
        RECT 126.995 212.765 127.995 212.935 ;
        RECT 125.475 204.510 125.645 212.550 ;
        RECT 126.765 204.510 126.935 212.550 ;
        RECT 128.055 204.510 128.225 212.550 ;
        RECT 125.705 204.125 126.705 204.295 ;
        RECT 126.995 204.125 127.995 204.295 ;
        RECT 128.780 203.605 128.950 213.455 ;
        RECT 129.735 212.765 130.735 212.935 ;
        RECT 131.025 212.765 132.025 212.935 ;
        RECT 129.505 204.510 129.675 212.550 ;
        RECT 130.795 204.510 130.965 212.550 ;
        RECT 132.085 204.510 132.255 212.550 ;
        RECT 129.735 204.125 130.735 204.295 ;
        RECT 131.025 204.125 132.025 204.295 ;
        RECT 132.810 203.605 132.980 213.455 ;
        RECT 133.765 212.765 134.765 212.935 ;
        RECT 135.055 212.765 136.055 212.935 ;
        RECT 133.535 204.510 133.705 212.550 ;
        RECT 134.825 204.510 134.995 212.550 ;
        RECT 136.115 204.510 136.285 212.550 ;
        RECT 133.765 204.125 134.765 204.295 ;
        RECT 135.055 204.125 136.055 204.295 ;
        RECT 136.840 203.605 137.010 213.455 ;
        RECT 137.795 212.765 138.795 212.935 ;
        RECT 139.085 212.765 140.085 212.935 ;
        RECT 137.565 204.510 137.735 212.550 ;
        RECT 138.855 204.510 139.025 212.550 ;
        RECT 140.145 204.510 140.315 212.550 ;
        RECT 137.795 204.125 138.795 204.295 ;
        RECT 139.085 204.125 140.085 204.295 ;
        RECT 140.870 203.605 141.040 213.455 ;
        RECT 141.825 212.765 142.825 212.935 ;
        RECT 143.115 212.765 144.115 212.935 ;
        RECT 141.595 204.510 141.765 212.550 ;
        RECT 142.885 204.510 143.055 212.550 ;
        RECT 144.175 204.510 144.345 212.550 ;
        RECT 141.825 204.125 142.825 204.295 ;
        RECT 143.115 204.125 144.115 204.295 ;
        RECT 144.900 203.605 145.070 213.455 ;
        RECT 145.855 212.765 146.855 212.935 ;
        RECT 147.145 212.765 148.145 212.935 ;
        RECT 145.625 204.510 145.795 212.550 ;
        RECT 146.915 204.510 147.085 212.550 ;
        RECT 148.205 204.510 148.375 212.550 ;
        RECT 145.855 204.125 146.855 204.295 ;
        RECT 147.145 204.125 148.145 204.295 ;
        RECT 148.930 203.605 149.100 213.455 ;
        RECT 149.885 212.765 150.885 212.935 ;
        RECT 151.175 212.765 152.175 212.935 ;
        RECT 149.655 204.510 149.825 212.550 ;
        RECT 150.945 204.510 151.115 212.550 ;
        RECT 152.235 204.510 152.405 212.550 ;
        RECT 149.885 204.125 150.885 204.295 ;
        RECT 151.175 204.125 152.175 204.295 ;
        RECT 152.960 203.605 153.130 213.455 ;
        RECT 108.630 203.435 153.130 203.605 ;
        RECT 162.095 201.405 236.155 201.575 ;
        RECT 108.630 200.740 153.130 200.910 ;
        RECT 108.630 194.980 108.800 200.740 ;
        RECT 109.585 200.050 110.585 200.220 ;
        RECT 110.875 200.050 111.875 200.220 ;
        RECT 109.355 195.840 109.525 199.880 ;
        RECT 110.645 195.840 110.815 199.880 ;
        RECT 111.935 195.840 112.105 199.880 ;
        RECT 109.585 195.500 110.585 195.670 ;
        RECT 110.875 195.500 111.875 195.670 ;
        RECT 112.660 194.980 112.830 200.740 ;
        RECT 113.615 200.050 114.615 200.220 ;
        RECT 114.905 200.050 115.905 200.220 ;
        RECT 113.385 195.840 113.555 199.880 ;
        RECT 114.675 195.840 114.845 199.880 ;
        RECT 115.965 195.840 116.135 199.880 ;
        RECT 113.615 195.500 114.615 195.670 ;
        RECT 114.905 195.500 115.905 195.670 ;
        RECT 116.690 194.980 116.860 200.740 ;
        RECT 117.645 200.050 118.645 200.220 ;
        RECT 118.935 200.050 119.935 200.220 ;
        RECT 117.415 195.840 117.585 199.880 ;
        RECT 118.705 195.840 118.875 199.880 ;
        RECT 119.995 195.840 120.165 199.880 ;
        RECT 117.645 195.500 118.645 195.670 ;
        RECT 118.935 195.500 119.935 195.670 ;
        RECT 120.720 194.980 120.890 200.740 ;
        RECT 121.675 200.050 122.675 200.220 ;
        RECT 122.965 200.050 123.965 200.220 ;
        RECT 121.445 195.840 121.615 199.880 ;
        RECT 122.735 195.840 122.905 199.880 ;
        RECT 124.025 195.840 124.195 199.880 ;
        RECT 121.675 195.500 122.675 195.670 ;
        RECT 122.965 195.500 123.965 195.670 ;
        RECT 124.750 194.980 124.920 200.740 ;
        RECT 125.705 200.050 126.705 200.220 ;
        RECT 126.995 200.050 127.995 200.220 ;
        RECT 125.475 195.840 125.645 199.880 ;
        RECT 126.765 195.840 126.935 199.880 ;
        RECT 128.055 195.840 128.225 199.880 ;
        RECT 125.705 195.500 126.705 195.670 ;
        RECT 126.995 195.500 127.995 195.670 ;
        RECT 128.780 194.980 128.950 200.740 ;
        RECT 129.735 200.050 130.735 200.220 ;
        RECT 131.025 200.050 132.025 200.220 ;
        RECT 129.505 195.840 129.675 199.880 ;
        RECT 130.795 195.840 130.965 199.880 ;
        RECT 132.085 195.840 132.255 199.880 ;
        RECT 129.735 195.500 130.735 195.670 ;
        RECT 131.025 195.500 132.025 195.670 ;
        RECT 132.810 194.980 132.980 200.740 ;
        RECT 133.765 200.050 134.765 200.220 ;
        RECT 135.055 200.050 136.055 200.220 ;
        RECT 133.535 195.840 133.705 199.880 ;
        RECT 134.825 195.840 134.995 199.880 ;
        RECT 136.115 195.840 136.285 199.880 ;
        RECT 133.765 195.500 134.765 195.670 ;
        RECT 135.055 195.500 136.055 195.670 ;
        RECT 136.840 194.980 137.010 200.740 ;
        RECT 137.795 200.050 138.795 200.220 ;
        RECT 139.085 200.050 140.085 200.220 ;
        RECT 137.565 195.840 137.735 199.880 ;
        RECT 138.855 195.840 139.025 199.880 ;
        RECT 140.145 195.840 140.315 199.880 ;
        RECT 137.795 195.500 138.795 195.670 ;
        RECT 139.085 195.500 140.085 195.670 ;
        RECT 140.870 194.980 141.040 200.740 ;
        RECT 141.825 200.050 142.825 200.220 ;
        RECT 143.115 200.050 144.115 200.220 ;
        RECT 141.595 195.840 141.765 199.880 ;
        RECT 142.885 195.840 143.055 199.880 ;
        RECT 144.175 195.840 144.345 199.880 ;
        RECT 141.825 195.500 142.825 195.670 ;
        RECT 143.115 195.500 144.115 195.670 ;
        RECT 144.900 194.980 145.070 200.740 ;
        RECT 145.855 200.050 146.855 200.220 ;
        RECT 147.145 200.050 148.145 200.220 ;
        RECT 145.625 195.840 145.795 199.880 ;
        RECT 146.915 195.840 147.085 199.880 ;
        RECT 148.205 195.840 148.375 199.880 ;
        RECT 145.855 195.500 146.855 195.670 ;
        RECT 147.145 195.500 148.145 195.670 ;
        RECT 148.930 194.980 149.100 200.740 ;
        RECT 149.885 200.050 150.885 200.220 ;
        RECT 151.175 200.050 152.175 200.220 ;
        RECT 149.655 195.840 149.825 199.880 ;
        RECT 150.945 195.840 151.115 199.880 ;
        RECT 152.235 195.840 152.405 199.880 ;
        RECT 149.885 195.500 150.885 195.670 ;
        RECT 151.175 195.500 152.175 195.670 ;
        RECT 152.960 194.980 153.130 200.740 ;
        RECT 162.180 200.315 163.390 201.405 ;
        RECT 162.180 199.605 162.700 200.145 ;
        RECT 162.870 199.775 163.390 200.315 ;
        RECT 163.560 200.435 163.830 201.205 ;
        RECT 164.000 200.625 164.330 201.405 ;
        RECT 164.535 200.800 164.720 201.205 ;
        RECT 164.890 200.980 165.225 201.405 ;
        RECT 164.535 200.625 165.200 200.800 ;
        RECT 163.560 200.265 164.690 200.435 ;
        RECT 162.180 198.855 163.390 199.605 ;
        RECT 163.560 199.355 163.730 200.265 ;
        RECT 163.900 199.515 164.260 200.095 ;
        RECT 164.440 199.765 164.690 200.265 ;
        RECT 164.860 199.595 165.200 200.625 ;
        RECT 165.865 200.255 166.125 201.405 ;
        RECT 166.300 200.330 166.555 201.235 ;
        RECT 166.725 200.645 167.055 201.405 ;
        RECT 167.270 200.475 167.440 201.235 ;
        RECT 167.700 200.970 173.045 201.405 ;
        RECT 164.515 199.425 165.200 199.595 ;
        RECT 163.560 199.025 163.820 199.355 ;
        RECT 164.030 198.855 164.305 199.335 ;
        RECT 164.515 199.025 164.720 199.425 ;
        RECT 164.890 198.855 165.225 199.255 ;
        RECT 165.865 198.855 166.125 199.695 ;
        RECT 166.300 199.600 166.470 200.330 ;
        RECT 166.725 200.305 167.440 200.475 ;
        RECT 166.725 200.095 166.895 200.305 ;
        RECT 166.640 199.765 166.895 200.095 ;
        RECT 166.300 199.025 166.555 199.600 ;
        RECT 166.725 199.575 166.895 199.765 ;
        RECT 167.175 199.755 167.530 200.125 ;
        RECT 166.725 199.405 167.440 199.575 ;
        RECT 166.725 198.855 167.055 199.235 ;
        RECT 167.270 199.025 167.440 199.405 ;
        RECT 169.285 199.400 169.625 200.230 ;
        RECT 171.105 199.720 171.455 200.970 ;
        RECT 173.220 200.315 174.890 201.405 ;
        RECT 173.220 199.625 173.970 200.145 ;
        RECT 174.140 199.795 174.890 200.315 ;
        RECT 175.060 200.240 175.350 201.405 ;
        RECT 175.610 200.475 175.780 201.235 ;
        RECT 175.995 200.645 176.325 201.405 ;
        RECT 175.610 200.305 176.325 200.475 ;
        RECT 176.495 200.330 176.750 201.235 ;
        RECT 175.520 199.755 175.875 200.125 ;
        RECT 176.155 200.095 176.325 200.305 ;
        RECT 176.155 199.765 176.410 200.095 ;
        RECT 167.700 198.855 173.045 199.400 ;
        RECT 173.220 198.855 174.890 199.625 ;
        RECT 175.060 198.855 175.350 199.580 ;
        RECT 176.155 199.575 176.325 199.765 ;
        RECT 176.580 199.600 176.750 200.330 ;
        RECT 176.925 200.255 177.185 201.405 ;
        RECT 177.360 200.970 182.705 201.405 ;
        RECT 175.610 199.405 176.325 199.575 ;
        RECT 175.610 199.025 175.780 199.405 ;
        RECT 175.995 198.855 176.325 199.235 ;
        RECT 176.495 199.025 176.750 199.600 ;
        RECT 176.925 198.855 177.185 199.695 ;
        RECT 178.945 199.400 179.285 200.230 ;
        RECT 180.765 199.720 181.115 200.970 ;
        RECT 182.880 200.315 184.550 201.405 ;
        RECT 182.880 199.625 183.630 200.145 ;
        RECT 183.800 199.795 184.550 200.315 ;
        RECT 185.270 200.475 185.440 201.235 ;
        RECT 185.655 200.645 185.985 201.405 ;
        RECT 185.270 200.305 185.985 200.475 ;
        RECT 186.155 200.330 186.410 201.235 ;
        RECT 185.180 199.755 185.535 200.125 ;
        RECT 185.815 200.095 185.985 200.305 ;
        RECT 185.815 199.765 186.070 200.095 ;
        RECT 177.360 198.855 182.705 199.400 ;
        RECT 182.880 198.855 184.550 199.625 ;
        RECT 185.815 199.575 185.985 199.765 ;
        RECT 186.240 199.600 186.410 200.330 ;
        RECT 186.585 200.255 186.845 201.405 ;
        RECT 187.940 200.240 188.230 201.405 ;
        RECT 188.400 200.970 193.745 201.405 ;
        RECT 185.270 199.405 185.985 199.575 ;
        RECT 185.270 199.025 185.440 199.405 ;
        RECT 185.655 198.855 185.985 199.235 ;
        RECT 186.155 199.025 186.410 199.600 ;
        RECT 186.585 198.855 186.845 199.695 ;
        RECT 187.940 198.855 188.230 199.580 ;
        RECT 189.985 199.400 190.325 200.230 ;
        RECT 191.805 199.720 192.155 200.970 ;
        RECT 194.930 200.475 195.100 201.235 ;
        RECT 195.315 200.645 195.645 201.405 ;
        RECT 194.930 200.305 195.645 200.475 ;
        RECT 195.815 200.330 196.070 201.235 ;
        RECT 194.840 199.755 195.195 200.125 ;
        RECT 195.475 200.095 195.645 200.305 ;
        RECT 195.475 199.765 195.730 200.095 ;
        RECT 195.475 199.575 195.645 199.765 ;
        RECT 195.900 199.600 196.070 200.330 ;
        RECT 196.245 200.255 196.505 201.405 ;
        RECT 196.680 200.315 200.190 201.405 ;
        RECT 194.930 199.405 195.645 199.575 ;
        RECT 188.400 198.855 193.745 199.400 ;
        RECT 194.930 199.025 195.100 199.405 ;
        RECT 195.315 198.855 195.645 199.235 ;
        RECT 195.815 199.025 196.070 199.600 ;
        RECT 196.245 198.855 196.505 199.695 ;
        RECT 196.680 199.625 198.330 200.145 ;
        RECT 198.500 199.795 200.190 200.315 ;
        RECT 200.820 200.240 201.110 201.405 ;
        RECT 201.280 200.315 203.870 201.405 ;
        RECT 201.280 199.625 202.490 200.145 ;
        RECT 202.660 199.795 203.870 200.315 ;
        RECT 204.590 200.475 204.760 201.235 ;
        RECT 204.975 200.645 205.305 201.405 ;
        RECT 204.590 200.305 205.305 200.475 ;
        RECT 205.475 200.330 205.730 201.235 ;
        RECT 204.500 199.755 204.855 200.125 ;
        RECT 205.135 200.095 205.305 200.305 ;
        RECT 205.135 199.765 205.390 200.095 ;
        RECT 196.680 198.855 200.190 199.625 ;
        RECT 200.820 198.855 201.110 199.580 ;
        RECT 201.280 198.855 203.870 199.625 ;
        RECT 205.135 199.575 205.305 199.765 ;
        RECT 205.560 199.600 205.730 200.330 ;
        RECT 205.905 200.255 206.165 201.405 ;
        RECT 206.340 200.970 211.685 201.405 ;
        RECT 204.590 199.405 205.305 199.575 ;
        RECT 204.590 199.025 204.760 199.405 ;
        RECT 204.975 198.855 205.305 199.235 ;
        RECT 205.475 199.025 205.730 199.600 ;
        RECT 205.905 198.855 206.165 199.695 ;
        RECT 207.925 199.400 208.265 200.230 ;
        RECT 209.745 199.720 210.095 200.970 ;
        RECT 211.860 200.315 213.530 201.405 ;
        RECT 211.860 199.625 212.610 200.145 ;
        RECT 212.780 199.795 213.530 200.315 ;
        RECT 213.700 200.240 213.990 201.405 ;
        RECT 214.250 200.475 214.420 201.235 ;
        RECT 214.635 200.645 214.965 201.405 ;
        RECT 214.250 200.305 214.965 200.475 ;
        RECT 215.135 200.330 215.390 201.235 ;
        RECT 214.160 199.755 214.515 200.125 ;
        RECT 214.795 200.095 214.965 200.305 ;
        RECT 214.795 199.765 215.050 200.095 ;
        RECT 206.340 198.855 211.685 199.400 ;
        RECT 211.860 198.855 213.530 199.625 ;
        RECT 213.700 198.855 213.990 199.580 ;
        RECT 214.795 199.575 214.965 199.765 ;
        RECT 215.220 199.600 215.390 200.330 ;
        RECT 215.565 200.255 215.825 201.405 ;
        RECT 216.000 200.970 221.345 201.405 ;
        RECT 214.250 199.405 214.965 199.575 ;
        RECT 214.250 199.025 214.420 199.405 ;
        RECT 214.635 198.855 214.965 199.235 ;
        RECT 215.135 199.025 215.390 199.600 ;
        RECT 215.565 198.855 215.825 199.695 ;
        RECT 217.585 199.400 217.925 200.230 ;
        RECT 219.405 199.720 219.755 200.970 ;
        RECT 221.520 200.315 223.190 201.405 ;
        RECT 221.520 199.625 222.270 200.145 ;
        RECT 222.440 199.795 223.190 200.315 ;
        RECT 223.910 200.475 224.080 201.235 ;
        RECT 224.295 200.645 224.625 201.405 ;
        RECT 223.910 200.305 224.625 200.475 ;
        RECT 224.795 200.330 225.050 201.235 ;
        RECT 223.820 199.755 224.175 200.125 ;
        RECT 224.455 200.095 224.625 200.305 ;
        RECT 224.455 199.765 224.710 200.095 ;
        RECT 216.000 198.855 221.345 199.400 ;
        RECT 221.520 198.855 223.190 199.625 ;
        RECT 224.455 199.575 224.625 199.765 ;
        RECT 224.880 199.600 225.050 200.330 ;
        RECT 225.225 200.255 225.485 201.405 ;
        RECT 226.580 200.240 226.870 201.405 ;
        RECT 227.040 200.970 232.385 201.405 ;
        RECT 223.910 199.405 224.625 199.575 ;
        RECT 223.910 199.025 224.080 199.405 ;
        RECT 224.295 198.855 224.625 199.235 ;
        RECT 224.795 199.025 225.050 199.600 ;
        RECT 225.225 198.855 225.485 199.695 ;
        RECT 226.580 198.855 226.870 199.580 ;
        RECT 228.625 199.400 228.965 200.230 ;
        RECT 230.445 199.720 230.795 200.970 ;
        RECT 233.110 200.475 233.280 201.235 ;
        RECT 233.495 200.645 233.825 201.405 ;
        RECT 233.110 200.305 233.825 200.475 ;
        RECT 233.995 200.330 234.250 201.235 ;
        RECT 233.020 199.755 233.375 200.125 ;
        RECT 233.655 200.095 233.825 200.305 ;
        RECT 233.655 199.765 233.910 200.095 ;
        RECT 233.655 199.575 233.825 199.765 ;
        RECT 234.080 199.600 234.250 200.330 ;
        RECT 234.425 200.255 234.685 201.405 ;
        RECT 234.860 200.315 236.070 201.405 ;
        RECT 234.860 199.775 235.380 200.315 ;
        RECT 233.110 199.405 233.825 199.575 ;
        RECT 227.040 198.855 232.385 199.400 ;
        RECT 233.110 199.025 233.280 199.405 ;
        RECT 233.495 198.855 233.825 199.235 ;
        RECT 233.995 199.025 234.250 199.600 ;
        RECT 234.425 198.855 234.685 199.695 ;
        RECT 235.550 199.605 236.070 200.145 ;
        RECT 234.860 198.855 236.070 199.605 ;
        RECT 162.095 198.685 236.155 198.855 ;
        RECT 162.180 197.935 163.390 198.685 ;
        RECT 163.560 198.140 168.905 198.685 ;
        RECT 169.080 198.140 174.425 198.685 ;
        RECT 174.600 198.140 179.945 198.685 ;
        RECT 180.120 198.140 185.465 198.685 ;
        RECT 162.180 197.395 162.700 197.935 ;
        RECT 162.870 197.225 163.390 197.765 ;
        RECT 165.145 197.310 165.485 198.140 ;
        RECT 162.180 196.135 163.390 197.225 ;
        RECT 166.965 196.570 167.315 197.820 ;
        RECT 170.665 197.310 171.005 198.140 ;
        RECT 172.485 196.570 172.835 197.820 ;
        RECT 176.185 197.310 176.525 198.140 ;
        RECT 178.005 196.570 178.355 197.820 ;
        RECT 181.705 197.310 182.045 198.140 ;
        RECT 185.640 197.915 187.310 198.685 ;
        RECT 187.940 197.960 188.230 198.685 ;
        RECT 188.400 198.140 193.745 198.685 ;
        RECT 193.920 198.140 199.265 198.685 ;
        RECT 199.440 198.140 204.785 198.685 ;
        RECT 204.960 198.140 210.305 198.685 ;
        RECT 183.525 196.570 183.875 197.820 ;
        RECT 185.640 197.395 186.390 197.915 ;
        RECT 186.560 197.225 187.310 197.745 ;
        RECT 189.985 197.310 190.325 198.140 ;
        RECT 163.560 196.135 168.905 196.570 ;
        RECT 169.080 196.135 174.425 196.570 ;
        RECT 174.600 196.135 179.945 196.570 ;
        RECT 180.120 196.135 185.465 196.570 ;
        RECT 185.640 196.135 187.310 197.225 ;
        RECT 187.940 196.135 188.230 197.300 ;
        RECT 191.805 196.570 192.155 197.820 ;
        RECT 195.505 197.310 195.845 198.140 ;
        RECT 197.325 196.570 197.675 197.820 ;
        RECT 201.025 197.310 201.365 198.140 ;
        RECT 202.845 196.570 203.195 197.820 ;
        RECT 206.545 197.310 206.885 198.140 ;
        RECT 210.480 197.915 213.070 198.685 ;
        RECT 213.700 197.960 213.990 198.685 ;
        RECT 214.160 198.140 219.505 198.685 ;
        RECT 219.680 198.140 225.025 198.685 ;
        RECT 225.200 198.140 230.545 198.685 ;
        RECT 208.365 196.570 208.715 197.820 ;
        RECT 210.480 197.395 211.690 197.915 ;
        RECT 211.860 197.225 213.070 197.745 ;
        RECT 215.745 197.310 216.085 198.140 ;
        RECT 188.400 196.135 193.745 196.570 ;
        RECT 193.920 196.135 199.265 196.570 ;
        RECT 199.440 196.135 204.785 196.570 ;
        RECT 204.960 196.135 210.305 196.570 ;
        RECT 210.480 196.135 213.070 197.225 ;
        RECT 213.700 196.135 213.990 197.300 ;
        RECT 217.565 196.570 217.915 197.820 ;
        RECT 221.265 197.310 221.605 198.140 ;
        RECT 223.085 196.570 223.435 197.820 ;
        RECT 226.785 197.310 227.125 198.140 ;
        RECT 230.720 197.915 234.230 198.685 ;
        RECT 234.860 197.935 236.070 198.685 ;
        RECT 228.605 196.570 228.955 197.820 ;
        RECT 230.720 197.395 232.370 197.915 ;
        RECT 232.540 197.225 234.230 197.745 ;
        RECT 214.160 196.135 219.505 196.570 ;
        RECT 219.680 196.135 225.025 196.570 ;
        RECT 225.200 196.135 230.545 196.570 ;
        RECT 230.720 196.135 234.230 197.225 ;
        RECT 234.860 197.225 235.380 197.765 ;
        RECT 235.550 197.395 236.070 197.935 ;
        RECT 234.860 196.135 236.070 197.225 ;
        RECT 162.095 195.965 236.155 196.135 ;
        RECT 108.630 194.810 153.130 194.980 ;
        RECT 162.180 194.875 163.390 195.965 ;
        RECT 163.560 195.530 168.905 195.965 ;
        RECT 169.080 195.530 174.425 195.965 ;
        RECT 108.630 185.050 108.800 194.810 ;
        RECT 109.585 194.120 110.585 194.290 ;
        RECT 110.875 194.120 111.875 194.290 ;
        RECT 109.355 185.910 109.525 193.950 ;
        RECT 110.645 185.910 110.815 193.950 ;
        RECT 111.935 185.910 112.105 193.950 ;
        RECT 109.585 185.570 110.585 185.740 ;
        RECT 110.875 185.570 111.875 185.740 ;
        RECT 112.660 185.050 112.830 194.810 ;
        RECT 113.615 194.120 114.615 194.290 ;
        RECT 114.905 194.120 115.905 194.290 ;
        RECT 113.385 185.910 113.555 193.950 ;
        RECT 114.675 185.910 114.845 193.950 ;
        RECT 115.965 185.910 116.135 193.950 ;
        RECT 113.615 185.570 114.615 185.740 ;
        RECT 114.905 185.570 115.905 185.740 ;
        RECT 116.690 185.050 116.860 194.810 ;
        RECT 117.645 194.120 118.645 194.290 ;
        RECT 118.935 194.120 119.935 194.290 ;
        RECT 117.415 185.910 117.585 193.950 ;
        RECT 118.705 185.910 118.875 193.950 ;
        RECT 119.995 185.910 120.165 193.950 ;
        RECT 117.645 185.570 118.645 185.740 ;
        RECT 118.935 185.570 119.935 185.740 ;
        RECT 120.720 185.050 120.890 194.810 ;
        RECT 121.675 194.120 122.675 194.290 ;
        RECT 122.965 194.120 123.965 194.290 ;
        RECT 121.445 185.910 121.615 193.950 ;
        RECT 122.735 185.910 122.905 193.950 ;
        RECT 124.025 185.910 124.195 193.950 ;
        RECT 121.675 185.570 122.675 185.740 ;
        RECT 122.965 185.570 123.965 185.740 ;
        RECT 124.750 185.050 124.920 194.810 ;
        RECT 125.705 194.120 126.705 194.290 ;
        RECT 126.995 194.120 127.995 194.290 ;
        RECT 125.475 185.910 125.645 193.950 ;
        RECT 126.765 185.910 126.935 193.950 ;
        RECT 128.055 185.910 128.225 193.950 ;
        RECT 125.705 185.570 126.705 185.740 ;
        RECT 126.995 185.570 127.995 185.740 ;
        RECT 128.780 185.050 128.950 194.810 ;
        RECT 129.735 194.120 130.735 194.290 ;
        RECT 131.025 194.120 132.025 194.290 ;
        RECT 129.505 185.910 129.675 193.950 ;
        RECT 130.795 185.910 130.965 193.950 ;
        RECT 132.085 185.910 132.255 193.950 ;
        RECT 129.735 185.570 130.735 185.740 ;
        RECT 131.025 185.570 132.025 185.740 ;
        RECT 132.810 185.050 132.980 194.810 ;
        RECT 133.765 194.120 134.765 194.290 ;
        RECT 135.055 194.120 136.055 194.290 ;
        RECT 133.535 185.910 133.705 193.950 ;
        RECT 134.825 185.910 134.995 193.950 ;
        RECT 136.115 185.910 136.285 193.950 ;
        RECT 133.765 185.570 134.765 185.740 ;
        RECT 135.055 185.570 136.055 185.740 ;
        RECT 136.840 185.050 137.010 194.810 ;
        RECT 137.795 194.120 138.795 194.290 ;
        RECT 139.085 194.120 140.085 194.290 ;
        RECT 137.565 185.910 137.735 193.950 ;
        RECT 138.855 185.910 139.025 193.950 ;
        RECT 140.145 185.910 140.315 193.950 ;
        RECT 137.795 185.570 138.795 185.740 ;
        RECT 139.085 185.570 140.085 185.740 ;
        RECT 140.870 185.050 141.040 194.810 ;
        RECT 141.825 194.120 142.825 194.290 ;
        RECT 143.115 194.120 144.115 194.290 ;
        RECT 141.595 185.910 141.765 193.950 ;
        RECT 142.885 185.910 143.055 193.950 ;
        RECT 144.175 185.910 144.345 193.950 ;
        RECT 141.825 185.570 142.825 185.740 ;
        RECT 143.115 185.570 144.115 185.740 ;
        RECT 144.900 185.050 145.070 194.810 ;
        RECT 145.855 194.120 146.855 194.290 ;
        RECT 147.145 194.120 148.145 194.290 ;
        RECT 145.625 185.910 145.795 193.950 ;
        RECT 146.915 185.910 147.085 193.950 ;
        RECT 148.205 185.910 148.375 193.950 ;
        RECT 145.855 185.570 146.855 185.740 ;
        RECT 147.145 185.570 148.145 185.740 ;
        RECT 148.930 185.050 149.100 194.810 ;
        RECT 149.885 194.120 150.885 194.290 ;
        RECT 151.175 194.120 152.175 194.290 ;
        RECT 149.655 185.910 149.825 193.950 ;
        RECT 150.945 185.910 151.115 193.950 ;
        RECT 152.235 185.910 152.405 193.950 ;
        RECT 149.885 185.570 150.885 185.740 ;
        RECT 151.175 185.570 152.175 185.740 ;
        RECT 152.960 185.050 153.130 194.810 ;
        RECT 162.180 194.165 162.700 194.705 ;
        RECT 162.870 194.335 163.390 194.875 ;
        RECT 162.180 193.415 163.390 194.165 ;
        RECT 165.145 193.960 165.485 194.790 ;
        RECT 166.965 194.280 167.315 195.530 ;
        RECT 170.665 193.960 171.005 194.790 ;
        RECT 172.485 194.280 172.835 195.530 ;
        RECT 175.060 194.800 175.350 195.965 ;
        RECT 175.580 194.825 175.790 195.965 ;
        RECT 175.960 194.815 176.290 195.795 ;
        RECT 176.460 194.825 176.690 195.965 ;
        RECT 176.900 195.530 182.245 195.965 ;
        RECT 182.420 195.530 187.765 195.965 ;
        RECT 187.940 195.530 193.285 195.965 ;
        RECT 193.460 195.530 198.805 195.965 ;
        RECT 163.560 193.415 168.905 193.960 ;
        RECT 169.080 193.415 174.425 193.960 ;
        RECT 175.060 193.415 175.350 194.140 ;
        RECT 175.580 193.415 175.790 194.235 ;
        RECT 175.960 194.215 176.210 194.815 ;
        RECT 176.380 194.405 176.710 194.655 ;
        RECT 175.960 193.585 176.290 194.215 ;
        RECT 176.460 193.415 176.690 194.235 ;
        RECT 178.485 193.960 178.825 194.790 ;
        RECT 180.305 194.280 180.655 195.530 ;
        RECT 184.005 193.960 184.345 194.790 ;
        RECT 185.825 194.280 186.175 195.530 ;
        RECT 189.525 193.960 189.865 194.790 ;
        RECT 191.345 194.280 191.695 195.530 ;
        RECT 195.045 193.960 195.385 194.790 ;
        RECT 196.865 194.280 197.215 195.530 ;
        RECT 198.980 194.875 200.650 195.965 ;
        RECT 198.980 194.185 199.730 194.705 ;
        RECT 199.900 194.355 200.650 194.875 ;
        RECT 200.820 194.800 201.110 195.965 ;
        RECT 201.280 195.530 206.625 195.965 ;
        RECT 206.800 195.530 212.145 195.965 ;
        RECT 212.320 195.530 217.665 195.965 ;
        RECT 217.840 195.530 223.185 195.965 ;
        RECT 176.900 193.415 182.245 193.960 ;
        RECT 182.420 193.415 187.765 193.960 ;
        RECT 187.940 193.415 193.285 193.960 ;
        RECT 193.460 193.415 198.805 193.960 ;
        RECT 198.980 193.415 200.650 194.185 ;
        RECT 200.820 193.415 201.110 194.140 ;
        RECT 202.865 193.960 203.205 194.790 ;
        RECT 204.685 194.280 205.035 195.530 ;
        RECT 208.385 193.960 208.725 194.790 ;
        RECT 210.205 194.280 210.555 195.530 ;
        RECT 213.905 193.960 214.245 194.790 ;
        RECT 215.725 194.280 216.075 195.530 ;
        RECT 219.425 193.960 219.765 194.790 ;
        RECT 221.245 194.280 221.595 195.530 ;
        RECT 223.360 194.875 225.950 195.965 ;
        RECT 223.360 194.185 224.570 194.705 ;
        RECT 224.740 194.355 225.950 194.875 ;
        RECT 226.580 194.800 226.870 195.965 ;
        RECT 227.040 195.530 232.385 195.965 ;
        RECT 201.280 193.415 206.625 193.960 ;
        RECT 206.800 193.415 212.145 193.960 ;
        RECT 212.320 193.415 217.665 193.960 ;
        RECT 217.840 193.415 223.185 193.960 ;
        RECT 223.360 193.415 225.950 194.185 ;
        RECT 226.580 193.415 226.870 194.140 ;
        RECT 228.625 193.960 228.965 194.790 ;
        RECT 230.445 194.280 230.795 195.530 ;
        RECT 232.560 194.875 234.230 195.965 ;
        RECT 232.560 194.185 233.310 194.705 ;
        RECT 233.480 194.355 234.230 194.875 ;
        RECT 234.860 194.875 236.070 195.965 ;
        RECT 234.860 194.335 235.380 194.875 ;
        RECT 227.040 193.415 232.385 193.960 ;
        RECT 232.560 193.415 234.230 194.185 ;
        RECT 235.550 194.165 236.070 194.705 ;
        RECT 234.860 193.415 236.070 194.165 ;
        RECT 162.095 193.245 236.155 193.415 ;
        RECT 162.180 192.495 163.390 193.245 ;
        RECT 163.560 192.700 168.905 193.245 ;
        RECT 162.180 191.955 162.700 192.495 ;
        RECT 162.870 191.785 163.390 192.325 ;
        RECT 165.145 191.870 165.485 192.700 ;
        RECT 170.000 192.570 170.260 193.075 ;
        RECT 170.440 192.865 170.770 193.245 ;
        RECT 170.950 192.695 171.120 193.075 ;
        RECT 171.385 192.845 171.720 193.245 ;
        RECT 162.180 190.695 163.390 191.785 ;
        RECT 166.965 191.130 167.315 192.380 ;
        RECT 170.000 191.770 170.170 192.570 ;
        RECT 170.455 192.525 171.120 192.695 ;
        RECT 171.890 192.675 172.095 193.075 ;
        RECT 172.305 192.765 172.580 193.245 ;
        RECT 172.790 192.745 173.050 193.075 ;
        RECT 170.455 192.270 170.625 192.525 ;
        RECT 171.410 192.505 172.095 192.675 ;
        RECT 170.340 191.940 170.625 192.270 ;
        RECT 170.860 191.975 171.190 192.345 ;
        RECT 170.455 191.795 170.625 191.940 ;
        RECT 163.560 190.695 168.905 191.130 ;
        RECT 170.000 190.865 170.270 191.770 ;
        RECT 170.455 191.625 171.120 191.795 ;
        RECT 170.440 190.695 170.770 191.455 ;
        RECT 170.950 190.865 171.120 191.625 ;
        RECT 171.410 191.475 171.750 192.505 ;
        RECT 171.920 191.835 172.170 192.335 ;
        RECT 172.350 192.005 172.710 192.585 ;
        RECT 172.880 191.835 173.050 192.745 ;
        RECT 173.225 192.405 173.485 193.245 ;
        RECT 173.660 192.500 173.915 193.075 ;
        RECT 174.085 192.865 174.415 193.245 ;
        RECT 174.630 192.695 174.800 193.075 ;
        RECT 174.085 192.525 174.800 192.695 ;
        RECT 175.060 192.745 175.360 193.075 ;
        RECT 175.530 192.765 175.805 193.245 ;
        RECT 171.920 191.665 173.050 191.835 ;
        RECT 171.410 191.300 172.075 191.475 ;
        RECT 171.385 190.695 171.720 191.120 ;
        RECT 171.890 190.895 172.075 191.300 ;
        RECT 172.280 190.695 172.610 191.475 ;
        RECT 172.780 190.895 173.050 191.665 ;
        RECT 173.225 190.695 173.485 191.845 ;
        RECT 173.660 191.770 173.830 192.500 ;
        RECT 174.085 192.335 174.255 192.525 ;
        RECT 174.000 192.005 174.255 192.335 ;
        RECT 174.085 191.795 174.255 192.005 ;
        RECT 174.535 191.975 174.890 192.345 ;
        RECT 175.060 191.835 175.230 192.745 ;
        RECT 175.985 192.595 176.280 192.985 ;
        RECT 176.450 192.765 176.705 193.245 ;
        RECT 176.880 192.595 177.140 192.985 ;
        RECT 177.310 192.765 177.590 193.245 ;
        RECT 177.910 192.695 178.080 193.075 ;
        RECT 178.295 192.865 178.625 193.245 ;
        RECT 175.400 192.005 175.750 192.575 ;
        RECT 175.985 192.425 177.635 192.595 ;
        RECT 177.910 192.525 178.625 192.695 ;
        RECT 175.920 192.085 177.060 192.255 ;
        RECT 175.920 191.835 176.090 192.085 ;
        RECT 177.230 191.915 177.635 192.425 ;
        RECT 177.820 191.975 178.175 192.345 ;
        RECT 178.455 192.335 178.625 192.525 ;
        RECT 178.795 192.500 179.050 193.075 ;
        RECT 178.455 192.005 178.710 192.335 ;
        RECT 173.660 190.865 173.915 191.770 ;
        RECT 174.085 191.625 174.800 191.795 ;
        RECT 174.085 190.695 174.415 191.455 ;
        RECT 174.630 190.865 174.800 191.625 ;
        RECT 175.060 191.665 176.090 191.835 ;
        RECT 176.880 191.745 177.635 191.915 ;
        RECT 178.455 191.795 178.625 192.005 ;
        RECT 175.060 190.865 175.370 191.665 ;
        RECT 176.880 191.495 177.140 191.745 ;
        RECT 177.910 191.625 178.625 191.795 ;
        RECT 178.880 191.770 179.050 192.500 ;
        RECT 179.225 192.405 179.485 193.245 ;
        RECT 179.660 192.570 179.920 193.075 ;
        RECT 180.100 192.865 180.430 193.245 ;
        RECT 180.610 192.695 180.780 193.075 ;
        RECT 175.540 190.695 175.850 191.495 ;
        RECT 176.020 191.325 177.140 191.495 ;
        RECT 176.020 190.865 176.280 191.325 ;
        RECT 176.450 190.695 176.705 191.155 ;
        RECT 176.880 190.865 177.140 191.325 ;
        RECT 177.310 190.695 177.595 191.565 ;
        RECT 177.910 190.865 178.080 191.625 ;
        RECT 178.295 190.695 178.625 191.455 ;
        RECT 178.795 190.865 179.050 191.770 ;
        RECT 179.225 190.695 179.485 191.845 ;
        RECT 179.660 191.770 179.830 192.570 ;
        RECT 180.115 192.525 180.780 192.695 ;
        RECT 180.115 192.270 180.285 192.525 ;
        RECT 181.040 192.475 184.550 193.245 ;
        RECT 180.000 191.940 180.285 192.270 ;
        RECT 180.520 191.975 180.850 192.345 ;
        RECT 181.040 191.955 182.690 192.475 ;
        RECT 180.115 191.795 180.285 191.940 ;
        RECT 179.660 190.865 179.930 191.770 ;
        RECT 180.115 191.625 180.780 191.795 ;
        RECT 182.860 191.785 184.550 192.305 ;
        RECT 180.100 190.695 180.430 191.455 ;
        RECT 180.610 190.865 180.780 191.625 ;
        RECT 181.040 190.695 184.550 191.785 ;
        RECT 184.720 192.300 185.060 193.075 ;
        RECT 185.230 192.785 185.400 193.245 ;
        RECT 185.640 192.810 186.000 193.075 ;
        RECT 185.640 192.805 185.995 192.810 ;
        RECT 185.640 192.795 185.990 192.805 ;
        RECT 185.640 192.790 185.985 192.795 ;
        RECT 185.640 192.780 185.980 192.790 ;
        RECT 186.630 192.785 186.800 193.245 ;
        RECT 185.640 192.775 185.975 192.780 ;
        RECT 185.640 192.765 185.965 192.775 ;
        RECT 185.640 192.755 185.955 192.765 ;
        RECT 185.640 192.615 185.940 192.755 ;
        RECT 185.230 192.425 185.940 192.615 ;
        RECT 186.130 192.615 186.460 192.695 ;
        RECT 186.970 192.615 187.310 193.075 ;
        RECT 186.130 192.425 187.310 192.615 ;
        RECT 187.940 192.520 188.230 193.245 ;
        RECT 188.400 192.700 193.745 193.245 ;
        RECT 184.720 190.865 185.000 192.300 ;
        RECT 185.230 191.855 185.515 192.425 ;
        RECT 185.700 192.025 186.170 192.255 ;
        RECT 186.340 192.235 186.670 192.255 ;
        RECT 186.340 192.055 186.790 192.235 ;
        RECT 186.980 192.055 187.310 192.255 ;
        RECT 185.230 191.640 186.380 191.855 ;
        RECT 185.170 190.695 185.880 191.470 ;
        RECT 186.050 190.865 186.380 191.640 ;
        RECT 186.575 190.940 186.790 192.055 ;
        RECT 187.080 191.715 187.310 192.055 ;
        RECT 189.985 191.870 190.325 192.700 ;
        RECT 186.970 190.695 187.300 191.415 ;
        RECT 187.940 190.695 188.230 191.860 ;
        RECT 191.805 191.130 192.155 192.380 ;
        RECT 194.380 192.300 194.720 193.075 ;
        RECT 194.890 192.785 195.060 193.245 ;
        RECT 195.300 192.810 195.660 193.075 ;
        RECT 195.300 192.805 195.655 192.810 ;
        RECT 195.300 192.795 195.650 192.805 ;
        RECT 195.300 192.790 195.645 192.795 ;
        RECT 195.300 192.780 195.640 192.790 ;
        RECT 196.290 192.785 196.460 193.245 ;
        RECT 195.300 192.775 195.635 192.780 ;
        RECT 195.300 192.765 195.625 192.775 ;
        RECT 195.300 192.755 195.615 192.765 ;
        RECT 195.300 192.615 195.600 192.755 ;
        RECT 194.890 192.425 195.600 192.615 ;
        RECT 195.790 192.615 196.120 192.695 ;
        RECT 196.630 192.615 196.970 193.075 ;
        RECT 195.790 192.425 196.970 192.615 ;
        RECT 197.140 192.475 200.650 193.245 ;
        RECT 200.820 192.495 202.030 193.245 ;
        RECT 202.200 192.615 202.540 193.075 ;
        RECT 202.710 192.785 202.880 193.245 ;
        RECT 203.510 192.810 203.870 193.075 ;
        RECT 203.515 192.805 203.870 192.810 ;
        RECT 203.520 192.795 203.870 192.805 ;
        RECT 203.525 192.790 203.870 192.795 ;
        RECT 203.530 192.780 203.870 192.790 ;
        RECT 204.110 192.785 204.280 193.245 ;
        RECT 203.535 192.775 203.870 192.780 ;
        RECT 203.545 192.765 203.870 192.775 ;
        RECT 203.555 192.755 203.870 192.765 ;
        RECT 203.050 192.615 203.380 192.695 ;
        RECT 188.400 190.695 193.745 191.130 ;
        RECT 194.380 190.865 194.660 192.300 ;
        RECT 194.890 191.855 195.175 192.425 ;
        RECT 195.360 192.025 195.830 192.255 ;
        RECT 196.000 192.235 196.330 192.255 ;
        RECT 196.000 192.055 196.450 192.235 ;
        RECT 196.640 192.055 196.970 192.255 ;
        RECT 194.890 191.640 196.040 191.855 ;
        RECT 194.830 190.695 195.540 191.470 ;
        RECT 195.710 190.865 196.040 191.640 ;
        RECT 196.235 190.940 196.450 192.055 ;
        RECT 196.740 191.715 196.970 192.055 ;
        RECT 197.140 191.955 198.790 192.475 ;
        RECT 198.960 191.785 200.650 192.305 ;
        RECT 200.820 191.955 201.340 192.495 ;
        RECT 202.200 192.425 203.380 192.615 ;
        RECT 203.570 192.615 203.870 192.755 ;
        RECT 203.570 192.425 204.280 192.615 ;
        RECT 201.510 191.785 202.030 192.325 ;
        RECT 196.630 190.695 196.960 191.415 ;
        RECT 197.140 190.695 200.650 191.785 ;
        RECT 200.820 190.695 202.030 191.785 ;
        RECT 202.200 192.055 202.530 192.255 ;
        RECT 202.840 192.235 203.170 192.255 ;
        RECT 202.720 192.055 203.170 192.235 ;
        RECT 202.200 191.715 202.430 192.055 ;
        RECT 202.210 190.695 202.540 191.415 ;
        RECT 202.720 190.940 202.935 192.055 ;
        RECT 203.340 192.025 203.810 192.255 ;
        RECT 203.995 191.855 204.280 192.425 ;
        RECT 204.450 192.300 204.790 193.075 ;
        RECT 204.960 192.700 210.305 193.245 ;
        RECT 203.130 191.640 204.280 191.855 ;
        RECT 203.130 190.865 203.460 191.640 ;
        RECT 203.630 190.695 204.340 191.470 ;
        RECT 204.510 190.865 204.790 192.300 ;
        RECT 206.545 191.870 206.885 192.700 ;
        RECT 210.480 192.475 213.070 193.245 ;
        RECT 213.700 192.520 213.990 193.245 ;
        RECT 214.160 192.700 219.505 193.245 ;
        RECT 219.680 192.700 225.025 193.245 ;
        RECT 225.200 192.700 230.545 193.245 ;
        RECT 208.365 191.130 208.715 192.380 ;
        RECT 210.480 191.955 211.690 192.475 ;
        RECT 211.860 191.785 213.070 192.305 ;
        RECT 215.745 191.870 216.085 192.700 ;
        RECT 204.960 190.695 210.305 191.130 ;
        RECT 210.480 190.695 213.070 191.785 ;
        RECT 213.700 190.695 213.990 191.860 ;
        RECT 217.565 191.130 217.915 192.380 ;
        RECT 221.265 191.870 221.605 192.700 ;
        RECT 223.085 191.130 223.435 192.380 ;
        RECT 226.785 191.870 227.125 192.700 ;
        RECT 230.720 192.475 234.230 193.245 ;
        RECT 234.860 192.495 236.070 193.245 ;
        RECT 228.605 191.130 228.955 192.380 ;
        RECT 230.720 191.955 232.370 192.475 ;
        RECT 232.540 191.785 234.230 192.305 ;
        RECT 214.160 190.695 219.505 191.130 ;
        RECT 219.680 190.695 225.025 191.130 ;
        RECT 225.200 190.695 230.545 191.130 ;
        RECT 230.720 190.695 234.230 191.785 ;
        RECT 234.860 191.785 235.380 192.325 ;
        RECT 235.550 191.955 236.070 192.495 ;
        RECT 234.860 190.695 236.070 191.785 ;
        RECT 162.095 190.525 236.155 190.695 ;
        RECT 162.180 189.435 163.390 190.525 ;
        RECT 162.180 188.725 162.700 189.265 ;
        RECT 162.870 188.895 163.390 189.435 ;
        RECT 163.650 189.595 163.820 190.355 ;
        RECT 164.000 189.765 164.330 190.525 ;
        RECT 163.650 189.425 164.315 189.595 ;
        RECT 164.500 189.450 164.770 190.355 ;
        RECT 164.145 189.280 164.315 189.425 ;
        RECT 163.580 188.875 163.910 189.245 ;
        RECT 164.145 188.950 164.430 189.280 ;
        RECT 162.180 187.975 163.390 188.725 ;
        RECT 164.145 188.695 164.315 188.950 ;
        RECT 163.650 188.525 164.315 188.695 ;
        RECT 164.600 188.650 164.770 189.450 ;
        RECT 164.940 189.435 166.610 190.525 ;
        RECT 163.650 188.145 163.820 188.525 ;
        RECT 164.000 187.975 164.330 188.355 ;
        RECT 164.510 188.145 164.770 188.650 ;
        RECT 164.940 188.745 165.690 189.265 ;
        RECT 165.860 188.915 166.610 189.435 ;
        RECT 166.870 189.595 167.040 190.355 ;
        RECT 167.220 189.765 167.550 190.525 ;
        RECT 166.870 189.425 167.535 189.595 ;
        RECT 167.720 189.450 167.990 190.355 ;
        RECT 167.365 189.280 167.535 189.425 ;
        RECT 166.800 188.875 167.130 189.245 ;
        RECT 167.365 188.950 167.650 189.280 ;
        RECT 164.940 187.975 166.610 188.745 ;
        RECT 167.365 188.695 167.535 188.950 ;
        RECT 166.870 188.525 167.535 188.695 ;
        RECT 167.820 188.650 167.990 189.450 ;
        RECT 168.250 189.595 168.420 190.355 ;
        RECT 168.600 189.765 168.930 190.525 ;
        RECT 168.250 189.425 168.915 189.595 ;
        RECT 169.100 189.450 169.370 190.355 ;
        RECT 169.545 190.100 169.880 190.525 ;
        RECT 170.050 189.920 170.235 190.325 ;
        RECT 168.745 189.280 168.915 189.425 ;
        RECT 168.180 188.875 168.510 189.245 ;
        RECT 168.745 188.950 169.030 189.280 ;
        RECT 168.745 188.695 168.915 188.950 ;
        RECT 166.870 188.145 167.040 188.525 ;
        RECT 167.220 187.975 167.550 188.355 ;
        RECT 167.730 188.145 167.990 188.650 ;
        RECT 168.250 188.525 168.915 188.695 ;
        RECT 169.200 188.650 169.370 189.450 ;
        RECT 168.250 188.145 168.420 188.525 ;
        RECT 168.600 187.975 168.930 188.355 ;
        RECT 169.110 188.145 169.370 188.650 ;
        RECT 169.570 189.745 170.235 189.920 ;
        RECT 170.440 189.745 170.770 190.525 ;
        RECT 169.570 188.715 169.910 189.745 ;
        RECT 170.940 189.555 171.210 190.325 ;
        RECT 170.080 189.385 171.210 189.555 ;
        RECT 171.595 189.425 171.925 190.525 ;
        RECT 172.400 189.925 172.725 190.355 ;
        RECT 172.895 190.105 173.225 190.525 ;
        RECT 173.970 190.095 174.380 190.525 ;
        RECT 172.400 189.755 174.380 189.925 ;
        RECT 170.080 188.885 170.330 189.385 ;
        RECT 169.570 188.545 170.255 188.715 ;
        RECT 170.510 188.635 170.870 189.215 ;
        RECT 169.545 187.975 169.880 188.375 ;
        RECT 170.050 188.145 170.255 188.545 ;
        RECT 171.040 188.475 171.210 189.385 ;
        RECT 172.400 189.345 173.105 189.755 ;
        RECT 171.380 188.965 172.025 189.175 ;
        RECT 172.195 188.965 172.765 189.175 ;
        RECT 170.465 187.975 170.740 188.455 ;
        RECT 170.950 188.145 171.210 188.475 ;
        RECT 171.535 188.625 172.705 188.795 ;
        RECT 171.535 188.160 171.865 188.625 ;
        RECT 172.035 187.975 172.205 188.445 ;
        RECT 172.375 188.145 172.705 188.625 ;
        RECT 172.935 188.145 173.105 189.345 ;
        RECT 173.275 189.415 173.900 189.585 ;
        RECT 173.275 188.715 173.445 189.415 ;
        RECT 174.115 189.215 174.380 189.755 ;
        RECT 174.550 189.370 174.890 190.355 ;
        RECT 173.615 188.885 173.945 189.215 ;
        RECT 174.115 188.885 174.465 189.215 ;
        RECT 174.635 188.715 174.890 189.370 ;
        RECT 175.060 189.360 175.350 190.525 ;
        RECT 175.735 189.425 176.065 190.525 ;
        RECT 176.540 189.925 176.865 190.355 ;
        RECT 177.035 190.105 177.365 190.525 ;
        RECT 178.110 190.095 178.520 190.525 ;
        RECT 176.540 189.755 178.520 189.925 ;
        RECT 176.540 189.345 177.245 189.755 ;
        RECT 175.520 188.965 176.165 189.175 ;
        RECT 176.335 188.965 176.905 189.175 ;
        RECT 173.275 188.545 173.815 188.715 ;
        RECT 173.645 188.340 173.815 188.545 ;
        RECT 174.095 187.975 174.265 188.715 ;
        RECT 174.530 188.340 174.890 188.715 ;
        RECT 175.060 187.975 175.350 188.700 ;
        RECT 175.675 188.625 176.845 188.795 ;
        RECT 175.675 188.160 176.005 188.625 ;
        RECT 176.175 187.975 176.345 188.445 ;
        RECT 176.515 188.145 176.845 188.625 ;
        RECT 177.075 188.145 177.245 189.345 ;
        RECT 177.415 189.415 178.040 189.585 ;
        RECT 177.415 188.715 177.585 189.415 ;
        RECT 178.255 189.215 178.520 189.755 ;
        RECT 178.690 189.370 179.030 190.355 ;
        RECT 177.755 188.885 178.085 189.215 ;
        RECT 178.255 188.885 178.605 189.215 ;
        RECT 178.775 188.715 179.030 189.370 ;
        RECT 179.750 189.515 179.920 190.355 ;
        RECT 180.090 190.185 181.260 190.355 ;
        RECT 180.090 189.685 180.420 190.185 ;
        RECT 180.930 190.145 181.260 190.185 ;
        RECT 181.450 190.105 181.805 190.525 ;
        RECT 180.590 189.925 180.820 190.015 ;
        RECT 181.975 189.925 182.225 190.355 ;
        RECT 180.590 189.685 182.225 189.925 ;
        RECT 182.395 189.765 182.725 190.525 ;
        RECT 182.895 189.685 183.150 190.355 ;
        RECT 183.835 189.725 184.085 190.525 ;
        RECT 184.255 189.895 184.585 190.355 ;
        RECT 184.755 190.065 184.970 190.525 ;
        RECT 184.255 189.725 185.425 189.895 ;
        RECT 182.940 189.675 183.150 189.685 ;
        RECT 179.750 189.345 182.810 189.515 ;
        RECT 179.665 188.965 180.015 189.175 ;
        RECT 180.185 188.965 180.630 189.165 ;
        RECT 180.800 188.965 181.275 189.165 ;
        RECT 177.415 188.545 177.955 188.715 ;
        RECT 177.785 188.340 177.955 188.545 ;
        RECT 178.235 187.975 178.405 188.715 ;
        RECT 178.670 188.340 179.030 188.715 ;
        RECT 179.750 188.625 180.815 188.795 ;
        RECT 179.750 188.145 179.920 188.625 ;
        RECT 180.090 187.975 180.420 188.455 ;
        RECT 180.645 188.395 180.815 188.625 ;
        RECT 180.995 188.565 181.275 188.965 ;
        RECT 181.545 188.965 181.875 189.165 ;
        RECT 182.045 188.995 182.420 189.165 ;
        RECT 182.045 188.965 182.410 188.995 ;
        RECT 181.545 188.565 181.830 188.965 ;
        RECT 182.640 188.795 182.810 189.345 ;
        RECT 182.010 188.625 182.810 188.795 ;
        RECT 182.010 188.395 182.180 188.625 ;
        RECT 182.980 188.555 183.150 189.675 ;
        RECT 183.345 189.555 183.625 189.715 ;
        RECT 183.345 189.385 184.680 189.555 ;
        RECT 184.510 189.215 184.680 189.385 ;
        RECT 183.345 188.965 183.695 189.205 ;
        RECT 183.865 188.965 184.340 189.205 ;
        RECT 184.510 188.965 184.885 189.215 ;
        RECT 184.510 188.795 184.680 188.965 ;
        RECT 182.965 188.475 183.150 188.555 ;
        RECT 180.645 188.145 182.180 188.395 ;
        RECT 182.350 187.975 182.680 188.455 ;
        RECT 182.895 188.145 183.150 188.475 ;
        RECT 183.345 188.625 184.680 188.795 ;
        RECT 183.345 188.415 183.615 188.625 ;
        RECT 185.055 188.435 185.425 189.725 ;
        RECT 186.190 189.515 186.360 190.355 ;
        RECT 186.530 190.185 187.700 190.355 ;
        RECT 186.530 189.685 186.860 190.185 ;
        RECT 187.370 190.145 187.700 190.185 ;
        RECT 187.890 190.105 188.245 190.525 ;
        RECT 187.030 189.925 187.260 190.015 ;
        RECT 188.415 189.925 188.665 190.355 ;
        RECT 187.030 189.685 188.665 189.925 ;
        RECT 188.835 189.765 189.165 190.525 ;
        RECT 189.335 189.685 189.590 190.355 ;
        RECT 190.735 189.725 190.985 190.525 ;
        RECT 191.155 189.895 191.485 190.355 ;
        RECT 191.655 190.065 191.870 190.525 ;
        RECT 191.155 189.725 192.325 189.895 ;
        RECT 186.190 189.345 189.250 189.515 ;
        RECT 186.105 188.965 186.455 189.175 ;
        RECT 186.625 188.965 187.070 189.165 ;
        RECT 187.240 188.965 187.715 189.165 ;
        RECT 183.835 187.975 184.165 188.435 ;
        RECT 184.675 188.145 185.425 188.435 ;
        RECT 186.190 188.625 187.255 188.795 ;
        RECT 186.190 188.145 186.360 188.625 ;
        RECT 186.530 187.975 186.860 188.455 ;
        RECT 187.085 188.395 187.255 188.625 ;
        RECT 187.435 188.565 187.715 188.965 ;
        RECT 187.985 188.965 188.315 189.165 ;
        RECT 188.485 188.995 188.860 189.165 ;
        RECT 188.485 188.965 188.850 188.995 ;
        RECT 187.985 188.565 188.270 188.965 ;
        RECT 189.080 188.795 189.250 189.345 ;
        RECT 188.450 188.625 189.250 188.795 ;
        RECT 188.450 188.395 188.620 188.625 ;
        RECT 189.420 188.555 189.590 189.685 ;
        RECT 190.245 189.555 190.525 189.715 ;
        RECT 190.245 189.385 191.580 189.555 ;
        RECT 191.410 189.215 191.580 189.385 ;
        RECT 190.245 188.965 190.595 189.205 ;
        RECT 190.765 188.965 191.240 189.205 ;
        RECT 191.410 188.965 191.785 189.215 ;
        RECT 191.410 188.795 191.580 188.965 ;
        RECT 189.405 188.475 189.590 188.555 ;
        RECT 187.085 188.145 188.620 188.395 ;
        RECT 188.790 187.975 189.120 188.455 ;
        RECT 189.335 188.145 189.590 188.475 ;
        RECT 190.245 188.625 191.580 188.795 ;
        RECT 190.245 188.415 190.515 188.625 ;
        RECT 191.955 188.435 192.325 189.725 ;
        RECT 192.540 189.435 195.130 190.525 ;
        RECT 190.735 187.975 191.065 188.435 ;
        RECT 191.575 188.145 192.325 188.435 ;
        RECT 192.540 188.745 193.750 189.265 ;
        RECT 193.920 188.915 195.130 189.435 ;
        RECT 195.765 189.385 196.100 190.355 ;
        RECT 196.270 189.385 196.440 190.525 ;
        RECT 196.610 190.185 198.640 190.355 ;
        RECT 192.540 187.975 195.130 188.745 ;
        RECT 195.765 188.715 195.935 189.385 ;
        RECT 196.610 189.215 196.780 190.185 ;
        RECT 196.105 188.885 196.360 189.215 ;
        RECT 196.585 188.885 196.780 189.215 ;
        RECT 196.950 189.845 198.075 190.015 ;
        RECT 196.190 188.715 196.360 188.885 ;
        RECT 196.950 188.715 197.120 189.845 ;
        RECT 195.765 188.145 196.020 188.715 ;
        RECT 196.190 188.545 197.120 188.715 ;
        RECT 197.290 189.505 198.300 189.675 ;
        RECT 197.290 188.705 197.460 189.505 ;
        RECT 197.665 189.165 197.940 189.305 ;
        RECT 197.660 188.995 197.940 189.165 ;
        RECT 196.945 188.510 197.120 188.545 ;
        RECT 196.190 187.975 196.520 188.375 ;
        RECT 196.945 188.145 197.475 188.510 ;
        RECT 197.665 188.145 197.940 188.995 ;
        RECT 198.110 188.145 198.300 189.505 ;
        RECT 198.470 189.520 198.640 190.185 ;
        RECT 198.810 189.765 198.980 190.525 ;
        RECT 199.215 189.765 199.730 190.175 ;
        RECT 198.470 189.330 199.220 189.520 ;
        RECT 199.390 188.955 199.730 189.765 ;
        RECT 200.820 189.360 201.110 190.525 ;
        RECT 201.280 190.090 206.625 190.525 ;
        RECT 198.500 188.785 199.730 188.955 ;
        RECT 198.480 187.975 198.990 188.510 ;
        RECT 199.210 188.180 199.455 188.785 ;
        RECT 200.820 187.975 201.110 188.700 ;
        RECT 202.865 188.520 203.205 189.350 ;
        RECT 204.685 188.840 205.035 190.090 ;
        RECT 206.800 189.435 210.310 190.525 ;
        RECT 211.410 189.805 211.740 190.525 ;
        RECT 206.800 188.745 208.450 189.265 ;
        RECT 208.620 188.915 210.310 189.435 ;
        RECT 211.400 189.165 211.630 189.505 ;
        RECT 211.920 189.165 212.135 190.280 ;
        RECT 212.330 189.580 212.660 190.355 ;
        RECT 212.830 189.750 213.540 190.525 ;
        RECT 212.330 189.365 213.480 189.580 ;
        RECT 211.400 188.965 211.730 189.165 ;
        RECT 211.920 188.985 212.370 189.165 ;
        RECT 212.040 188.965 212.370 188.985 ;
        RECT 212.540 188.965 213.010 189.195 ;
        RECT 213.195 188.795 213.480 189.365 ;
        RECT 213.710 188.920 213.990 190.355 ;
        RECT 214.160 190.090 219.505 190.525 ;
        RECT 201.280 187.975 206.625 188.520 ;
        RECT 206.800 187.975 210.310 188.745 ;
        RECT 211.400 188.605 212.580 188.795 ;
        RECT 211.400 188.145 211.740 188.605 ;
        RECT 212.250 188.525 212.580 188.605 ;
        RECT 212.770 188.605 213.480 188.795 ;
        RECT 212.770 188.465 213.070 188.605 ;
        RECT 212.755 188.455 213.070 188.465 ;
        RECT 212.745 188.445 213.070 188.455 ;
        RECT 212.735 188.440 213.070 188.445 ;
        RECT 211.910 187.975 212.080 188.435 ;
        RECT 212.730 188.430 213.070 188.440 ;
        RECT 212.725 188.425 213.070 188.430 ;
        RECT 212.720 188.415 213.070 188.425 ;
        RECT 212.715 188.410 213.070 188.415 ;
        RECT 212.710 188.145 213.070 188.410 ;
        RECT 213.310 187.975 213.480 188.435 ;
        RECT 213.650 188.145 213.990 188.920 ;
        RECT 215.745 188.520 216.085 189.350 ;
        RECT 217.565 188.840 217.915 190.090 ;
        RECT 219.680 189.435 222.270 190.525 ;
        RECT 219.680 188.745 220.890 189.265 ;
        RECT 221.060 188.915 222.270 189.435 ;
        RECT 222.900 188.920 223.180 190.355 ;
        RECT 223.350 189.750 224.060 190.525 ;
        RECT 224.230 189.580 224.560 190.355 ;
        RECT 223.410 189.365 224.560 189.580 ;
        RECT 214.160 187.975 219.505 188.520 ;
        RECT 219.680 187.975 222.270 188.745 ;
        RECT 222.900 188.145 223.240 188.920 ;
        RECT 223.410 188.795 223.695 189.365 ;
        RECT 223.880 188.965 224.350 189.195 ;
        RECT 224.755 189.165 224.970 190.280 ;
        RECT 225.150 189.805 225.480 190.525 ;
        RECT 225.260 189.165 225.490 189.505 ;
        RECT 226.580 189.360 226.870 190.525 ;
        RECT 227.130 189.595 227.300 190.355 ;
        RECT 227.480 189.765 227.810 190.525 ;
        RECT 227.130 189.425 227.795 189.595 ;
        RECT 227.980 189.450 228.250 190.355 ;
        RECT 227.625 189.280 227.795 189.425 ;
        RECT 224.520 188.985 224.970 189.165 ;
        RECT 224.520 188.965 224.850 188.985 ;
        RECT 225.160 188.965 225.490 189.165 ;
        RECT 227.060 188.875 227.390 189.245 ;
        RECT 227.625 188.950 227.910 189.280 ;
        RECT 223.410 188.605 224.120 188.795 ;
        RECT 223.820 188.465 224.120 188.605 ;
        RECT 224.310 188.605 225.490 188.795 ;
        RECT 224.310 188.525 224.640 188.605 ;
        RECT 223.820 188.455 224.135 188.465 ;
        RECT 223.820 188.445 224.145 188.455 ;
        RECT 223.820 188.440 224.155 188.445 ;
        RECT 223.410 187.975 223.580 188.435 ;
        RECT 223.820 188.430 224.160 188.440 ;
        RECT 223.820 188.425 224.165 188.430 ;
        RECT 223.820 188.415 224.170 188.425 ;
        RECT 223.820 188.410 224.175 188.415 ;
        RECT 223.820 188.145 224.180 188.410 ;
        RECT 224.810 187.975 224.980 188.435 ;
        RECT 225.150 188.145 225.490 188.605 ;
        RECT 226.580 187.975 226.870 188.700 ;
        RECT 227.625 188.695 227.795 188.950 ;
        RECT 227.130 188.525 227.795 188.695 ;
        RECT 228.080 188.650 228.250 189.450 ;
        RECT 227.130 188.145 227.300 188.525 ;
        RECT 227.480 187.975 227.810 188.355 ;
        RECT 227.990 188.145 228.250 188.650 ;
        RECT 228.420 189.450 228.690 190.355 ;
        RECT 228.860 189.765 229.190 190.525 ;
        RECT 229.370 189.595 229.540 190.355 ;
        RECT 228.420 188.650 228.590 189.450 ;
        RECT 228.875 189.425 229.540 189.595 ;
        RECT 229.800 189.450 230.070 190.355 ;
        RECT 230.240 189.765 230.570 190.525 ;
        RECT 230.750 189.595 230.920 190.355 ;
        RECT 228.875 189.280 229.045 189.425 ;
        RECT 228.760 188.950 229.045 189.280 ;
        RECT 228.875 188.695 229.045 188.950 ;
        RECT 229.280 188.875 229.610 189.245 ;
        RECT 228.420 188.145 228.680 188.650 ;
        RECT 228.875 188.525 229.540 188.695 ;
        RECT 228.860 187.975 229.190 188.355 ;
        RECT 229.370 188.145 229.540 188.525 ;
        RECT 229.800 188.650 229.970 189.450 ;
        RECT 230.255 189.425 230.920 189.595 ;
        RECT 231.180 189.435 234.690 190.525 ;
        RECT 230.255 189.280 230.425 189.425 ;
        RECT 230.140 188.950 230.425 189.280 ;
        RECT 230.255 188.695 230.425 188.950 ;
        RECT 230.660 188.875 230.990 189.245 ;
        RECT 231.180 188.745 232.830 189.265 ;
        RECT 233.000 188.915 234.690 189.435 ;
        RECT 234.860 189.435 236.070 190.525 ;
        RECT 234.860 188.895 235.380 189.435 ;
        RECT 229.800 188.145 230.060 188.650 ;
        RECT 230.255 188.525 230.920 188.695 ;
        RECT 230.240 187.975 230.570 188.355 ;
        RECT 230.750 188.145 230.920 188.525 ;
        RECT 231.180 187.975 234.690 188.745 ;
        RECT 235.550 188.725 236.070 189.265 ;
        RECT 234.860 187.975 236.070 188.725 ;
        RECT 162.095 187.805 236.155 187.975 ;
        RECT 162.180 187.055 163.390 187.805 ;
        RECT 163.650 187.255 163.820 187.635 ;
        RECT 164.000 187.425 164.330 187.805 ;
        RECT 163.650 187.085 164.315 187.255 ;
        RECT 164.510 187.130 164.770 187.635 ;
        RECT 162.180 186.515 162.700 187.055 ;
        RECT 162.870 186.345 163.390 186.885 ;
        RECT 163.580 186.535 163.910 186.905 ;
        RECT 164.145 186.830 164.315 187.085 ;
        RECT 164.145 186.500 164.430 186.830 ;
        RECT 164.145 186.355 164.315 186.500 ;
        RECT 162.180 185.255 163.390 186.345 ;
        RECT 163.650 186.185 164.315 186.355 ;
        RECT 164.600 186.330 164.770 187.130 ;
        RECT 165.030 187.255 165.200 187.635 ;
        RECT 165.380 187.425 165.710 187.805 ;
        RECT 165.030 187.085 165.695 187.255 ;
        RECT 165.890 187.130 166.150 187.635 ;
        RECT 164.960 186.535 165.290 186.905 ;
        RECT 165.525 186.830 165.695 187.085 ;
        RECT 165.525 186.500 165.810 186.830 ;
        RECT 165.525 186.355 165.695 186.500 ;
        RECT 163.650 185.425 163.820 186.185 ;
        RECT 164.000 185.255 164.330 186.015 ;
        RECT 164.500 185.425 164.770 186.330 ;
        RECT 165.030 186.185 165.695 186.355 ;
        RECT 165.980 186.330 166.150 187.130 ;
        RECT 166.410 187.255 166.580 187.635 ;
        RECT 166.760 187.425 167.090 187.805 ;
        RECT 166.410 187.085 167.075 187.255 ;
        RECT 167.270 187.130 167.530 187.635 ;
        RECT 166.340 186.535 166.670 186.905 ;
        RECT 166.905 186.830 167.075 187.085 ;
        RECT 166.905 186.500 167.190 186.830 ;
        RECT 166.905 186.355 167.075 186.500 ;
        RECT 165.030 185.425 165.200 186.185 ;
        RECT 165.380 185.255 165.710 186.015 ;
        RECT 165.880 185.425 166.150 186.330 ;
        RECT 166.410 186.185 167.075 186.355 ;
        RECT 167.360 186.330 167.530 187.130 ;
        RECT 166.410 185.425 166.580 186.185 ;
        RECT 166.760 185.255 167.090 186.015 ;
        RECT 167.260 185.425 167.530 186.330 ;
        RECT 167.700 186.860 168.040 187.635 ;
        RECT 168.210 187.345 168.380 187.805 ;
        RECT 168.620 187.370 168.980 187.635 ;
        RECT 168.620 187.365 168.975 187.370 ;
        RECT 168.620 187.355 168.970 187.365 ;
        RECT 168.620 187.350 168.965 187.355 ;
        RECT 168.620 187.340 168.960 187.350 ;
        RECT 169.610 187.345 169.780 187.805 ;
        RECT 168.620 187.335 168.955 187.340 ;
        RECT 168.620 187.325 168.945 187.335 ;
        RECT 168.620 187.315 168.935 187.325 ;
        RECT 168.620 187.175 168.920 187.315 ;
        RECT 168.210 186.985 168.920 187.175 ;
        RECT 169.110 187.175 169.440 187.255 ;
        RECT 169.950 187.175 170.290 187.635 ;
        RECT 169.110 186.985 170.290 187.175 ;
        RECT 170.615 187.155 170.945 187.620 ;
        RECT 171.115 187.335 171.285 187.805 ;
        RECT 171.455 187.155 171.785 187.635 ;
        RECT 170.615 186.985 171.785 187.155 ;
        RECT 167.700 185.425 167.980 186.860 ;
        RECT 168.210 186.415 168.495 186.985 ;
        RECT 168.680 186.585 169.150 186.815 ;
        RECT 169.320 186.795 169.650 186.815 ;
        RECT 169.320 186.615 169.770 186.795 ;
        RECT 169.960 186.615 170.290 186.815 ;
        RECT 168.210 186.200 169.360 186.415 ;
        RECT 168.150 185.255 168.860 186.030 ;
        RECT 169.030 185.425 169.360 186.200 ;
        RECT 169.555 185.500 169.770 186.615 ;
        RECT 170.060 186.275 170.290 186.615 ;
        RECT 170.460 186.605 171.105 186.815 ;
        RECT 171.275 186.605 171.845 186.815 ;
        RECT 172.015 186.435 172.185 187.635 ;
        RECT 172.725 187.235 172.895 187.440 ;
        RECT 169.950 185.255 170.280 185.975 ;
        RECT 170.675 185.255 171.005 186.355 ;
        RECT 171.480 186.025 172.185 186.435 ;
        RECT 172.355 187.065 172.895 187.235 ;
        RECT 173.175 187.065 173.345 187.805 ;
        RECT 173.610 187.065 173.970 187.440 ;
        RECT 172.355 186.365 172.525 187.065 ;
        RECT 172.695 186.565 173.025 186.895 ;
        RECT 173.195 186.565 173.545 186.895 ;
        RECT 172.355 186.195 172.980 186.365 ;
        RECT 173.195 186.025 173.460 186.565 ;
        RECT 173.715 186.410 173.970 187.065 ;
        RECT 171.480 185.855 173.460 186.025 ;
        RECT 171.480 185.425 171.805 185.855 ;
        RECT 171.975 185.255 172.305 185.675 ;
        RECT 173.050 185.255 173.460 185.685 ;
        RECT 173.630 185.425 173.970 186.410 ;
        RECT 175.060 186.860 175.400 187.635 ;
        RECT 175.570 187.345 175.740 187.805 ;
        RECT 175.980 187.370 176.340 187.635 ;
        RECT 175.980 187.365 176.335 187.370 ;
        RECT 175.980 187.355 176.330 187.365 ;
        RECT 175.980 187.350 176.325 187.355 ;
        RECT 175.980 187.340 176.320 187.350 ;
        RECT 176.970 187.345 177.140 187.805 ;
        RECT 175.980 187.335 176.315 187.340 ;
        RECT 175.980 187.325 176.305 187.335 ;
        RECT 175.980 187.315 176.295 187.325 ;
        RECT 175.980 187.175 176.280 187.315 ;
        RECT 175.570 186.985 176.280 187.175 ;
        RECT 176.470 187.175 176.800 187.255 ;
        RECT 177.310 187.175 177.650 187.635 ;
        RECT 176.470 186.985 177.650 187.175 ;
        RECT 178.745 187.155 179.015 187.365 ;
        RECT 179.235 187.345 179.565 187.805 ;
        RECT 180.075 187.345 180.825 187.635 ;
        RECT 178.745 186.985 180.080 187.155 ;
        RECT 175.060 185.425 175.340 186.860 ;
        RECT 175.570 186.415 175.855 186.985 ;
        RECT 179.910 186.815 180.080 186.985 ;
        RECT 176.040 186.585 176.510 186.815 ;
        RECT 176.680 186.795 177.010 186.815 ;
        RECT 176.680 186.615 177.130 186.795 ;
        RECT 177.320 186.615 177.650 186.815 ;
        RECT 175.570 186.200 176.720 186.415 ;
        RECT 175.510 185.255 176.220 186.030 ;
        RECT 176.390 185.425 176.720 186.200 ;
        RECT 176.915 185.500 177.130 186.615 ;
        RECT 177.420 186.275 177.650 186.615 ;
        RECT 178.745 186.575 179.095 186.815 ;
        RECT 179.265 186.575 179.740 186.815 ;
        RECT 179.910 186.565 180.285 186.815 ;
        RECT 179.910 186.395 180.080 186.565 ;
        RECT 178.745 186.225 180.080 186.395 ;
        RECT 178.745 186.065 179.025 186.225 ;
        RECT 180.455 186.055 180.825 187.345 ;
        RECT 181.130 187.255 181.300 187.635 ;
        RECT 181.480 187.425 181.810 187.805 ;
        RECT 181.130 187.085 181.795 187.255 ;
        RECT 181.990 187.130 182.250 187.635 ;
        RECT 181.060 186.535 181.390 186.905 ;
        RECT 181.625 186.830 181.795 187.085 ;
        RECT 181.625 186.500 181.910 186.830 ;
        RECT 181.625 186.355 181.795 186.500 ;
        RECT 177.310 185.255 177.640 185.975 ;
        RECT 179.235 185.255 179.485 186.055 ;
        RECT 179.655 185.885 180.825 186.055 ;
        RECT 181.130 186.185 181.795 186.355 ;
        RECT 182.080 186.330 182.250 187.130 ;
        RECT 182.510 187.255 182.680 187.635 ;
        RECT 182.860 187.425 183.190 187.805 ;
        RECT 182.510 187.085 183.175 187.255 ;
        RECT 183.370 187.130 183.630 187.635 ;
        RECT 182.440 186.535 182.770 186.905 ;
        RECT 183.005 186.830 183.175 187.085 ;
        RECT 183.005 186.500 183.290 186.830 ;
        RECT 183.005 186.355 183.175 186.500 ;
        RECT 179.655 185.425 179.985 185.885 ;
        RECT 180.155 185.255 180.370 185.715 ;
        RECT 181.130 185.425 181.300 186.185 ;
        RECT 181.480 185.255 181.810 186.015 ;
        RECT 181.980 185.425 182.250 186.330 ;
        RECT 182.510 186.185 183.175 186.355 ;
        RECT 183.460 186.330 183.630 187.130 ;
        RECT 183.890 187.255 184.060 187.635 ;
        RECT 184.275 187.425 184.605 187.805 ;
        RECT 183.890 187.085 184.605 187.255 ;
        RECT 183.800 186.535 184.155 186.905 ;
        RECT 184.435 186.895 184.605 187.085 ;
        RECT 184.775 187.060 185.030 187.635 ;
        RECT 184.435 186.565 184.690 186.895 ;
        RECT 184.435 186.355 184.605 186.565 ;
        RECT 182.510 185.425 182.680 186.185 ;
        RECT 182.860 185.255 183.190 186.015 ;
        RECT 183.360 185.425 183.630 186.330 ;
        RECT 183.890 186.185 184.605 186.355 ;
        RECT 184.860 186.330 185.030 187.060 ;
        RECT 185.205 186.965 185.465 187.805 ;
        RECT 186.650 187.255 186.820 187.635 ;
        RECT 187.000 187.425 187.330 187.805 ;
        RECT 186.650 187.085 187.315 187.255 ;
        RECT 187.510 187.130 187.770 187.635 ;
        RECT 186.580 186.535 186.910 186.905 ;
        RECT 187.145 186.830 187.315 187.085 ;
        RECT 187.145 186.500 187.430 186.830 ;
        RECT 183.890 185.425 184.060 186.185 ;
        RECT 184.275 185.255 184.605 186.015 ;
        RECT 184.775 185.425 185.030 186.330 ;
        RECT 185.205 185.255 185.465 186.405 ;
        RECT 187.145 186.355 187.315 186.500 ;
        RECT 186.650 186.185 187.315 186.355 ;
        RECT 187.600 186.330 187.770 187.130 ;
        RECT 187.940 187.080 188.230 187.805 ;
        RECT 188.950 187.255 189.120 187.635 ;
        RECT 189.300 187.425 189.630 187.805 ;
        RECT 188.950 187.085 189.615 187.255 ;
        RECT 189.810 187.130 190.070 187.635 ;
        RECT 188.880 186.535 189.210 186.905 ;
        RECT 189.445 186.830 189.615 187.085 ;
        RECT 189.445 186.500 189.730 186.830 ;
        RECT 186.650 185.425 186.820 186.185 ;
        RECT 187.000 185.255 187.330 186.015 ;
        RECT 187.500 185.425 187.770 186.330 ;
        RECT 187.940 185.255 188.230 186.420 ;
        RECT 189.445 186.355 189.615 186.500 ;
        RECT 188.950 186.185 189.615 186.355 ;
        RECT 189.900 186.330 190.070 187.130 ;
        RECT 190.330 187.155 190.500 187.635 ;
        RECT 190.670 187.325 191.000 187.805 ;
        RECT 191.225 187.385 192.760 187.635 ;
        RECT 191.225 187.155 191.395 187.385 ;
        RECT 190.330 186.985 191.395 187.155 ;
        RECT 191.575 186.815 191.855 187.215 ;
        RECT 190.245 186.605 190.595 186.815 ;
        RECT 190.765 186.615 191.210 186.815 ;
        RECT 191.380 186.615 191.855 186.815 ;
        RECT 192.125 186.815 192.410 187.215 ;
        RECT 192.590 187.155 192.760 187.385 ;
        RECT 192.930 187.325 193.260 187.805 ;
        RECT 193.475 187.305 193.730 187.635 ;
        RECT 193.545 187.225 193.730 187.305 ;
        RECT 192.590 186.985 193.390 187.155 ;
        RECT 192.125 186.615 192.455 186.815 ;
        RECT 192.625 186.615 192.990 186.815 ;
        RECT 193.220 186.435 193.390 186.985 ;
        RECT 188.950 185.425 189.120 186.185 ;
        RECT 189.300 185.255 189.630 186.015 ;
        RECT 189.800 185.425 190.070 186.330 ;
        RECT 190.330 186.265 193.390 186.435 ;
        RECT 190.330 185.425 190.500 186.265 ;
        RECT 193.560 186.095 193.730 187.225 ;
        RECT 190.670 185.595 191.000 186.095 ;
        RECT 191.170 185.855 192.805 186.095 ;
        RECT 191.170 185.765 191.400 185.855 ;
        RECT 191.510 185.595 191.840 185.635 ;
        RECT 190.670 185.425 191.840 185.595 ;
        RECT 192.030 185.255 192.385 185.675 ;
        RECT 192.555 185.425 192.805 185.855 ;
        RECT 192.975 185.255 193.305 186.015 ;
        RECT 193.475 185.425 193.730 186.095 ;
        RECT 193.920 187.130 194.180 187.635 ;
        RECT 194.360 187.425 194.690 187.805 ;
        RECT 194.870 187.255 195.040 187.635 ;
        RECT 193.920 186.330 194.090 187.130 ;
        RECT 194.375 187.085 195.040 187.255 ;
        RECT 195.390 187.155 195.560 187.635 ;
        RECT 195.730 187.325 196.060 187.805 ;
        RECT 196.285 187.385 197.820 187.635 ;
        RECT 196.285 187.155 196.455 187.385 ;
        RECT 194.375 186.830 194.545 187.085 ;
        RECT 195.390 186.985 196.455 187.155 ;
        RECT 194.260 186.500 194.545 186.830 ;
        RECT 194.780 186.535 195.110 186.905 ;
        RECT 196.635 186.815 196.915 187.215 ;
        RECT 195.305 186.605 195.655 186.815 ;
        RECT 195.825 186.615 196.270 186.815 ;
        RECT 196.440 186.615 196.915 186.815 ;
        RECT 197.185 186.815 197.470 187.215 ;
        RECT 197.650 187.155 197.820 187.385 ;
        RECT 197.990 187.325 198.320 187.805 ;
        RECT 198.535 187.305 198.790 187.635 ;
        RECT 198.580 187.295 198.790 187.305 ;
        RECT 198.605 187.225 198.790 187.295 ;
        RECT 197.650 186.985 198.450 187.155 ;
        RECT 197.185 186.615 197.515 186.815 ;
        RECT 197.685 186.615 198.050 186.815 ;
        RECT 194.375 186.355 194.545 186.500 ;
        RECT 198.280 186.435 198.450 186.985 ;
        RECT 193.920 185.425 194.190 186.330 ;
        RECT 194.375 186.185 195.040 186.355 ;
        RECT 194.360 185.255 194.690 186.015 ;
        RECT 194.870 185.425 195.040 186.185 ;
        RECT 195.390 186.265 198.450 186.435 ;
        RECT 195.390 185.425 195.560 186.265 ;
        RECT 198.620 186.095 198.790 187.225 ;
        RECT 195.730 185.595 196.060 186.095 ;
        RECT 196.230 185.855 197.865 186.095 ;
        RECT 196.230 185.765 196.460 185.855 ;
        RECT 196.570 185.595 196.900 185.635 ;
        RECT 195.730 185.425 196.900 185.595 ;
        RECT 197.090 185.255 197.445 185.675 ;
        RECT 197.615 185.425 197.865 185.855 ;
        RECT 198.035 185.255 198.365 186.015 ;
        RECT 198.535 185.425 198.790 186.095 ;
        RECT 198.980 187.130 199.240 187.635 ;
        RECT 199.420 187.425 199.750 187.805 ;
        RECT 199.930 187.255 200.100 187.635 ;
        RECT 200.360 187.260 205.705 187.805 ;
        RECT 198.980 186.330 199.150 187.130 ;
        RECT 199.435 187.085 200.100 187.255 ;
        RECT 199.435 186.830 199.605 187.085 ;
        RECT 199.320 186.500 199.605 186.830 ;
        RECT 199.840 186.535 200.170 186.905 ;
        RECT 199.435 186.355 199.605 186.500 ;
        RECT 201.945 186.430 202.285 187.260 ;
        RECT 205.880 187.055 207.090 187.805 ;
        RECT 207.260 187.130 207.520 187.635 ;
        RECT 207.700 187.425 208.030 187.805 ;
        RECT 208.210 187.255 208.380 187.635 ;
        RECT 198.980 185.425 199.250 186.330 ;
        RECT 199.435 186.185 200.100 186.355 ;
        RECT 199.420 185.255 199.750 186.015 ;
        RECT 199.930 185.425 200.100 186.185 ;
        RECT 203.765 185.690 204.115 186.940 ;
        RECT 205.880 186.515 206.400 187.055 ;
        RECT 206.570 186.345 207.090 186.885 ;
        RECT 200.360 185.255 205.705 185.690 ;
        RECT 205.880 185.255 207.090 186.345 ;
        RECT 207.260 186.330 207.430 187.130 ;
        RECT 207.715 187.085 208.380 187.255 ;
        RECT 208.640 187.130 208.900 187.635 ;
        RECT 209.080 187.425 209.410 187.805 ;
        RECT 209.590 187.255 209.760 187.635 ;
        RECT 207.715 186.830 207.885 187.085 ;
        RECT 207.600 186.500 207.885 186.830 ;
        RECT 208.120 186.535 208.450 186.905 ;
        RECT 207.715 186.355 207.885 186.500 ;
        RECT 207.260 185.425 207.530 186.330 ;
        RECT 207.715 186.185 208.380 186.355 ;
        RECT 207.700 185.255 208.030 186.015 ;
        RECT 208.210 185.425 208.380 186.185 ;
        RECT 208.640 186.330 208.810 187.130 ;
        RECT 209.095 187.085 209.760 187.255 ;
        RECT 210.110 187.255 210.280 187.635 ;
        RECT 210.460 187.425 210.790 187.805 ;
        RECT 210.110 187.085 210.775 187.255 ;
        RECT 210.970 187.130 211.230 187.635 ;
        RECT 209.095 186.830 209.265 187.085 ;
        RECT 208.980 186.500 209.265 186.830 ;
        RECT 209.500 186.535 209.830 186.905 ;
        RECT 210.040 186.535 210.370 186.905 ;
        RECT 210.605 186.830 210.775 187.085 ;
        RECT 209.095 186.355 209.265 186.500 ;
        RECT 210.605 186.500 210.890 186.830 ;
        RECT 210.605 186.355 210.775 186.500 ;
        RECT 208.640 185.425 208.910 186.330 ;
        RECT 209.095 186.185 209.760 186.355 ;
        RECT 209.080 185.255 209.410 186.015 ;
        RECT 209.590 185.425 209.760 186.185 ;
        RECT 210.110 186.185 210.775 186.355 ;
        RECT 211.060 186.330 211.230 187.130 ;
        RECT 211.490 187.255 211.660 187.635 ;
        RECT 211.840 187.425 212.170 187.805 ;
        RECT 211.490 187.085 212.155 187.255 ;
        RECT 212.350 187.130 212.610 187.635 ;
        RECT 211.420 186.535 211.750 186.905 ;
        RECT 211.985 186.830 212.155 187.085 ;
        RECT 211.985 186.500 212.270 186.830 ;
        RECT 211.985 186.355 212.155 186.500 ;
        RECT 210.110 185.425 210.280 186.185 ;
        RECT 210.460 185.255 210.790 186.015 ;
        RECT 210.960 185.425 211.230 186.330 ;
        RECT 211.490 186.185 212.155 186.355 ;
        RECT 212.440 186.330 212.610 187.130 ;
        RECT 213.700 187.080 213.990 187.805 ;
        RECT 214.250 187.255 214.420 187.635 ;
        RECT 214.600 187.425 214.930 187.805 ;
        RECT 214.250 187.085 214.915 187.255 ;
        RECT 215.110 187.130 215.370 187.635 ;
        RECT 214.180 186.535 214.510 186.905 ;
        RECT 214.745 186.830 214.915 187.085 ;
        RECT 214.745 186.500 215.030 186.830 ;
        RECT 211.490 185.425 211.660 186.185 ;
        RECT 211.840 185.255 212.170 186.015 ;
        RECT 212.340 185.425 212.610 186.330 ;
        RECT 213.700 185.255 213.990 186.420 ;
        RECT 214.745 186.355 214.915 186.500 ;
        RECT 214.250 186.185 214.915 186.355 ;
        RECT 215.200 186.330 215.370 187.130 ;
        RECT 215.630 187.255 215.800 187.635 ;
        RECT 215.980 187.425 216.310 187.805 ;
        RECT 215.630 187.085 216.295 187.255 ;
        RECT 216.490 187.130 216.750 187.635 ;
        RECT 215.560 186.535 215.890 186.905 ;
        RECT 216.125 186.830 216.295 187.085 ;
        RECT 216.125 186.500 216.410 186.830 ;
        RECT 216.125 186.355 216.295 186.500 ;
        RECT 214.250 185.425 214.420 186.185 ;
        RECT 214.600 185.255 214.930 186.015 ;
        RECT 215.100 185.425 215.370 186.330 ;
        RECT 215.630 186.185 216.295 186.355 ;
        RECT 216.580 186.330 216.750 187.130 ;
        RECT 215.630 185.425 215.800 186.185 ;
        RECT 215.980 185.255 216.310 186.015 ;
        RECT 216.480 185.425 216.750 186.330 ;
        RECT 216.920 187.130 217.180 187.635 ;
        RECT 217.360 187.425 217.690 187.805 ;
        RECT 217.870 187.255 218.040 187.635 ;
        RECT 216.920 186.330 217.090 187.130 ;
        RECT 217.375 187.085 218.040 187.255 ;
        RECT 218.300 187.130 218.560 187.635 ;
        RECT 218.740 187.425 219.070 187.805 ;
        RECT 219.250 187.255 219.420 187.635 ;
        RECT 217.375 186.830 217.545 187.085 ;
        RECT 217.260 186.500 217.545 186.830 ;
        RECT 217.780 186.535 218.110 186.905 ;
        RECT 217.375 186.355 217.545 186.500 ;
        RECT 216.920 185.425 217.190 186.330 ;
        RECT 217.375 186.185 218.040 186.355 ;
        RECT 217.360 185.255 217.690 186.015 ;
        RECT 217.870 185.425 218.040 186.185 ;
        RECT 218.300 186.330 218.470 187.130 ;
        RECT 218.755 187.085 219.420 187.255 ;
        RECT 220.230 187.255 220.400 187.630 ;
        RECT 220.570 187.425 220.900 187.805 ;
        RECT 221.070 187.465 222.145 187.635 ;
        RECT 221.070 187.255 221.240 187.465 ;
        RECT 220.230 187.085 221.240 187.255 ;
        RECT 221.465 187.125 221.805 187.295 ;
        RECT 221.975 187.130 222.145 187.465 ;
        RECT 218.755 186.830 218.925 187.085 ;
        RECT 221.465 186.955 221.755 187.125 ;
        RECT 218.640 186.500 218.925 186.830 ;
        RECT 219.160 186.535 219.490 186.905 ;
        RECT 218.755 186.355 218.925 186.500 ;
        RECT 220.205 186.445 220.550 186.895 ;
        RECT 218.300 185.425 218.570 186.330 ;
        RECT 218.755 186.185 219.420 186.355 ;
        RECT 220.200 186.275 220.550 186.445 ;
        RECT 220.860 186.275 221.295 186.895 ;
        RECT 221.465 186.435 221.635 186.955 ;
        RECT 222.315 186.785 222.675 187.460 ;
        RECT 222.855 187.085 223.145 187.805 ;
        RECT 223.435 187.465 225.035 187.635 ;
        RECT 223.435 187.095 223.605 187.465 ;
        RECT 224.680 187.425 225.035 187.465 ;
        RECT 225.205 187.345 225.375 187.805 ;
        RECT 223.775 187.045 224.105 187.295 ;
        RECT 223.790 186.970 224.105 187.045 ;
        RECT 224.275 187.175 224.445 187.295 ;
        RECT 225.550 187.175 225.795 187.595 ;
        RECT 226.065 187.425 226.395 187.805 ;
        RECT 226.565 187.235 226.740 187.565 ;
        RECT 227.085 187.475 227.255 187.635 ;
        RECT 227.085 187.305 227.615 187.475 ;
        RECT 227.785 187.465 228.780 187.635 ;
        RECT 227.785 187.305 227.955 187.465 ;
        RECT 224.275 187.005 225.795 187.175 ;
        RECT 222.135 186.605 222.675 186.785 ;
        RECT 222.315 186.495 222.675 186.605 ;
        RECT 221.465 186.265 222.100 186.435 ;
        RECT 222.315 186.265 223.120 186.495 ;
        RECT 218.740 185.255 219.070 186.015 ;
        RECT 219.250 185.425 219.420 186.185 ;
        RECT 220.230 185.925 221.760 186.095 ;
        RECT 220.230 185.425 220.400 185.925 ;
        RECT 221.590 185.765 221.760 185.925 ;
        RECT 221.930 185.935 222.100 186.265 ;
        RECT 221.930 185.765 222.260 185.935 ;
        RECT 220.570 185.255 220.900 185.635 ;
        RECT 221.070 185.595 221.240 185.755 ;
        RECT 222.430 185.595 222.600 186.095 ;
        RECT 221.070 185.425 222.600 185.595 ;
        RECT 222.770 185.425 223.120 186.265 ;
        RECT 223.320 185.895 223.620 186.895 ;
        RECT 223.790 186.445 223.960 186.970 ;
        RECT 224.275 186.965 224.445 187.005 ;
        RECT 224.130 186.785 224.460 186.795 ;
        RECT 224.130 186.625 224.515 186.785 ;
        RECT 224.345 186.615 224.515 186.625 ;
        RECT 224.855 186.445 225.100 186.835 ;
        RECT 223.790 186.275 224.550 186.445 ;
        RECT 224.800 186.275 225.100 186.445 ;
        RECT 223.290 185.255 223.620 185.635 ;
        RECT 223.880 185.595 224.050 186.105 ;
        RECT 224.220 185.765 224.550 186.275 ;
        RECT 224.855 186.215 225.100 186.275 ;
        RECT 225.305 186.445 225.635 186.835 ;
        RECT 225.305 186.275 225.660 186.445 ;
        RECT 225.305 186.215 225.635 186.275 ;
        RECT 226.110 186.215 226.400 186.895 ;
        RECT 226.570 186.785 226.740 187.235 ;
        RECT 227.035 186.955 227.275 187.125 ;
        RECT 226.570 186.615 226.860 186.785 ;
        RECT 224.720 185.805 225.785 185.975 ;
        RECT 224.720 185.595 224.890 185.805 ;
        RECT 223.880 185.425 224.890 185.595 ;
        RECT 225.115 185.255 225.445 185.635 ;
        RECT 225.615 185.425 225.785 185.805 ;
        RECT 226.570 185.755 226.740 186.615 ;
        RECT 226.035 185.255 226.385 185.635 ;
        RECT 226.555 185.425 226.740 185.755 ;
        RECT 227.035 185.755 227.205 186.955 ;
        RECT 227.445 186.135 227.615 187.305 ;
        RECT 228.265 187.125 228.440 187.295 ;
        RECT 228.025 186.965 228.440 187.125 ;
        RECT 228.610 187.175 228.780 187.465 ;
        RECT 228.950 187.345 229.120 187.805 ;
        RECT 228.610 187.005 229.180 187.175 ;
        RECT 228.025 186.955 228.435 186.965 ;
        RECT 228.245 186.615 228.700 186.785 ;
        RECT 229.010 186.225 229.180 187.005 ;
        RECT 227.445 185.905 228.230 186.135 ;
        RECT 227.900 185.765 228.230 185.905 ;
        RECT 228.530 186.055 229.180 186.225 ;
        RECT 227.035 185.425 227.245 185.755 ;
        RECT 227.415 185.595 227.745 185.635 ;
        RECT 228.530 185.595 228.700 186.055 ;
        RECT 227.415 185.425 228.700 185.595 ;
        RECT 228.870 185.255 229.200 185.635 ;
        RECT 229.370 185.425 229.630 187.635 ;
        RECT 229.800 187.175 230.140 187.635 ;
        RECT 230.310 187.345 230.480 187.805 ;
        RECT 231.110 187.370 231.470 187.635 ;
        RECT 231.115 187.365 231.470 187.370 ;
        RECT 231.120 187.355 231.470 187.365 ;
        RECT 231.125 187.350 231.470 187.355 ;
        RECT 231.130 187.340 231.470 187.350 ;
        RECT 231.710 187.345 231.880 187.805 ;
        RECT 231.135 187.335 231.470 187.340 ;
        RECT 231.145 187.325 231.470 187.335 ;
        RECT 231.155 187.315 231.470 187.325 ;
        RECT 230.650 187.175 230.980 187.255 ;
        RECT 229.800 186.985 230.980 187.175 ;
        RECT 231.170 187.175 231.470 187.315 ;
        RECT 231.170 186.985 231.880 187.175 ;
        RECT 229.800 186.615 230.130 186.815 ;
        RECT 230.440 186.795 230.770 186.815 ;
        RECT 230.320 186.615 230.770 186.795 ;
        RECT 229.800 186.275 230.030 186.615 ;
        RECT 229.810 185.255 230.140 185.975 ;
        RECT 230.320 185.500 230.535 186.615 ;
        RECT 230.940 186.585 231.410 186.815 ;
        RECT 231.595 186.415 231.880 186.985 ;
        RECT 232.050 186.860 232.390 187.635 ;
        RECT 230.730 186.200 231.880 186.415 ;
        RECT 230.730 185.425 231.060 186.200 ;
        RECT 231.230 185.255 231.940 186.030 ;
        RECT 232.110 185.425 232.390 186.860 ;
        RECT 232.560 187.130 232.820 187.635 ;
        RECT 233.000 187.425 233.330 187.805 ;
        RECT 233.510 187.255 233.680 187.635 ;
        RECT 232.560 186.330 232.730 187.130 ;
        RECT 233.015 187.085 233.680 187.255 ;
        RECT 233.015 186.830 233.185 187.085 ;
        RECT 234.860 187.055 236.070 187.805 ;
        RECT 232.900 186.500 233.185 186.830 ;
        RECT 233.420 186.535 233.750 186.905 ;
        RECT 233.015 186.355 233.185 186.500 ;
        RECT 232.560 185.425 232.830 186.330 ;
        RECT 233.015 186.185 233.680 186.355 ;
        RECT 233.000 185.255 233.330 186.015 ;
        RECT 233.510 185.425 233.680 186.185 ;
        RECT 234.860 186.345 235.380 186.885 ;
        RECT 235.550 186.515 236.070 187.055 ;
        RECT 234.860 185.255 236.070 186.345 ;
        RECT 162.095 185.085 236.155 185.255 ;
        RECT 108.630 184.880 153.130 185.050 ;
        RECT 162.180 183.995 163.390 185.085 ;
        RECT 162.180 183.285 162.700 183.825 ;
        RECT 162.870 183.455 163.390 183.995 ;
        RECT 164.110 184.155 164.280 184.915 ;
        RECT 164.460 184.325 164.790 185.085 ;
        RECT 164.110 183.985 164.775 184.155 ;
        RECT 164.960 184.010 165.230 184.915 ;
        RECT 164.605 183.840 164.775 183.985 ;
        RECT 164.040 183.435 164.370 183.805 ;
        RECT 164.605 183.510 164.890 183.840 ;
        RECT 162.180 182.535 163.390 183.285 ;
        RECT 164.605 183.255 164.775 183.510 ;
        RECT 164.110 183.085 164.775 183.255 ;
        RECT 165.060 183.210 165.230 184.010 ;
        RECT 165.490 184.155 165.660 184.915 ;
        RECT 165.840 184.325 166.170 185.085 ;
        RECT 165.490 183.985 166.155 184.155 ;
        RECT 166.340 184.010 166.610 184.915 ;
        RECT 165.985 183.840 166.155 183.985 ;
        RECT 165.420 183.435 165.750 183.805 ;
        RECT 165.985 183.510 166.270 183.840 ;
        RECT 165.985 183.255 166.155 183.510 ;
        RECT 164.110 182.705 164.280 183.085 ;
        RECT 164.460 182.535 164.790 182.915 ;
        RECT 164.970 182.705 165.230 183.210 ;
        RECT 165.490 183.085 166.155 183.255 ;
        RECT 166.440 183.210 166.610 184.010 ;
        RECT 165.490 182.705 165.660 183.085 ;
        RECT 165.840 182.535 166.170 182.915 ;
        RECT 166.350 182.705 166.610 183.210 ;
        RECT 166.800 184.245 167.055 184.915 ;
        RECT 167.225 184.325 167.555 185.085 ;
        RECT 167.725 184.485 167.975 184.915 ;
        RECT 168.145 184.665 168.500 185.085 ;
        RECT 168.690 184.745 169.860 184.915 ;
        RECT 168.690 184.705 169.020 184.745 ;
        RECT 169.130 184.485 169.360 184.575 ;
        RECT 167.725 184.245 169.360 184.485 ;
        RECT 169.530 184.245 169.860 184.745 ;
        RECT 166.800 183.115 166.970 184.245 ;
        RECT 170.030 184.075 170.200 184.915 ;
        RECT 167.140 183.905 170.200 184.075 ;
        RECT 171.470 184.075 171.640 184.915 ;
        RECT 171.810 184.745 172.980 184.915 ;
        RECT 171.810 184.245 172.140 184.745 ;
        RECT 172.650 184.705 172.980 184.745 ;
        RECT 173.170 184.665 173.525 185.085 ;
        RECT 172.310 184.485 172.540 184.575 ;
        RECT 173.695 184.485 173.945 184.915 ;
        RECT 172.310 184.245 173.945 184.485 ;
        RECT 174.115 184.325 174.445 185.085 ;
        RECT 174.615 184.245 174.870 184.915 ;
        RECT 171.470 183.905 174.530 184.075 ;
        RECT 167.140 183.355 167.310 183.905 ;
        RECT 167.540 183.525 167.905 183.725 ;
        RECT 168.075 183.525 168.405 183.725 ;
        RECT 167.140 183.185 167.940 183.355 ;
        RECT 166.800 183.035 166.985 183.115 ;
        RECT 166.800 182.705 167.055 183.035 ;
        RECT 167.270 182.535 167.600 183.015 ;
        RECT 167.770 182.955 167.940 183.185 ;
        RECT 168.120 183.125 168.405 183.525 ;
        RECT 168.675 183.525 169.150 183.725 ;
        RECT 169.320 183.525 169.765 183.725 ;
        RECT 169.935 183.525 170.285 183.735 ;
        RECT 171.385 183.525 171.735 183.735 ;
        RECT 171.905 183.525 172.350 183.725 ;
        RECT 172.520 183.525 172.995 183.725 ;
        RECT 168.675 183.125 168.955 183.525 ;
        RECT 169.135 183.185 170.200 183.355 ;
        RECT 169.135 182.955 169.305 183.185 ;
        RECT 167.770 182.705 169.305 182.955 ;
        RECT 169.530 182.535 169.860 183.015 ;
        RECT 170.030 182.705 170.200 183.185 ;
        RECT 171.470 183.185 172.535 183.355 ;
        RECT 171.470 182.705 171.640 183.185 ;
        RECT 171.810 182.535 172.140 183.015 ;
        RECT 172.365 182.955 172.535 183.185 ;
        RECT 172.715 183.125 172.995 183.525 ;
        RECT 173.265 183.525 173.595 183.725 ;
        RECT 173.765 183.525 174.130 183.725 ;
        RECT 173.265 183.125 173.550 183.525 ;
        RECT 174.360 183.355 174.530 183.905 ;
        RECT 173.730 183.185 174.530 183.355 ;
        RECT 173.730 182.955 173.900 183.185 ;
        RECT 174.700 183.115 174.870 184.245 ;
        RECT 175.060 183.920 175.350 185.085 ;
        RECT 175.735 183.985 176.065 185.085 ;
        RECT 176.540 184.485 176.865 184.915 ;
        RECT 177.035 184.665 177.365 185.085 ;
        RECT 178.110 184.655 178.520 185.085 ;
        RECT 176.540 184.315 178.520 184.485 ;
        RECT 176.540 183.905 177.245 184.315 ;
        RECT 175.520 183.525 176.165 183.735 ;
        RECT 176.335 183.525 176.905 183.735 ;
        RECT 174.685 183.035 174.870 183.115 ;
        RECT 172.365 182.705 173.900 182.955 ;
        RECT 174.070 182.535 174.400 183.015 ;
        RECT 174.615 182.705 174.870 183.035 ;
        RECT 175.060 182.535 175.350 183.260 ;
        RECT 175.675 183.185 176.845 183.355 ;
        RECT 175.675 182.720 176.005 183.185 ;
        RECT 176.175 182.535 176.345 183.005 ;
        RECT 176.515 182.705 176.845 183.185 ;
        RECT 177.075 182.705 177.245 183.905 ;
        RECT 177.415 183.975 178.040 184.145 ;
        RECT 177.415 183.275 177.585 183.975 ;
        RECT 178.255 183.775 178.520 184.315 ;
        RECT 178.690 183.930 179.030 184.915 ;
        RECT 179.750 184.155 179.920 184.915 ;
        RECT 180.100 184.325 180.430 185.085 ;
        RECT 179.750 183.985 180.415 184.155 ;
        RECT 180.600 184.010 180.870 184.915 ;
        RECT 177.755 183.445 178.085 183.775 ;
        RECT 178.255 183.445 178.605 183.775 ;
        RECT 178.775 183.275 179.030 183.930 ;
        RECT 180.245 183.840 180.415 183.985 ;
        RECT 179.680 183.435 180.010 183.805 ;
        RECT 180.245 183.510 180.530 183.840 ;
        RECT 177.415 183.105 177.955 183.275 ;
        RECT 177.785 182.900 177.955 183.105 ;
        RECT 178.235 182.535 178.405 183.275 ;
        RECT 178.670 182.900 179.030 183.275 ;
        RECT 180.245 183.255 180.415 183.510 ;
        RECT 179.750 183.085 180.415 183.255 ;
        RECT 180.700 183.210 180.870 184.010 ;
        RECT 179.750 182.705 179.920 183.085 ;
        RECT 180.100 182.535 180.430 182.915 ;
        RECT 180.610 182.705 180.870 183.210 ;
        RECT 181.040 184.010 181.310 184.915 ;
        RECT 181.480 184.325 181.810 185.085 ;
        RECT 181.990 184.155 182.160 184.915 ;
        RECT 181.040 183.210 181.210 184.010 ;
        RECT 181.495 183.985 182.160 184.155 ;
        RECT 182.510 184.155 182.680 184.915 ;
        RECT 182.860 184.325 183.190 185.085 ;
        RECT 182.510 183.985 183.175 184.155 ;
        RECT 183.360 184.010 183.630 184.915 ;
        RECT 181.495 183.840 181.665 183.985 ;
        RECT 181.380 183.510 181.665 183.840 ;
        RECT 183.005 183.840 183.175 183.985 ;
        RECT 181.495 183.255 181.665 183.510 ;
        RECT 181.900 183.435 182.230 183.805 ;
        RECT 182.440 183.435 182.770 183.805 ;
        RECT 183.005 183.510 183.290 183.840 ;
        RECT 183.005 183.255 183.175 183.510 ;
        RECT 181.040 182.705 181.300 183.210 ;
        RECT 181.495 183.085 182.160 183.255 ;
        RECT 181.480 182.535 181.810 182.915 ;
        RECT 181.990 182.705 182.160 183.085 ;
        RECT 182.510 183.085 183.175 183.255 ;
        RECT 183.460 183.210 183.630 184.010 ;
        RECT 183.890 184.155 184.060 184.915 ;
        RECT 184.240 184.325 184.570 185.085 ;
        RECT 183.890 183.985 184.555 184.155 ;
        RECT 184.740 184.010 185.010 184.915 ;
        RECT 184.385 183.840 184.555 183.985 ;
        RECT 183.820 183.435 184.150 183.805 ;
        RECT 184.385 183.510 184.670 183.840 ;
        RECT 184.385 183.255 184.555 183.510 ;
        RECT 182.510 182.705 182.680 183.085 ;
        RECT 182.860 182.535 183.190 182.915 ;
        RECT 183.370 182.705 183.630 183.210 ;
        RECT 183.890 183.085 184.555 183.255 ;
        RECT 184.840 183.210 185.010 184.010 ;
        RECT 185.270 184.155 185.440 184.915 ;
        RECT 185.620 184.325 185.950 185.085 ;
        RECT 185.270 183.985 185.935 184.155 ;
        RECT 186.120 184.010 186.390 184.915 ;
        RECT 187.055 184.285 187.305 185.085 ;
        RECT 187.475 184.455 187.805 184.915 ;
        RECT 187.975 184.625 188.190 185.085 ;
        RECT 187.475 184.285 188.645 184.455 ;
        RECT 185.765 183.840 185.935 183.985 ;
        RECT 185.200 183.435 185.530 183.805 ;
        RECT 185.765 183.510 186.050 183.840 ;
        RECT 185.765 183.255 185.935 183.510 ;
        RECT 183.890 182.705 184.060 183.085 ;
        RECT 184.240 182.535 184.570 182.915 ;
        RECT 184.750 182.705 185.010 183.210 ;
        RECT 185.270 183.085 185.935 183.255 ;
        RECT 186.220 183.210 186.390 184.010 ;
        RECT 186.565 184.115 186.845 184.275 ;
        RECT 186.565 183.945 187.900 184.115 ;
        RECT 187.730 183.775 187.900 183.945 ;
        RECT 186.565 183.525 186.915 183.765 ;
        RECT 187.085 183.525 187.560 183.765 ;
        RECT 187.730 183.525 188.105 183.775 ;
        RECT 187.730 183.355 187.900 183.525 ;
        RECT 185.270 182.705 185.440 183.085 ;
        RECT 185.620 182.535 185.950 182.915 ;
        RECT 186.130 182.705 186.390 183.210 ;
        RECT 186.565 183.185 187.900 183.355 ;
        RECT 186.565 182.975 186.835 183.185 ;
        RECT 188.275 182.995 188.645 184.285 ;
        RECT 188.950 184.075 189.120 184.915 ;
        RECT 189.290 184.745 190.460 184.915 ;
        RECT 189.290 184.245 189.620 184.745 ;
        RECT 190.130 184.705 190.460 184.745 ;
        RECT 190.650 184.665 191.005 185.085 ;
        RECT 189.790 184.485 190.020 184.575 ;
        RECT 191.175 184.485 191.425 184.915 ;
        RECT 189.790 184.245 191.425 184.485 ;
        RECT 191.595 184.325 191.925 185.085 ;
        RECT 192.095 184.245 192.350 184.915 ;
        RECT 188.950 183.905 192.010 184.075 ;
        RECT 188.865 183.525 189.215 183.735 ;
        RECT 189.385 183.525 189.830 183.725 ;
        RECT 190.000 183.525 190.475 183.725 ;
        RECT 187.055 182.535 187.385 182.995 ;
        RECT 187.895 182.705 188.645 182.995 ;
        RECT 188.950 183.185 190.015 183.355 ;
        RECT 188.950 182.705 189.120 183.185 ;
        RECT 189.290 182.535 189.620 183.015 ;
        RECT 189.845 182.955 190.015 183.185 ;
        RECT 190.195 183.125 190.475 183.525 ;
        RECT 190.745 183.525 191.075 183.725 ;
        RECT 191.245 183.555 191.620 183.725 ;
        RECT 191.245 183.525 191.610 183.555 ;
        RECT 190.745 183.125 191.030 183.525 ;
        RECT 191.840 183.355 192.010 183.905 ;
        RECT 191.210 183.185 192.010 183.355 ;
        RECT 191.210 182.955 191.380 183.185 ;
        RECT 192.180 183.115 192.350 184.245 ;
        RECT 192.630 184.075 192.800 184.915 ;
        RECT 192.970 184.745 194.140 184.915 ;
        RECT 192.970 184.245 193.300 184.745 ;
        RECT 193.810 184.705 194.140 184.745 ;
        RECT 194.330 184.665 194.685 185.085 ;
        RECT 193.470 184.485 193.700 184.575 ;
        RECT 194.855 184.485 195.105 184.915 ;
        RECT 193.470 184.245 195.105 184.485 ;
        RECT 195.275 184.325 195.605 185.085 ;
        RECT 195.775 184.245 196.030 184.915 ;
        RECT 195.820 184.235 196.030 184.245 ;
        RECT 192.630 183.905 195.690 184.075 ;
        RECT 192.545 183.525 192.895 183.735 ;
        RECT 193.065 183.525 193.510 183.725 ;
        RECT 193.680 183.525 194.155 183.725 ;
        RECT 192.165 183.045 192.350 183.115 ;
        RECT 192.140 183.035 192.350 183.045 ;
        RECT 189.845 182.705 191.380 182.955 ;
        RECT 191.550 182.535 191.880 183.015 ;
        RECT 192.095 182.705 192.350 183.035 ;
        RECT 192.630 183.185 193.695 183.355 ;
        RECT 192.630 182.705 192.800 183.185 ;
        RECT 192.970 182.535 193.300 183.015 ;
        RECT 193.525 182.955 193.695 183.185 ;
        RECT 193.875 183.125 194.155 183.525 ;
        RECT 194.425 183.525 194.755 183.725 ;
        RECT 194.925 183.555 195.300 183.725 ;
        RECT 194.925 183.525 195.290 183.555 ;
        RECT 194.425 183.125 194.710 183.525 ;
        RECT 195.520 183.355 195.690 183.905 ;
        RECT 194.890 183.185 195.690 183.355 ;
        RECT 194.890 182.955 195.060 183.185 ;
        RECT 195.860 183.115 196.030 184.235 ;
        RECT 195.845 183.035 196.030 183.115 ;
        RECT 193.525 182.705 195.060 182.955 ;
        RECT 195.230 182.535 195.560 183.015 ;
        RECT 195.775 182.705 196.030 183.035 ;
        RECT 196.225 183.945 196.560 184.915 ;
        RECT 196.730 183.945 196.900 185.085 ;
        RECT 197.070 184.745 199.100 184.915 ;
        RECT 196.225 183.275 196.395 183.945 ;
        RECT 197.070 183.775 197.240 184.745 ;
        RECT 196.565 183.445 196.820 183.775 ;
        RECT 197.045 183.445 197.240 183.775 ;
        RECT 197.410 184.405 198.535 184.575 ;
        RECT 196.650 183.275 196.820 183.445 ;
        RECT 197.410 183.275 197.580 184.405 ;
        RECT 196.225 182.705 196.480 183.275 ;
        RECT 196.650 183.105 197.580 183.275 ;
        RECT 197.750 184.065 198.760 184.235 ;
        RECT 197.750 183.265 197.920 184.065 ;
        RECT 198.125 183.725 198.400 183.865 ;
        RECT 198.120 183.555 198.400 183.725 ;
        RECT 197.405 183.070 197.580 183.105 ;
        RECT 196.650 182.535 196.980 182.935 ;
        RECT 197.405 182.705 197.935 183.070 ;
        RECT 198.125 182.705 198.400 183.555 ;
        RECT 198.570 182.705 198.760 184.065 ;
        RECT 198.930 184.080 199.100 184.745 ;
        RECT 199.270 184.325 199.440 185.085 ;
        RECT 199.675 184.325 200.190 184.735 ;
        RECT 198.930 183.890 199.680 184.080 ;
        RECT 199.850 183.515 200.190 184.325 ;
        RECT 200.820 183.920 201.110 185.085 ;
        RECT 201.280 184.010 201.550 184.915 ;
        RECT 201.720 184.325 202.050 185.085 ;
        RECT 202.230 184.155 202.400 184.915 ;
        RECT 198.960 183.345 200.190 183.515 ;
        RECT 198.940 182.535 199.450 183.070 ;
        RECT 199.670 182.740 199.915 183.345 ;
        RECT 200.820 182.535 201.110 183.260 ;
        RECT 201.280 183.210 201.450 184.010 ;
        RECT 201.735 183.985 202.400 184.155 ;
        RECT 202.660 184.010 202.930 184.915 ;
        RECT 203.100 184.325 203.430 185.085 ;
        RECT 203.610 184.155 203.780 184.915 ;
        RECT 201.735 183.840 201.905 183.985 ;
        RECT 201.620 183.510 201.905 183.840 ;
        RECT 201.735 183.255 201.905 183.510 ;
        RECT 202.140 183.435 202.470 183.805 ;
        RECT 201.280 182.705 201.540 183.210 ;
        RECT 201.735 183.085 202.400 183.255 ;
        RECT 201.720 182.535 202.050 182.915 ;
        RECT 202.230 182.705 202.400 183.085 ;
        RECT 202.660 183.210 202.830 184.010 ;
        RECT 203.115 183.985 203.780 184.155 ;
        RECT 204.040 183.995 205.250 185.085 ;
        RECT 205.510 184.415 205.680 184.915 ;
        RECT 205.850 184.705 206.180 185.085 ;
        RECT 206.350 184.745 207.880 184.915 ;
        RECT 206.350 184.585 206.520 184.745 ;
        RECT 206.870 184.415 207.040 184.575 ;
        RECT 205.510 184.245 207.040 184.415 ;
        RECT 207.210 184.405 207.540 184.575 ;
        RECT 207.210 184.075 207.380 184.405 ;
        RECT 207.710 184.245 207.880 184.745 ;
        RECT 208.050 184.075 208.400 184.915 ;
        RECT 208.570 184.705 208.900 185.085 ;
        RECT 209.160 184.745 210.170 184.915 ;
        RECT 203.115 183.840 203.285 183.985 ;
        RECT 203.000 183.510 203.285 183.840 ;
        RECT 203.115 183.255 203.285 183.510 ;
        RECT 203.520 183.435 203.850 183.805 ;
        RECT 204.040 183.285 204.560 183.825 ;
        RECT 204.730 183.455 205.250 183.995 ;
        RECT 205.480 183.895 205.830 184.065 ;
        RECT 205.485 183.445 205.830 183.895 ;
        RECT 206.140 183.445 206.575 184.065 ;
        RECT 206.745 183.905 207.380 184.075 ;
        RECT 206.745 183.385 206.915 183.905 ;
        RECT 207.595 183.845 208.400 184.075 ;
        RECT 207.595 183.735 207.955 183.845 ;
        RECT 207.415 183.555 207.955 183.735 ;
        RECT 202.660 182.705 202.920 183.210 ;
        RECT 203.115 183.085 203.780 183.255 ;
        RECT 203.100 182.535 203.430 182.915 ;
        RECT 203.610 182.705 203.780 183.085 ;
        RECT 204.040 182.535 205.250 183.285 ;
        RECT 205.510 183.085 206.520 183.255 ;
        RECT 205.510 182.710 205.680 183.085 ;
        RECT 205.850 182.535 206.180 182.915 ;
        RECT 206.350 182.875 206.520 183.085 ;
        RECT 206.745 183.215 207.035 183.385 ;
        RECT 206.745 183.045 207.085 183.215 ;
        RECT 207.255 182.875 207.425 183.210 ;
        RECT 207.595 182.880 207.955 183.555 ;
        RECT 208.600 183.445 208.900 184.445 ;
        RECT 209.160 184.235 209.330 184.745 ;
        RECT 209.500 184.065 209.830 184.575 ;
        RECT 210.000 184.535 210.170 184.745 ;
        RECT 210.395 184.705 210.725 185.085 ;
        RECT 210.895 184.535 211.065 184.915 ;
        RECT 211.315 184.705 211.665 185.085 ;
        RECT 211.835 184.585 212.020 184.915 ;
        RECT 210.000 184.365 211.065 184.535 ;
        RECT 210.135 184.065 210.380 184.125 ;
        RECT 209.070 183.895 209.830 184.065 ;
        RECT 210.080 183.895 210.380 184.065 ;
        RECT 209.070 183.370 209.240 183.895 ;
        RECT 209.625 183.715 209.795 183.725 ;
        RECT 209.410 183.555 209.795 183.715 ;
        RECT 209.410 183.545 209.740 183.555 ;
        RECT 210.135 183.505 210.380 183.895 ;
        RECT 210.585 183.505 210.915 184.125 ;
        RECT 211.390 183.445 211.680 184.125 ;
        RECT 211.850 183.725 212.020 184.585 ;
        RECT 212.315 184.585 212.525 184.915 ;
        RECT 212.695 184.745 213.980 184.915 ;
        RECT 212.695 184.705 213.025 184.745 ;
        RECT 211.850 183.555 212.140 183.725 ;
        RECT 209.070 183.295 209.385 183.370 ;
        RECT 206.350 182.705 207.425 182.875 ;
        RECT 208.135 182.535 208.425 183.255 ;
        RECT 208.715 182.875 208.885 183.245 ;
        RECT 209.055 183.045 209.385 183.295 ;
        RECT 209.555 183.335 209.725 183.375 ;
        RECT 209.555 183.165 211.075 183.335 ;
        RECT 209.555 183.045 209.725 183.165 ;
        RECT 209.960 182.875 210.315 182.915 ;
        RECT 208.715 182.705 210.315 182.875 ;
        RECT 210.485 182.535 210.655 182.995 ;
        RECT 210.830 182.745 211.075 183.165 ;
        RECT 211.850 183.105 212.020 183.555 ;
        RECT 212.315 183.385 212.485 184.585 ;
        RECT 213.180 184.435 213.510 184.575 ;
        RECT 212.725 184.205 213.510 184.435 ;
        RECT 213.810 184.285 213.980 184.745 ;
        RECT 214.150 184.705 214.480 185.085 ;
        RECT 212.315 183.215 212.555 183.385 ;
        RECT 211.345 182.535 211.675 182.915 ;
        RECT 211.845 182.775 212.020 183.105 ;
        RECT 212.725 183.035 212.895 184.205 ;
        RECT 213.810 184.115 214.460 184.285 ;
        RECT 213.525 183.555 213.980 183.725 ;
        RECT 213.305 183.375 213.715 183.385 ;
        RECT 213.305 183.215 213.720 183.375 ;
        RECT 214.290 183.335 214.460 184.115 ;
        RECT 213.545 183.045 213.720 183.215 ;
        RECT 213.890 183.165 214.460 183.335 ;
        RECT 212.365 182.865 212.895 183.035 ;
        RECT 213.065 182.875 213.235 183.035 ;
        RECT 213.890 182.875 214.060 183.165 ;
        RECT 212.365 182.705 212.535 182.865 ;
        RECT 213.065 182.705 214.060 182.875 ;
        RECT 214.230 182.535 214.400 182.995 ;
        RECT 214.650 182.705 214.910 184.915 ;
        RECT 215.170 184.155 215.340 184.915 ;
        RECT 215.520 184.325 215.850 185.085 ;
        RECT 215.170 183.985 215.835 184.155 ;
        RECT 216.020 184.010 216.290 184.915 ;
        RECT 217.010 184.415 217.180 184.915 ;
        RECT 217.350 184.705 217.680 185.085 ;
        RECT 217.850 184.745 219.380 184.915 ;
        RECT 217.850 184.585 218.020 184.745 ;
        RECT 218.370 184.415 218.540 184.575 ;
        RECT 217.010 184.245 218.540 184.415 ;
        RECT 218.710 184.405 219.040 184.575 ;
        RECT 218.710 184.075 218.880 184.405 ;
        RECT 219.210 184.245 219.380 184.745 ;
        RECT 219.550 184.075 219.900 184.915 ;
        RECT 220.070 184.705 220.400 185.085 ;
        RECT 220.660 184.745 221.670 184.915 ;
        RECT 215.665 183.840 215.835 183.985 ;
        RECT 215.100 183.435 215.430 183.805 ;
        RECT 215.665 183.510 215.950 183.840 ;
        RECT 215.665 183.255 215.835 183.510 ;
        RECT 215.170 183.085 215.835 183.255 ;
        RECT 216.120 183.210 216.290 184.010 ;
        RECT 216.985 183.725 217.330 184.065 ;
        RECT 216.980 183.555 217.330 183.725 ;
        RECT 216.985 183.445 217.330 183.555 ;
        RECT 217.640 183.445 218.075 184.065 ;
        RECT 218.245 183.905 218.880 184.075 ;
        RECT 218.245 183.385 218.415 183.905 ;
        RECT 219.095 183.845 219.900 184.075 ;
        RECT 219.095 183.735 219.455 183.845 ;
        RECT 218.915 183.555 219.455 183.735 ;
        RECT 215.170 182.705 215.340 183.085 ;
        RECT 215.520 182.535 215.850 182.915 ;
        RECT 216.030 182.705 216.290 183.210 ;
        RECT 217.010 183.085 218.020 183.255 ;
        RECT 217.010 182.710 217.180 183.085 ;
        RECT 217.350 182.535 217.680 182.915 ;
        RECT 217.850 182.875 218.020 183.085 ;
        RECT 218.245 183.215 218.535 183.385 ;
        RECT 218.245 183.045 218.585 183.215 ;
        RECT 218.755 182.875 218.925 183.210 ;
        RECT 219.095 182.880 219.455 183.555 ;
        RECT 220.100 183.445 220.400 184.445 ;
        RECT 220.660 184.235 220.830 184.745 ;
        RECT 221.000 184.065 221.330 184.575 ;
        RECT 221.500 184.535 221.670 184.745 ;
        RECT 221.895 184.705 222.225 185.085 ;
        RECT 222.395 184.535 222.565 184.915 ;
        RECT 222.815 184.705 223.165 185.085 ;
        RECT 223.335 184.585 223.520 184.915 ;
        RECT 221.500 184.365 222.565 184.535 ;
        RECT 220.570 183.895 221.330 184.065 ;
        RECT 220.570 183.370 220.740 183.895 ;
        RECT 221.635 183.725 221.880 184.125 ;
        RECT 221.125 183.715 221.295 183.725 ;
        RECT 220.910 183.555 221.295 183.715 ;
        RECT 221.580 183.555 221.880 183.725 ;
        RECT 220.910 183.545 221.240 183.555 ;
        RECT 221.635 183.505 221.880 183.555 ;
        RECT 222.085 183.505 222.415 184.125 ;
        RECT 222.890 183.445 223.180 184.125 ;
        RECT 223.350 183.725 223.520 184.585 ;
        RECT 223.815 184.585 224.025 184.915 ;
        RECT 224.195 184.745 225.480 184.915 ;
        RECT 224.195 184.705 224.525 184.745 ;
        RECT 223.350 183.555 223.640 183.725 ;
        RECT 220.570 183.295 220.885 183.370 ;
        RECT 217.850 182.705 218.925 182.875 ;
        RECT 219.635 182.535 219.925 183.255 ;
        RECT 220.215 182.875 220.385 183.245 ;
        RECT 220.555 183.045 220.885 183.295 ;
        RECT 221.055 183.335 221.225 183.375 ;
        RECT 221.055 183.165 222.575 183.335 ;
        RECT 221.055 183.045 221.225 183.165 ;
        RECT 221.460 182.875 221.815 182.915 ;
        RECT 220.215 182.705 221.815 182.875 ;
        RECT 221.985 182.535 222.155 182.995 ;
        RECT 222.330 182.745 222.575 183.165 ;
        RECT 223.350 183.105 223.520 183.555 ;
        RECT 223.815 183.385 223.985 184.585 ;
        RECT 224.680 184.435 225.010 184.575 ;
        RECT 224.225 184.205 225.010 184.435 ;
        RECT 225.310 184.285 225.480 184.745 ;
        RECT 225.650 184.705 225.980 185.085 ;
        RECT 223.815 183.215 224.055 183.385 ;
        RECT 222.845 182.535 223.175 182.915 ;
        RECT 223.345 182.775 223.520 183.105 ;
        RECT 224.225 183.035 224.395 184.205 ;
        RECT 225.310 184.115 225.960 184.285 ;
        RECT 225.025 183.555 225.480 183.725 ;
        RECT 224.805 183.375 225.215 183.385 ;
        RECT 224.805 183.215 225.220 183.375 ;
        RECT 225.790 183.335 225.960 184.115 ;
        RECT 225.045 183.045 225.220 183.215 ;
        RECT 225.390 183.165 225.960 183.335 ;
        RECT 223.865 182.865 224.395 183.035 ;
        RECT 224.565 182.875 224.735 183.035 ;
        RECT 225.390 182.875 225.560 183.165 ;
        RECT 223.865 182.705 224.035 182.865 ;
        RECT 224.565 182.705 225.560 182.875 ;
        RECT 225.730 182.535 225.900 182.995 ;
        RECT 226.150 182.705 226.410 184.915 ;
        RECT 226.580 183.920 226.870 185.085 ;
        RECT 227.040 184.010 227.310 184.915 ;
        RECT 227.480 184.325 227.810 185.085 ;
        RECT 227.990 184.155 228.160 184.915 ;
        RECT 226.580 182.535 226.870 183.260 ;
        RECT 227.040 183.210 227.210 184.010 ;
        RECT 227.495 183.985 228.160 184.155 ;
        RECT 228.420 184.010 228.690 184.915 ;
        RECT 228.860 184.325 229.190 185.085 ;
        RECT 229.370 184.155 229.540 184.915 ;
        RECT 227.495 183.840 227.665 183.985 ;
        RECT 227.380 183.510 227.665 183.840 ;
        RECT 227.495 183.255 227.665 183.510 ;
        RECT 227.900 183.435 228.230 183.805 ;
        RECT 227.040 182.705 227.300 183.210 ;
        RECT 227.495 183.085 228.160 183.255 ;
        RECT 227.480 182.535 227.810 182.915 ;
        RECT 227.990 182.705 228.160 183.085 ;
        RECT 228.420 183.210 228.590 184.010 ;
        RECT 228.875 183.985 229.540 184.155 ;
        RECT 229.800 184.010 230.070 184.915 ;
        RECT 230.240 184.325 230.570 185.085 ;
        RECT 230.750 184.155 230.920 184.915 ;
        RECT 228.875 183.840 229.045 183.985 ;
        RECT 228.760 183.510 229.045 183.840 ;
        RECT 228.875 183.255 229.045 183.510 ;
        RECT 229.280 183.435 229.610 183.805 ;
        RECT 228.420 182.705 228.680 183.210 ;
        RECT 228.875 183.085 229.540 183.255 ;
        RECT 228.860 182.535 229.190 182.915 ;
        RECT 229.370 182.705 229.540 183.085 ;
        RECT 229.800 183.210 229.970 184.010 ;
        RECT 230.255 183.985 230.920 184.155 ;
        RECT 231.180 184.010 231.450 184.915 ;
        RECT 231.620 184.325 231.950 185.085 ;
        RECT 232.130 184.155 232.300 184.915 ;
        RECT 230.255 183.840 230.425 183.985 ;
        RECT 230.140 183.510 230.425 183.840 ;
        RECT 230.255 183.255 230.425 183.510 ;
        RECT 230.660 183.435 230.990 183.805 ;
        RECT 229.800 182.705 230.060 183.210 ;
        RECT 230.255 183.085 230.920 183.255 ;
        RECT 230.240 182.535 230.570 182.915 ;
        RECT 230.750 182.705 230.920 183.085 ;
        RECT 231.180 183.210 231.350 184.010 ;
        RECT 231.635 183.985 232.300 184.155 ;
        RECT 232.560 184.010 232.830 184.915 ;
        RECT 233.000 184.325 233.330 185.085 ;
        RECT 233.510 184.155 233.680 184.915 ;
        RECT 231.635 183.840 231.805 183.985 ;
        RECT 231.520 183.510 231.805 183.840 ;
        RECT 231.635 183.255 231.805 183.510 ;
        RECT 232.040 183.435 232.370 183.805 ;
        RECT 231.180 182.705 231.440 183.210 ;
        RECT 231.635 183.085 232.300 183.255 ;
        RECT 231.620 182.535 231.950 182.915 ;
        RECT 232.130 182.705 232.300 183.085 ;
        RECT 232.560 183.210 232.730 184.010 ;
        RECT 233.015 183.985 233.680 184.155 ;
        RECT 234.860 183.995 236.070 185.085 ;
        RECT 233.015 183.840 233.185 183.985 ;
        RECT 232.900 183.510 233.185 183.840 ;
        RECT 233.015 183.255 233.185 183.510 ;
        RECT 233.420 183.435 233.750 183.805 ;
        RECT 234.860 183.455 235.380 183.995 ;
        RECT 235.550 183.285 236.070 183.825 ;
        RECT 232.560 182.705 232.820 183.210 ;
        RECT 233.015 183.085 233.680 183.255 ;
        RECT 233.000 182.535 233.330 182.915 ;
        RECT 233.510 182.705 233.680 183.085 ;
        RECT 234.860 182.535 236.070 183.285 ;
        RECT 162.095 182.365 236.155 182.535 ;
        RECT 162.180 181.615 163.390 182.365 ;
        RECT 164.635 181.715 164.965 182.180 ;
        RECT 165.135 181.895 165.305 182.365 ;
        RECT 165.475 181.715 165.805 182.195 ;
        RECT 162.180 181.075 162.700 181.615 ;
        RECT 164.635 181.545 165.805 181.715 ;
        RECT 102.225 180.620 155.700 181.020 ;
        RECT 162.870 180.905 163.390 181.445 ;
        RECT 164.480 181.165 165.125 181.375 ;
        RECT 165.295 181.165 165.865 181.375 ;
        RECT 166.035 180.995 166.205 182.195 ;
        RECT 166.745 181.795 166.915 182.000 ;
        RECT 62.895 180.305 99.045 180.475 ;
        RECT 9.330 178.450 52.060 178.620 ;
        RECT 9.330 168.690 9.500 178.450 ;
        RECT 10.230 177.760 12.230 177.930 ;
        RECT 12.520 177.760 14.520 177.930 ;
        RECT 14.810 177.760 16.810 177.930 ;
        RECT 17.100 177.760 19.100 177.930 ;
        RECT 19.390 177.760 21.390 177.930 ;
        RECT 21.680 177.760 23.680 177.930 ;
        RECT 23.970 177.760 25.970 177.930 ;
        RECT 26.260 177.760 28.260 177.930 ;
        RECT 28.550 177.760 30.550 177.930 ;
        RECT 30.840 177.760 32.840 177.930 ;
        RECT 33.130 177.760 35.130 177.930 ;
        RECT 35.420 177.760 37.420 177.930 ;
        RECT 37.710 177.760 39.710 177.930 ;
        RECT 40.000 177.760 42.000 177.930 ;
        RECT 42.290 177.760 44.290 177.930 ;
        RECT 44.580 177.760 46.580 177.930 ;
        RECT 46.870 177.760 48.870 177.930 ;
        RECT 49.160 177.760 51.160 177.930 ;
        RECT 10.000 169.550 10.170 177.590 ;
        RECT 12.290 169.550 12.460 177.590 ;
        RECT 14.580 169.550 14.750 177.590 ;
        RECT 16.870 169.550 17.040 177.590 ;
        RECT 19.160 169.550 19.330 177.590 ;
        RECT 21.450 169.550 21.620 177.590 ;
        RECT 23.740 169.550 23.910 177.590 ;
        RECT 26.030 169.550 26.200 177.590 ;
        RECT 28.320 169.550 28.490 177.590 ;
        RECT 30.610 169.550 30.780 177.590 ;
        RECT 32.900 169.550 33.070 177.590 ;
        RECT 35.190 169.550 35.360 177.590 ;
        RECT 37.480 169.550 37.650 177.590 ;
        RECT 39.770 169.550 39.940 177.590 ;
        RECT 42.060 169.550 42.230 177.590 ;
        RECT 44.350 169.550 44.520 177.590 ;
        RECT 46.640 169.550 46.810 177.590 ;
        RECT 48.930 169.550 49.100 177.590 ;
        RECT 51.220 169.550 51.390 177.590 ;
        RECT 10.230 169.210 12.230 169.380 ;
        RECT 12.520 169.210 14.520 169.380 ;
        RECT 14.810 169.210 16.810 169.380 ;
        RECT 17.100 169.210 19.100 169.380 ;
        RECT 19.390 169.210 21.390 169.380 ;
        RECT 21.680 169.210 23.680 169.380 ;
        RECT 23.970 169.210 25.970 169.380 ;
        RECT 26.260 169.210 28.260 169.380 ;
        RECT 28.550 169.210 30.550 169.380 ;
        RECT 30.840 169.210 32.840 169.380 ;
        RECT 33.130 169.210 35.130 169.380 ;
        RECT 35.420 169.210 37.420 169.380 ;
        RECT 37.710 169.210 39.710 169.380 ;
        RECT 40.000 169.210 42.000 169.380 ;
        RECT 42.290 169.210 44.290 169.380 ;
        RECT 44.580 169.210 46.580 169.380 ;
        RECT 46.870 169.210 48.870 169.380 ;
        RECT 49.160 169.210 51.160 169.380 ;
        RECT 51.890 168.690 52.060 178.450 ;
        RECT 62.895 177.455 63.425 180.305 ;
        RECT 64.155 179.615 80.155 179.785 ;
        RECT 63.925 178.360 64.095 179.400 ;
        RECT 80.215 178.360 80.385 179.400 ;
        RECT 64.155 177.975 80.155 178.145 ;
        RECT 80.885 177.455 81.055 180.305 ;
        RECT 81.785 179.615 97.785 179.785 ;
        RECT 81.555 178.360 81.725 179.400 ;
        RECT 97.845 178.360 98.015 179.400 ;
        RECT 81.785 177.975 97.785 178.145 ;
        RECT 98.515 177.455 99.045 180.305 ;
        RECT 62.895 177.285 99.045 177.455 ;
        RECT 62.895 174.435 63.425 177.285 ;
        RECT 64.155 176.595 80.155 176.765 ;
        RECT 63.925 175.340 64.095 176.380 ;
        RECT 80.215 175.340 80.385 176.380 ;
        RECT 64.155 174.955 80.155 175.125 ;
        RECT 80.885 174.435 81.055 177.285 ;
        RECT 81.785 176.595 97.785 176.765 ;
        RECT 81.555 175.340 81.725 176.380 ;
        RECT 97.845 175.340 98.015 176.380 ;
        RECT 81.785 174.955 97.785 175.125 ;
        RECT 98.515 174.435 99.045 177.285 ;
        RECT 62.895 174.265 99.045 174.435 ;
        RECT 62.895 171.415 63.425 174.265 ;
        RECT 63.925 173.575 80.385 173.745 ;
        RECT 63.925 172.105 64.155 173.575 ;
        RECT 80.155 172.105 80.385 173.575 ;
        RECT 63.925 171.935 80.385 172.105 ;
        RECT 80.885 171.415 81.055 174.265 ;
        RECT 81.555 173.575 98.015 173.745 ;
        RECT 81.555 172.105 81.785 173.575 ;
        RECT 97.785 172.105 98.015 173.575 ;
        RECT 81.555 171.935 98.015 172.105 ;
        RECT 98.515 171.415 99.045 174.265 ;
        RECT 113.860 176.355 151.710 176.885 ;
        RECT 62.895 170.885 99.045 171.415 ;
        RECT 102.740 172.330 110.970 172.500 ;
        RECT 9.330 168.520 52.060 168.690 ;
        RECT 9.330 167.860 51.780 168.030 ;
        RECT 9.330 158.100 9.500 167.860 ;
        RECT 10.290 167.170 12.290 167.340 ;
        RECT 12.580 167.170 14.580 167.340 ;
        RECT 10.060 158.960 10.230 167.000 ;
        RECT 12.350 158.960 12.520 167.000 ;
        RECT 14.640 158.960 14.810 167.000 ;
        RECT 10.290 158.620 12.290 158.790 ;
        RECT 12.580 158.620 14.580 158.790 ;
        RECT 15.370 158.100 15.540 167.860 ;
        RECT 16.330 167.170 18.330 167.340 ;
        RECT 18.620 167.170 20.620 167.340 ;
        RECT 16.100 158.960 16.270 167.000 ;
        RECT 18.390 158.960 18.560 167.000 ;
        RECT 20.680 158.960 20.850 167.000 ;
        RECT 16.330 158.620 18.330 158.790 ;
        RECT 18.620 158.620 20.620 158.790 ;
        RECT 21.410 158.100 21.580 167.860 ;
        RECT 22.370 167.170 24.370 167.340 ;
        RECT 24.660 167.170 26.660 167.340 ;
        RECT 22.140 158.960 22.310 167.000 ;
        RECT 24.430 158.960 24.600 167.000 ;
        RECT 26.720 158.960 26.890 167.000 ;
        RECT 22.370 158.620 24.370 158.790 ;
        RECT 24.660 158.620 26.660 158.790 ;
        RECT 27.450 158.100 27.620 167.860 ;
        RECT 28.410 167.170 30.410 167.340 ;
        RECT 30.700 167.170 32.700 167.340 ;
        RECT 28.180 158.960 28.350 167.000 ;
        RECT 30.470 158.960 30.640 167.000 ;
        RECT 32.760 158.960 32.930 167.000 ;
        RECT 28.410 158.620 30.410 158.790 ;
        RECT 30.700 158.620 32.700 158.790 ;
        RECT 33.490 158.100 33.660 167.860 ;
        RECT 34.450 167.170 36.450 167.340 ;
        RECT 36.740 167.170 38.740 167.340 ;
        RECT 34.220 158.960 34.390 167.000 ;
        RECT 36.510 158.960 36.680 167.000 ;
        RECT 38.800 158.960 38.970 167.000 ;
        RECT 34.450 158.620 36.450 158.790 ;
        RECT 36.740 158.620 38.740 158.790 ;
        RECT 39.530 158.100 39.700 167.860 ;
        RECT 40.490 167.170 42.490 167.340 ;
        RECT 42.780 167.170 44.780 167.340 ;
        RECT 40.260 158.960 40.430 167.000 ;
        RECT 42.550 158.960 42.720 167.000 ;
        RECT 44.840 158.960 45.010 167.000 ;
        RECT 40.490 158.620 42.490 158.790 ;
        RECT 42.780 158.620 44.780 158.790 ;
        RECT 45.570 158.100 45.740 167.860 ;
        RECT 46.530 167.170 48.530 167.340 ;
        RECT 48.820 167.170 50.820 167.340 ;
        RECT 46.300 158.960 46.470 167.000 ;
        RECT 48.590 158.960 48.760 167.000 ;
        RECT 50.880 158.960 51.050 167.000 ;
        RECT 46.530 158.620 48.530 158.790 ;
        RECT 48.820 158.620 50.820 158.790 ;
        RECT 51.610 158.100 51.780 167.860 ;
        RECT 9.330 157.930 51.780 158.100 ;
        RECT 9.330 148.170 9.500 157.930 ;
        RECT 10.290 157.240 12.290 157.410 ;
        RECT 12.580 157.240 14.580 157.410 ;
        RECT 10.060 149.030 10.230 157.070 ;
        RECT 12.350 149.030 12.520 157.070 ;
        RECT 14.640 149.030 14.810 157.070 ;
        RECT 10.290 148.690 12.290 148.860 ;
        RECT 12.580 148.690 14.580 148.860 ;
        RECT 15.370 148.170 15.540 157.930 ;
        RECT 16.330 157.240 18.330 157.410 ;
        RECT 18.620 157.240 20.620 157.410 ;
        RECT 16.100 149.030 16.270 157.070 ;
        RECT 18.390 149.030 18.560 157.070 ;
        RECT 20.680 149.030 20.850 157.070 ;
        RECT 16.330 148.690 18.330 148.860 ;
        RECT 18.620 148.690 20.620 148.860 ;
        RECT 21.410 148.170 21.580 157.930 ;
        RECT 22.370 157.240 24.370 157.410 ;
        RECT 24.660 157.240 26.660 157.410 ;
        RECT 22.140 149.030 22.310 157.070 ;
        RECT 24.430 149.030 24.600 157.070 ;
        RECT 26.720 149.030 26.890 157.070 ;
        RECT 22.370 148.690 24.370 148.860 ;
        RECT 24.660 148.690 26.660 148.860 ;
        RECT 27.450 148.170 27.620 157.930 ;
        RECT 28.410 157.240 30.410 157.410 ;
        RECT 30.700 157.240 32.700 157.410 ;
        RECT 28.180 149.030 28.350 157.070 ;
        RECT 30.470 149.030 30.640 157.070 ;
        RECT 32.760 149.030 32.930 157.070 ;
        RECT 28.410 148.690 30.410 148.860 ;
        RECT 30.700 148.690 32.700 148.860 ;
        RECT 33.490 148.170 33.660 157.930 ;
        RECT 34.450 157.240 36.450 157.410 ;
        RECT 36.740 157.240 38.740 157.410 ;
        RECT 34.220 149.030 34.390 157.070 ;
        RECT 36.510 149.030 36.680 157.070 ;
        RECT 38.800 149.030 38.970 157.070 ;
        RECT 34.450 148.690 36.450 148.860 ;
        RECT 36.740 148.690 38.740 148.860 ;
        RECT 39.530 148.170 39.700 157.930 ;
        RECT 40.490 157.240 42.490 157.410 ;
        RECT 42.780 157.240 44.780 157.410 ;
        RECT 40.260 149.030 40.430 157.070 ;
        RECT 42.550 149.030 42.720 157.070 ;
        RECT 44.840 149.030 45.010 157.070 ;
        RECT 40.490 148.690 42.490 148.860 ;
        RECT 42.780 148.690 44.780 148.860 ;
        RECT 45.570 148.170 45.740 157.930 ;
        RECT 46.530 157.240 48.530 157.410 ;
        RECT 48.820 157.240 50.820 157.410 ;
        RECT 46.300 149.030 46.470 157.070 ;
        RECT 48.590 149.030 48.760 157.070 ;
        RECT 50.880 149.030 51.050 157.070 ;
        RECT 46.530 148.690 48.530 148.860 ;
        RECT 48.820 148.690 50.820 148.860 ;
        RECT 51.610 148.170 51.780 157.930 ;
        RECT 9.330 148.000 51.780 148.170 ;
        RECT 64.100 166.025 96.940 166.425 ;
        RECT 23.195 143.155 58.705 143.745 ;
        RECT 23.195 140.745 23.785 143.155 ;
        RECT 24.515 142.465 32.515 142.635 ;
        RECT 32.805 142.465 40.805 142.635 ;
        RECT 41.095 142.465 49.095 142.635 ;
        RECT 49.385 142.465 57.385 142.635 ;
        RECT 24.285 141.255 24.455 142.295 ;
        RECT 32.575 141.255 32.745 142.295 ;
        RECT 40.865 141.255 41.035 142.295 ;
        RECT 49.155 141.255 49.325 142.295 ;
        RECT 57.445 141.255 57.615 142.295 ;
        RECT 24.515 140.915 32.515 141.085 ;
        RECT 32.805 140.915 40.805 141.085 ;
        RECT 41.095 140.915 49.095 141.085 ;
        RECT 49.385 140.915 57.385 141.085 ;
        RECT 23.195 139.705 24.455 140.745 ;
        RECT 32.575 139.705 32.745 140.745 ;
        RECT 40.865 139.705 41.035 140.745 ;
        RECT 49.155 139.705 49.325 140.745 ;
        RECT 57.445 139.705 57.615 140.745 ;
        RECT 23.195 139.195 23.785 139.705 ;
        RECT 24.515 139.365 32.515 139.535 ;
        RECT 32.805 139.365 40.805 139.535 ;
        RECT 41.095 139.365 49.095 139.535 ;
        RECT 49.385 139.365 57.385 139.535 ;
        RECT 9.430 137.955 20.720 138.485 ;
        RECT 9.430 135.195 9.960 137.955 ;
        RECT 10.995 137.265 11.995 137.435 ;
        RECT 10.765 136.055 10.935 137.095 ;
        RECT 12.055 136.055 12.225 137.095 ;
        RECT 13.030 135.195 13.200 137.955 ;
        RECT 13.930 137.265 14.930 137.435 ;
        RECT 15.220 137.265 16.220 137.435 ;
        RECT 13.700 136.055 13.870 137.095 ;
        RECT 14.990 136.055 15.160 137.095 ;
        RECT 16.280 136.055 16.450 137.095 ;
        RECT 16.950 135.195 17.120 137.955 ;
        RECT 18.155 137.265 19.155 137.435 ;
        RECT 17.925 136.055 18.095 137.095 ;
        RECT 19.215 136.055 19.385 137.095 ;
        RECT 20.190 135.195 20.720 137.955 ;
        RECT 9.430 134.665 20.720 135.195 ;
        RECT 23.195 138.155 24.455 139.195 ;
        RECT 32.575 138.155 32.745 139.195 ;
        RECT 40.865 138.155 41.035 139.195 ;
        RECT 49.155 138.155 49.325 139.195 ;
        RECT 57.445 138.155 57.615 139.195 ;
        RECT 23.195 135.745 23.785 138.155 ;
        RECT 24.515 137.815 32.515 137.985 ;
        RECT 32.805 137.815 40.805 137.985 ;
        RECT 41.095 137.815 49.095 137.985 ;
        RECT 49.385 137.815 57.385 137.985 ;
        RECT 24.285 136.605 24.455 137.645 ;
        RECT 32.575 136.605 32.745 137.645 ;
        RECT 40.865 136.605 41.035 137.645 ;
        RECT 49.155 136.605 49.325 137.645 ;
        RECT 57.445 136.605 57.615 137.645 ;
        RECT 24.515 136.265 32.515 136.435 ;
        RECT 32.805 136.265 40.805 136.435 ;
        RECT 41.095 136.265 49.095 136.435 ;
        RECT 49.385 136.265 57.385 136.435 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 23.195 135.155 58.705 135.745 ;
        RECT 64.100 133.985 64.500 166.025 ;
        RECT 69.635 160.720 91.405 160.890 ;
        RECT 69.635 139.290 69.805 160.720 ;
        RECT 71.220 158.800 89.820 159.305 ;
        RECT 71.220 156.090 71.725 158.800 ;
        RECT 72.035 158.130 74.125 158.490 ;
        RECT 72.035 156.760 72.395 158.130 ;
        RECT 72.685 157.050 73.475 157.840 ;
        RECT 73.765 156.760 74.125 158.130 ;
        RECT 72.035 156.400 74.125 156.760 ;
        RECT 74.435 156.090 75.445 158.800 ;
        RECT 75.755 158.130 77.845 158.490 ;
        RECT 75.755 156.760 76.115 158.130 ;
        RECT 76.405 157.050 77.195 157.840 ;
        RECT 77.485 156.760 77.845 158.130 ;
        RECT 75.755 156.400 77.845 156.760 ;
        RECT 78.155 156.090 79.165 158.800 ;
        RECT 79.475 158.130 81.565 158.490 ;
        RECT 79.475 156.760 79.835 158.130 ;
        RECT 80.125 157.050 80.915 157.840 ;
        RECT 81.205 156.760 81.565 158.130 ;
        RECT 79.475 156.400 81.565 156.760 ;
        RECT 81.875 156.090 82.885 158.800 ;
        RECT 83.195 158.130 85.285 158.490 ;
        RECT 83.195 156.760 83.555 158.130 ;
        RECT 83.845 157.050 84.635 157.840 ;
        RECT 84.925 156.760 85.285 158.130 ;
        RECT 83.195 156.400 85.285 156.760 ;
        RECT 85.595 156.090 86.605 158.800 ;
        RECT 86.915 158.130 89.005 158.490 ;
        RECT 86.915 156.760 87.275 158.130 ;
        RECT 87.565 157.050 88.355 157.840 ;
        RECT 88.645 156.760 89.005 158.130 ;
        RECT 86.915 156.400 89.005 156.760 ;
        RECT 89.315 156.090 89.820 158.800 ;
        RECT 71.220 155.080 89.820 156.090 ;
        RECT 71.220 152.370 71.725 155.080 ;
        RECT 72.035 154.410 74.125 154.770 ;
        RECT 72.035 153.040 72.395 154.410 ;
        RECT 72.685 153.330 73.475 154.120 ;
        RECT 73.765 153.040 74.125 154.410 ;
        RECT 72.035 152.680 74.125 153.040 ;
        RECT 74.435 152.370 75.445 155.080 ;
        RECT 75.755 154.410 77.845 154.770 ;
        RECT 75.755 153.040 76.115 154.410 ;
        RECT 76.405 153.330 77.195 154.120 ;
        RECT 77.485 153.040 77.845 154.410 ;
        RECT 75.755 152.680 77.845 153.040 ;
        RECT 78.155 152.370 79.165 155.080 ;
        RECT 79.475 154.410 81.565 154.770 ;
        RECT 79.475 153.040 79.835 154.410 ;
        RECT 80.125 153.330 80.915 154.120 ;
        RECT 81.205 153.040 81.565 154.410 ;
        RECT 79.475 152.680 81.565 153.040 ;
        RECT 81.875 152.370 82.885 155.080 ;
        RECT 83.195 154.410 85.285 154.770 ;
        RECT 83.195 153.040 83.555 154.410 ;
        RECT 83.845 153.330 84.635 154.120 ;
        RECT 84.925 153.040 85.285 154.410 ;
        RECT 83.195 152.680 85.285 153.040 ;
        RECT 85.595 152.370 86.605 155.080 ;
        RECT 86.915 154.410 89.005 154.770 ;
        RECT 86.915 153.040 87.275 154.410 ;
        RECT 87.565 153.330 88.355 154.120 ;
        RECT 88.645 153.040 89.005 154.410 ;
        RECT 86.915 152.680 89.005 153.040 ;
        RECT 89.315 152.370 89.820 155.080 ;
        RECT 71.220 151.360 89.820 152.370 ;
        RECT 71.220 148.650 71.725 151.360 ;
        RECT 72.035 150.690 74.125 151.050 ;
        RECT 72.035 149.320 72.395 150.690 ;
        RECT 72.685 149.610 73.475 150.400 ;
        RECT 73.765 149.320 74.125 150.690 ;
        RECT 72.035 148.960 74.125 149.320 ;
        RECT 74.435 148.650 75.445 151.360 ;
        RECT 75.755 150.690 77.845 151.050 ;
        RECT 75.755 149.320 76.115 150.690 ;
        RECT 76.405 149.610 77.195 150.400 ;
        RECT 77.485 149.320 77.845 150.690 ;
        RECT 75.755 148.960 77.845 149.320 ;
        RECT 78.155 148.650 79.165 151.360 ;
        RECT 79.475 150.690 81.565 151.050 ;
        RECT 79.475 149.320 79.835 150.690 ;
        RECT 80.125 149.610 80.915 150.400 ;
        RECT 81.205 149.320 81.565 150.690 ;
        RECT 79.475 148.960 81.565 149.320 ;
        RECT 81.875 148.650 82.885 151.360 ;
        RECT 83.195 150.690 85.285 151.050 ;
        RECT 83.195 149.320 83.555 150.690 ;
        RECT 83.845 149.610 84.635 150.400 ;
        RECT 84.925 149.320 85.285 150.690 ;
        RECT 83.195 148.960 85.285 149.320 ;
        RECT 85.595 148.650 86.605 151.360 ;
        RECT 86.915 150.690 89.005 151.050 ;
        RECT 86.915 149.320 87.275 150.690 ;
        RECT 87.565 149.610 88.355 150.400 ;
        RECT 88.645 149.320 89.005 150.690 ;
        RECT 86.915 148.960 89.005 149.320 ;
        RECT 89.315 148.650 89.820 151.360 ;
        RECT 71.220 147.640 89.820 148.650 ;
        RECT 71.220 144.930 71.725 147.640 ;
        RECT 72.035 146.970 74.125 147.330 ;
        RECT 72.035 145.600 72.395 146.970 ;
        RECT 72.685 145.890 73.475 146.680 ;
        RECT 73.765 145.600 74.125 146.970 ;
        RECT 72.035 145.240 74.125 145.600 ;
        RECT 74.435 144.930 75.445 147.640 ;
        RECT 75.755 146.970 77.845 147.330 ;
        RECT 75.755 145.600 76.115 146.970 ;
        RECT 76.405 145.890 77.195 146.680 ;
        RECT 77.485 145.600 77.845 146.970 ;
        RECT 75.755 145.240 77.845 145.600 ;
        RECT 78.155 144.930 79.165 147.640 ;
        RECT 79.475 146.970 81.565 147.330 ;
        RECT 79.475 145.600 79.835 146.970 ;
        RECT 80.125 145.890 80.915 146.680 ;
        RECT 81.205 145.600 81.565 146.970 ;
        RECT 79.475 145.240 81.565 145.600 ;
        RECT 81.875 144.930 82.885 147.640 ;
        RECT 83.195 146.970 85.285 147.330 ;
        RECT 83.195 145.600 83.555 146.970 ;
        RECT 83.845 145.890 84.635 146.680 ;
        RECT 84.925 145.600 85.285 146.970 ;
        RECT 83.195 145.240 85.285 145.600 ;
        RECT 85.595 144.930 86.605 147.640 ;
        RECT 86.915 146.970 89.005 147.330 ;
        RECT 86.915 145.600 87.275 146.970 ;
        RECT 87.565 145.890 88.355 146.680 ;
        RECT 88.645 145.600 89.005 146.970 ;
        RECT 86.915 145.240 89.005 145.600 ;
        RECT 89.315 144.930 89.820 147.640 ;
        RECT 71.220 143.920 89.820 144.930 ;
        RECT 71.220 141.210 71.725 143.920 ;
        RECT 72.035 143.250 74.125 143.610 ;
        RECT 72.035 141.880 72.395 143.250 ;
        RECT 72.685 142.170 73.475 142.960 ;
        RECT 73.765 141.880 74.125 143.250 ;
        RECT 72.035 141.520 74.125 141.880 ;
        RECT 74.435 141.210 75.445 143.920 ;
        RECT 75.755 143.250 77.845 143.610 ;
        RECT 75.755 141.880 76.115 143.250 ;
        RECT 76.405 142.170 77.195 142.960 ;
        RECT 77.485 141.880 77.845 143.250 ;
        RECT 75.755 141.520 77.845 141.880 ;
        RECT 78.155 141.210 79.165 143.920 ;
        RECT 79.475 143.250 81.565 143.610 ;
        RECT 79.475 141.880 79.835 143.250 ;
        RECT 80.125 142.170 80.915 142.960 ;
        RECT 81.205 141.880 81.565 143.250 ;
        RECT 79.475 141.520 81.565 141.880 ;
        RECT 81.875 141.210 82.885 143.920 ;
        RECT 83.195 143.250 85.285 143.610 ;
        RECT 83.195 141.880 83.555 143.250 ;
        RECT 83.845 142.170 84.635 142.960 ;
        RECT 84.925 141.880 85.285 143.250 ;
        RECT 83.195 141.520 85.285 141.880 ;
        RECT 85.595 141.210 86.605 143.920 ;
        RECT 86.915 143.250 89.005 143.610 ;
        RECT 86.915 141.880 87.275 143.250 ;
        RECT 87.565 142.170 88.355 142.960 ;
        RECT 88.645 141.880 89.005 143.250 ;
        RECT 86.915 141.520 89.005 141.880 ;
        RECT 89.315 141.210 89.820 143.920 ;
        RECT 71.220 140.705 89.820 141.210 ;
        RECT 91.235 139.290 91.405 160.720 ;
        RECT 69.635 139.120 91.405 139.290 ;
        RECT 96.540 133.985 96.940 166.025 ;
        RECT 102.740 162.570 102.910 172.330 ;
        RECT 103.695 171.640 104.695 171.810 ;
        RECT 104.985 171.640 105.985 171.810 ;
        RECT 103.465 163.430 103.635 171.470 ;
        RECT 104.755 163.430 104.925 171.470 ;
        RECT 106.045 163.430 106.215 171.470 ;
        RECT 103.695 163.090 104.695 163.260 ;
        RECT 104.985 163.090 105.985 163.260 ;
        RECT 106.770 162.570 106.940 172.330 ;
        RECT 107.725 171.640 108.725 171.810 ;
        RECT 109.015 171.640 110.015 171.810 ;
        RECT 107.495 163.430 107.665 171.470 ;
        RECT 108.785 163.430 108.955 171.470 ;
        RECT 110.075 163.430 110.245 171.470 ;
        RECT 107.725 163.090 108.725 163.260 ;
        RECT 109.015 163.090 110.015 163.260 ;
        RECT 110.800 162.570 110.970 172.330 ;
        RECT 113.860 166.595 114.390 176.355 ;
        RECT 115.180 175.665 115.680 175.835 ;
        RECT 115.970 175.665 116.470 175.835 ;
        RECT 116.760 175.665 117.260 175.835 ;
        RECT 117.550 175.665 118.050 175.835 ;
        RECT 114.950 167.455 115.120 175.495 ;
        RECT 115.740 167.455 115.910 175.495 ;
        RECT 116.530 167.455 116.700 175.495 ;
        RECT 117.320 167.455 117.490 175.495 ;
        RECT 118.110 167.455 118.280 175.495 ;
        RECT 115.180 167.115 115.680 167.285 ;
        RECT 115.970 167.115 116.470 167.285 ;
        RECT 116.760 167.115 117.260 167.285 ;
        RECT 117.550 167.115 118.050 167.285 ;
        RECT 118.840 166.595 119.010 176.355 ;
        RECT 119.800 175.665 120.300 175.835 ;
        RECT 120.590 175.665 121.090 175.835 ;
        RECT 121.380 175.665 121.880 175.835 ;
        RECT 122.170 175.665 122.670 175.835 ;
        RECT 119.570 167.455 119.740 175.495 ;
        RECT 120.360 167.455 120.530 175.495 ;
        RECT 121.150 167.455 121.320 175.495 ;
        RECT 121.940 167.455 122.110 175.495 ;
        RECT 122.730 167.455 122.900 175.495 ;
        RECT 119.800 167.115 120.300 167.285 ;
        RECT 120.590 167.115 121.090 167.285 ;
        RECT 121.380 167.115 121.880 167.285 ;
        RECT 122.170 167.115 122.670 167.285 ;
        RECT 123.460 166.595 123.630 176.355 ;
        RECT 124.420 175.665 124.920 175.835 ;
        RECT 125.210 175.665 125.710 175.835 ;
        RECT 126.000 175.665 126.500 175.835 ;
        RECT 126.790 175.665 127.290 175.835 ;
        RECT 124.190 167.455 124.360 175.495 ;
        RECT 124.980 167.455 125.150 175.495 ;
        RECT 125.770 167.455 125.940 175.495 ;
        RECT 126.560 167.455 126.730 175.495 ;
        RECT 127.350 167.455 127.520 175.495 ;
        RECT 124.420 167.115 124.920 167.285 ;
        RECT 125.210 167.115 125.710 167.285 ;
        RECT 126.000 167.115 126.500 167.285 ;
        RECT 126.790 167.115 127.290 167.285 ;
        RECT 128.080 166.595 128.250 176.355 ;
        RECT 129.040 175.665 129.540 175.835 ;
        RECT 129.830 175.665 130.330 175.835 ;
        RECT 130.620 175.665 131.120 175.835 ;
        RECT 131.410 175.665 131.910 175.835 ;
        RECT 128.810 167.455 128.980 175.495 ;
        RECT 129.600 167.455 129.770 175.495 ;
        RECT 130.390 167.455 130.560 175.495 ;
        RECT 131.180 167.455 131.350 175.495 ;
        RECT 131.970 167.455 132.140 175.495 ;
        RECT 129.040 167.115 129.540 167.285 ;
        RECT 129.830 167.115 130.330 167.285 ;
        RECT 130.620 167.115 131.120 167.285 ;
        RECT 131.410 167.115 131.910 167.285 ;
        RECT 132.700 166.595 132.870 176.355 ;
        RECT 133.660 175.665 134.160 175.835 ;
        RECT 134.450 175.665 134.950 175.835 ;
        RECT 135.240 175.665 135.740 175.835 ;
        RECT 136.030 175.665 136.530 175.835 ;
        RECT 133.430 167.455 133.600 175.495 ;
        RECT 134.220 167.455 134.390 175.495 ;
        RECT 135.010 167.455 135.180 175.495 ;
        RECT 135.800 167.455 135.970 175.495 ;
        RECT 136.590 167.455 136.760 175.495 ;
        RECT 133.660 167.115 134.160 167.285 ;
        RECT 134.450 167.115 134.950 167.285 ;
        RECT 135.240 167.115 135.740 167.285 ;
        RECT 136.030 167.115 136.530 167.285 ;
        RECT 137.320 166.595 137.490 176.355 ;
        RECT 138.280 175.665 138.780 175.835 ;
        RECT 139.070 175.665 139.570 175.835 ;
        RECT 139.860 175.665 140.360 175.835 ;
        RECT 140.650 175.665 141.150 175.835 ;
        RECT 138.050 167.455 138.220 175.495 ;
        RECT 138.840 167.455 139.010 175.495 ;
        RECT 139.630 167.455 139.800 175.495 ;
        RECT 140.420 167.455 140.590 175.495 ;
        RECT 141.210 167.455 141.380 175.495 ;
        RECT 138.280 167.115 138.780 167.285 ;
        RECT 139.070 167.115 139.570 167.285 ;
        RECT 139.860 167.115 140.360 167.285 ;
        RECT 140.650 167.115 141.150 167.285 ;
        RECT 141.940 166.595 142.110 176.355 ;
        RECT 142.900 175.665 143.400 175.835 ;
        RECT 143.690 175.665 144.190 175.835 ;
        RECT 144.480 175.665 144.980 175.835 ;
        RECT 145.270 175.665 145.770 175.835 ;
        RECT 142.670 167.455 142.840 175.495 ;
        RECT 143.460 167.455 143.630 175.495 ;
        RECT 144.250 167.455 144.420 175.495 ;
        RECT 145.040 167.455 145.210 175.495 ;
        RECT 145.830 167.455 146.000 175.495 ;
        RECT 142.900 167.115 143.400 167.285 ;
        RECT 143.690 167.115 144.190 167.285 ;
        RECT 144.480 167.115 144.980 167.285 ;
        RECT 145.270 167.115 145.770 167.285 ;
        RECT 146.560 166.595 146.730 176.355 ;
        RECT 147.520 175.665 148.020 175.835 ;
        RECT 148.310 175.665 148.810 175.835 ;
        RECT 149.100 175.665 149.600 175.835 ;
        RECT 149.890 175.665 150.390 175.835 ;
        RECT 147.290 167.455 147.460 175.495 ;
        RECT 148.080 167.455 148.250 175.495 ;
        RECT 148.870 167.455 149.040 175.495 ;
        RECT 149.660 167.455 149.830 175.495 ;
        RECT 150.450 167.455 150.620 175.495 ;
        RECT 147.520 167.115 148.020 167.285 ;
        RECT 148.310 167.115 148.810 167.285 ;
        RECT 149.100 167.115 149.600 167.285 ;
        RECT 149.890 167.115 150.390 167.285 ;
        RECT 151.180 166.595 151.710 176.355 ;
        RECT 113.860 166.065 151.710 166.595 ;
        RECT 102.740 162.400 110.970 162.570 ;
        RECT 102.740 158.640 102.910 162.400 ;
        RECT 103.465 159.500 103.635 161.540 ;
        RECT 104.755 159.500 104.925 161.540 ;
        RECT 106.045 159.500 106.215 161.540 ;
        RECT 103.695 159.160 104.695 159.330 ;
        RECT 104.985 159.160 105.985 159.330 ;
        RECT 106.770 158.640 106.940 162.400 ;
        RECT 107.495 159.500 107.665 161.540 ;
        RECT 108.785 159.500 108.955 161.540 ;
        RECT 110.075 159.500 110.245 161.540 ;
        RECT 107.725 159.160 108.725 159.330 ;
        RECT 109.015 159.160 110.015 159.330 ;
        RECT 110.800 158.640 110.970 162.400 ;
        RECT 102.740 158.470 110.970 158.640 ;
        RECT 116.015 157.500 149.445 158.030 ;
        RECT 102.740 155.775 110.970 155.945 ;
        RECT 102.740 151.925 102.910 155.775 ;
        RECT 103.695 155.085 104.695 155.255 ;
        RECT 104.985 155.085 105.985 155.255 ;
        RECT 103.465 152.830 103.635 154.870 ;
        RECT 104.755 152.830 104.925 154.870 ;
        RECT 106.045 152.830 106.215 154.870 ;
        RECT 106.770 151.925 106.940 155.775 ;
        RECT 107.725 155.085 108.725 155.255 ;
        RECT 109.015 155.085 110.015 155.255 ;
        RECT 107.495 152.830 107.665 154.870 ;
        RECT 108.785 152.830 108.955 154.870 ;
        RECT 110.075 152.830 110.245 154.870 ;
        RECT 110.800 151.925 110.970 155.775 ;
        RECT 102.740 151.755 110.970 151.925 ;
        RECT 102.740 141.905 102.910 151.755 ;
        RECT 103.695 151.065 104.695 151.235 ;
        RECT 104.985 151.065 105.985 151.235 ;
        RECT 103.465 142.810 103.635 150.850 ;
        RECT 104.755 142.810 104.925 150.850 ;
        RECT 106.045 142.810 106.215 150.850 ;
        RECT 103.695 142.425 104.695 142.595 ;
        RECT 104.985 142.425 105.985 142.595 ;
        RECT 106.770 141.905 106.940 151.755 ;
        RECT 107.725 151.065 108.725 151.235 ;
        RECT 109.015 151.065 110.015 151.235 ;
        RECT 107.495 142.810 107.665 150.850 ;
        RECT 108.785 142.810 108.955 150.850 ;
        RECT 110.075 142.810 110.245 150.850 ;
        RECT 107.725 142.425 108.725 142.595 ;
        RECT 109.015 142.425 110.015 142.595 ;
        RECT 110.800 141.905 110.970 151.755 ;
        RECT 102.740 141.735 110.970 141.905 ;
        RECT 116.015 140.250 116.545 157.500 ;
        RECT 117.130 156.135 119.290 156.825 ;
        RECT 117.130 154.965 119.290 155.655 ;
        RECT 117.130 153.795 119.290 154.485 ;
        RECT 117.130 152.625 119.290 153.315 ;
        RECT 117.130 151.455 119.290 152.145 ;
        RECT 117.130 150.285 119.290 150.975 ;
        RECT 117.130 149.115 119.290 149.805 ;
        RECT 117.130 147.945 119.290 148.635 ;
        RECT 117.130 146.775 119.290 147.465 ;
        RECT 117.130 145.605 119.290 146.295 ;
        RECT 117.130 144.435 119.290 145.125 ;
        RECT 117.130 143.265 119.290 143.955 ;
        RECT 117.130 142.095 119.290 142.785 ;
        RECT 117.130 140.925 119.290 141.615 ;
        RECT 119.595 140.250 122.075 157.500 ;
        RECT 122.380 156.135 124.540 156.825 ;
        RECT 125.060 156.135 127.220 156.825 ;
        RECT 122.380 154.965 124.540 155.655 ;
        RECT 125.060 154.965 127.220 155.655 ;
        RECT 122.380 153.795 124.540 154.485 ;
        RECT 125.060 153.795 127.220 154.485 ;
        RECT 122.380 152.625 124.540 153.315 ;
        RECT 125.060 152.625 127.220 153.315 ;
        RECT 122.380 151.455 124.540 152.145 ;
        RECT 125.060 151.455 127.220 152.145 ;
        RECT 122.380 150.285 124.540 150.975 ;
        RECT 125.060 150.285 127.220 150.975 ;
        RECT 122.380 149.115 124.540 149.805 ;
        RECT 125.060 149.115 127.220 149.805 ;
        RECT 122.380 147.945 124.540 148.635 ;
        RECT 125.060 147.945 127.220 148.635 ;
        RECT 122.380 146.775 124.540 147.465 ;
        RECT 125.060 146.775 127.220 147.465 ;
        RECT 122.380 145.605 124.540 146.295 ;
        RECT 125.060 145.605 127.220 146.295 ;
        RECT 122.380 144.435 124.540 145.125 ;
        RECT 125.060 144.435 127.220 145.125 ;
        RECT 122.380 143.265 124.540 143.955 ;
        RECT 125.060 143.265 127.220 143.955 ;
        RECT 122.380 142.095 124.540 142.785 ;
        RECT 125.060 142.095 127.220 142.785 ;
        RECT 122.380 140.925 124.540 141.615 ;
        RECT 125.060 140.925 127.220 141.615 ;
        RECT 127.525 140.250 130.005 157.500 ;
        RECT 130.310 156.135 132.470 156.825 ;
        RECT 132.990 156.135 135.150 156.825 ;
        RECT 130.310 154.965 132.470 155.655 ;
        RECT 132.990 154.965 135.150 155.655 ;
        RECT 130.310 153.795 132.470 154.485 ;
        RECT 132.990 153.795 135.150 154.485 ;
        RECT 130.310 152.625 132.470 153.315 ;
        RECT 132.990 152.625 135.150 153.315 ;
        RECT 130.310 151.455 132.470 152.145 ;
        RECT 132.990 151.455 135.150 152.145 ;
        RECT 130.310 150.285 132.470 150.975 ;
        RECT 132.990 150.285 135.150 150.975 ;
        RECT 130.310 149.115 132.470 149.805 ;
        RECT 132.990 149.115 135.150 149.805 ;
        RECT 130.310 147.945 132.470 148.635 ;
        RECT 132.990 147.945 135.150 148.635 ;
        RECT 130.310 146.775 132.470 147.465 ;
        RECT 132.990 146.775 135.150 147.465 ;
        RECT 130.310 145.605 132.470 146.295 ;
        RECT 132.990 145.605 135.150 146.295 ;
        RECT 130.310 144.435 132.470 145.125 ;
        RECT 132.990 144.435 135.150 145.125 ;
        RECT 130.310 143.265 132.470 143.955 ;
        RECT 132.990 143.265 135.150 143.955 ;
        RECT 130.310 142.095 132.470 142.785 ;
        RECT 132.990 142.095 135.150 142.785 ;
        RECT 130.310 140.925 132.470 141.615 ;
        RECT 132.990 140.925 135.150 141.615 ;
        RECT 135.455 140.250 137.935 157.500 ;
        RECT 138.240 156.135 140.400 156.825 ;
        RECT 140.920 156.135 143.080 156.825 ;
        RECT 138.240 154.965 140.400 155.655 ;
        RECT 140.920 154.965 143.080 155.655 ;
        RECT 138.240 153.795 140.400 154.485 ;
        RECT 140.920 153.795 143.080 154.485 ;
        RECT 138.240 152.625 140.400 153.315 ;
        RECT 140.920 152.625 143.080 153.315 ;
        RECT 138.240 151.455 140.400 152.145 ;
        RECT 140.920 151.455 143.080 152.145 ;
        RECT 138.240 150.285 140.400 150.975 ;
        RECT 140.920 150.285 143.080 150.975 ;
        RECT 138.240 149.115 140.400 149.805 ;
        RECT 140.920 149.115 143.080 149.805 ;
        RECT 138.240 147.945 140.400 148.635 ;
        RECT 140.920 147.945 143.080 148.635 ;
        RECT 138.240 146.775 140.400 147.465 ;
        RECT 140.920 146.775 143.080 147.465 ;
        RECT 138.240 145.605 140.400 146.295 ;
        RECT 140.920 145.605 143.080 146.295 ;
        RECT 138.240 144.435 140.400 145.125 ;
        RECT 140.920 144.435 143.080 145.125 ;
        RECT 138.240 143.265 140.400 143.955 ;
        RECT 140.920 143.265 143.080 143.955 ;
        RECT 138.240 142.095 140.400 142.785 ;
        RECT 140.920 142.095 143.080 142.785 ;
        RECT 138.240 140.925 140.400 141.615 ;
        RECT 140.920 140.925 143.080 141.615 ;
        RECT 143.385 140.250 145.865 157.500 ;
        RECT 146.170 156.135 148.330 156.825 ;
        RECT 146.170 154.965 148.330 155.655 ;
        RECT 146.170 153.795 148.330 154.485 ;
        RECT 146.170 152.625 148.330 153.315 ;
        RECT 146.170 151.455 148.330 152.145 ;
        RECT 146.170 150.285 148.330 150.975 ;
        RECT 146.170 149.115 148.330 149.805 ;
        RECT 146.170 147.945 148.330 148.635 ;
        RECT 146.170 146.775 148.330 147.465 ;
        RECT 146.170 145.605 148.330 146.295 ;
        RECT 146.170 144.435 148.330 145.125 ;
        RECT 146.170 143.265 148.330 143.955 ;
        RECT 146.170 142.095 148.330 142.785 ;
        RECT 146.170 140.925 148.330 141.615 ;
        RECT 148.915 140.250 149.445 157.500 ;
        RECT 116.015 139.720 149.445 140.250 ;
        RECT 64.100 133.585 96.940 133.985 ;
        RECT 138.110 134.130 145.930 134.660 ;
        RECT 138.110 130.280 138.640 134.130 ;
        RECT 139.465 133.440 140.465 133.610 ;
        RECT 140.755 133.440 141.755 133.610 ;
        RECT 139.235 131.185 139.405 133.225 ;
        RECT 140.525 131.185 140.695 133.225 ;
        RECT 141.815 131.185 141.985 133.225 ;
        RECT 142.580 130.280 142.750 134.130 ;
        RECT 143.345 131.185 143.515 133.225 ;
        RECT 144.635 131.185 144.805 133.225 ;
        RECT 143.575 130.800 144.575 130.970 ;
        RECT 145.400 130.280 145.930 134.130 ;
        RECT 138.110 129.750 145.930 130.280 ;
        RECT 138.110 128.410 145.930 128.940 ;
        RECT 138.110 124.650 138.640 128.410 ;
        RECT 139.235 125.510 139.405 127.550 ;
        RECT 140.525 125.510 140.695 127.550 ;
        RECT 141.815 125.510 141.985 127.550 ;
        RECT 139.465 125.170 140.465 125.340 ;
        RECT 140.755 125.170 141.755 125.340 ;
        RECT 142.580 124.650 142.750 128.410 ;
        RECT 143.575 127.720 144.575 127.890 ;
        RECT 143.345 125.510 143.515 127.550 ;
        RECT 144.635 125.510 144.805 127.550 ;
        RECT 145.400 124.650 145.930 128.410 ;
        RECT 10.055 123.725 70.145 124.255 ;
        RECT 10.055 113.875 10.585 123.725 ;
        RECT 11.315 123.035 13.315 123.205 ;
        RECT 13.605 123.035 15.605 123.205 ;
        RECT 11.085 114.780 11.255 122.820 ;
        RECT 13.375 114.780 13.545 122.820 ;
        RECT 15.665 114.780 15.835 122.820 ;
        RECT 11.315 114.395 13.315 114.565 ;
        RECT 13.605 114.395 15.605 114.565 ;
        RECT 16.335 113.875 16.505 123.725 ;
        RECT 17.235 123.035 19.235 123.205 ;
        RECT 19.525 123.035 21.525 123.205 ;
        RECT 17.005 114.780 17.175 122.820 ;
        RECT 19.295 114.780 19.465 122.820 ;
        RECT 21.585 114.780 21.755 122.820 ;
        RECT 17.235 114.395 19.235 114.565 ;
        RECT 19.525 114.395 21.525 114.565 ;
        RECT 22.255 113.875 22.425 123.725 ;
        RECT 23.155 123.035 25.155 123.205 ;
        RECT 25.445 123.035 27.445 123.205 ;
        RECT 22.925 114.780 23.095 122.820 ;
        RECT 25.215 114.780 25.385 122.820 ;
        RECT 27.505 114.780 27.675 122.820 ;
        RECT 23.155 114.395 25.155 114.565 ;
        RECT 25.445 114.395 27.445 114.565 ;
        RECT 28.175 113.875 28.345 123.725 ;
        RECT 29.075 123.035 31.075 123.205 ;
        RECT 31.365 123.035 33.365 123.205 ;
        RECT 28.845 114.780 29.015 122.820 ;
        RECT 31.135 114.780 31.305 122.820 ;
        RECT 33.425 114.780 33.595 122.820 ;
        RECT 29.075 114.395 31.075 114.565 ;
        RECT 31.365 114.395 33.365 114.565 ;
        RECT 34.095 113.875 34.265 123.725 ;
        RECT 34.995 123.035 36.995 123.205 ;
        RECT 37.285 123.035 39.285 123.205 ;
        RECT 34.765 114.780 34.935 122.820 ;
        RECT 37.055 114.780 37.225 122.820 ;
        RECT 39.345 114.780 39.515 122.820 ;
        RECT 34.995 114.395 36.995 114.565 ;
        RECT 37.285 114.395 39.285 114.565 ;
        RECT 40.015 113.875 40.185 123.725 ;
        RECT 40.915 123.035 42.915 123.205 ;
        RECT 43.205 123.035 45.205 123.205 ;
        RECT 40.685 114.780 40.855 122.820 ;
        RECT 42.975 114.780 43.145 122.820 ;
        RECT 45.265 114.780 45.435 122.820 ;
        RECT 40.915 114.395 42.915 114.565 ;
        RECT 43.205 114.395 45.205 114.565 ;
        RECT 45.935 113.875 46.105 123.725 ;
        RECT 46.835 123.035 48.835 123.205 ;
        RECT 49.125 123.035 51.125 123.205 ;
        RECT 46.605 114.780 46.775 122.820 ;
        RECT 48.895 114.780 49.065 122.820 ;
        RECT 51.185 114.780 51.355 122.820 ;
        RECT 46.835 114.395 48.835 114.565 ;
        RECT 49.125 114.395 51.125 114.565 ;
        RECT 51.855 113.875 52.025 123.725 ;
        RECT 52.755 123.035 54.755 123.205 ;
        RECT 55.045 123.035 57.045 123.205 ;
        RECT 52.525 114.780 52.695 122.820 ;
        RECT 54.815 114.780 54.985 122.820 ;
        RECT 57.105 114.780 57.275 122.820 ;
        RECT 52.755 114.395 54.755 114.565 ;
        RECT 55.045 114.395 57.045 114.565 ;
        RECT 57.775 113.875 57.945 123.725 ;
        RECT 58.675 123.035 60.675 123.205 ;
        RECT 60.965 123.035 62.965 123.205 ;
        RECT 58.445 114.780 58.615 122.820 ;
        RECT 60.735 114.780 60.905 122.820 ;
        RECT 63.025 114.780 63.195 122.820 ;
        RECT 58.675 114.395 60.675 114.565 ;
        RECT 60.965 114.395 62.965 114.565 ;
        RECT 63.695 113.875 63.865 123.725 ;
        RECT 64.595 123.035 66.595 123.205 ;
        RECT 66.885 123.035 68.885 123.205 ;
        RECT 64.365 114.780 64.535 122.820 ;
        RECT 66.655 114.780 66.825 122.820 ;
        RECT 68.945 114.780 69.115 122.820 ;
        RECT 64.595 114.395 66.595 114.565 ;
        RECT 66.885 114.395 68.885 114.565 ;
        RECT 69.615 113.875 70.145 123.725 ;
        RECT 10.055 113.705 70.145 113.875 ;
        RECT 10.055 103.855 10.585 113.705 ;
        RECT 11.315 113.015 13.315 113.185 ;
        RECT 13.605 113.015 15.605 113.185 ;
        RECT 11.085 104.760 11.255 112.800 ;
        RECT 13.375 104.760 13.545 112.800 ;
        RECT 15.665 104.760 15.835 112.800 ;
        RECT 11.315 104.375 13.315 104.545 ;
        RECT 13.605 104.375 15.605 104.545 ;
        RECT 16.335 103.855 16.505 113.705 ;
        RECT 17.235 113.015 19.235 113.185 ;
        RECT 19.525 113.015 21.525 113.185 ;
        RECT 17.005 104.760 17.175 112.800 ;
        RECT 19.295 104.760 19.465 112.800 ;
        RECT 21.585 104.760 21.755 112.800 ;
        RECT 17.235 104.375 19.235 104.545 ;
        RECT 19.525 104.375 21.525 104.545 ;
        RECT 22.255 103.855 22.425 113.705 ;
        RECT 23.155 113.015 25.155 113.185 ;
        RECT 25.445 113.015 27.445 113.185 ;
        RECT 22.925 104.760 23.095 112.800 ;
        RECT 25.215 104.760 25.385 112.800 ;
        RECT 27.505 104.760 27.675 112.800 ;
        RECT 23.155 104.375 25.155 104.545 ;
        RECT 25.445 104.375 27.445 104.545 ;
        RECT 28.175 103.855 28.345 113.705 ;
        RECT 29.075 113.015 31.075 113.185 ;
        RECT 31.365 113.015 33.365 113.185 ;
        RECT 28.845 104.760 29.015 112.800 ;
        RECT 31.135 104.760 31.305 112.800 ;
        RECT 33.425 104.760 33.595 112.800 ;
        RECT 29.075 104.375 31.075 104.545 ;
        RECT 31.365 104.375 33.365 104.545 ;
        RECT 34.095 103.855 34.265 113.705 ;
        RECT 34.995 113.015 36.995 113.185 ;
        RECT 37.285 113.015 39.285 113.185 ;
        RECT 34.765 104.760 34.935 112.800 ;
        RECT 37.055 104.760 37.225 112.800 ;
        RECT 39.345 104.760 39.515 112.800 ;
        RECT 34.995 104.375 36.995 104.545 ;
        RECT 37.285 104.375 39.285 104.545 ;
        RECT 40.015 103.855 40.185 113.705 ;
        RECT 40.915 113.015 42.915 113.185 ;
        RECT 43.205 113.015 45.205 113.185 ;
        RECT 40.685 104.760 40.855 112.800 ;
        RECT 42.975 104.760 43.145 112.800 ;
        RECT 45.265 104.760 45.435 112.800 ;
        RECT 40.915 104.375 42.915 104.545 ;
        RECT 43.205 104.375 45.205 104.545 ;
        RECT 45.935 103.855 46.105 113.705 ;
        RECT 46.835 113.015 48.835 113.185 ;
        RECT 49.125 113.015 51.125 113.185 ;
        RECT 46.605 104.760 46.775 112.800 ;
        RECT 48.895 104.760 49.065 112.800 ;
        RECT 51.185 104.760 51.355 112.800 ;
        RECT 46.835 104.375 48.835 104.545 ;
        RECT 49.125 104.375 51.125 104.545 ;
        RECT 51.855 103.855 52.025 113.705 ;
        RECT 52.755 113.015 54.755 113.185 ;
        RECT 55.045 113.015 57.045 113.185 ;
        RECT 52.525 104.760 52.695 112.800 ;
        RECT 54.815 104.760 54.985 112.800 ;
        RECT 57.105 104.760 57.275 112.800 ;
        RECT 52.755 104.375 54.755 104.545 ;
        RECT 55.045 104.375 57.045 104.545 ;
        RECT 57.775 103.855 57.945 113.705 ;
        RECT 58.675 113.015 60.675 113.185 ;
        RECT 60.965 113.015 62.965 113.185 ;
        RECT 58.445 104.760 58.615 112.800 ;
        RECT 60.735 104.760 60.905 112.800 ;
        RECT 63.025 104.760 63.195 112.800 ;
        RECT 58.675 104.375 60.675 104.545 ;
        RECT 60.965 104.375 62.965 104.545 ;
        RECT 63.695 103.855 63.865 113.705 ;
        RECT 64.595 113.015 66.595 113.185 ;
        RECT 66.885 113.015 68.885 113.185 ;
        RECT 64.365 104.760 64.535 112.800 ;
        RECT 66.655 104.760 66.825 112.800 ;
        RECT 68.945 104.760 69.115 112.800 ;
        RECT 64.595 104.375 66.595 104.545 ;
        RECT 66.885 104.375 68.885 104.545 ;
        RECT 69.615 103.855 70.145 113.705 ;
        RECT 10.055 103.325 70.145 103.855 ;
        RECT 71.805 123.725 114.135 124.255 ;
        RECT 138.110 124.120 145.930 124.650 ;
        RECT 71.805 113.875 72.335 123.725 ;
        RECT 72.835 122.820 77.585 123.725 ;
        RECT 72.835 114.780 73.005 122.820 ;
        RECT 75.125 114.780 75.295 122.820 ;
        RECT 77.415 114.780 77.585 122.820 ;
        RECT 73.065 114.395 75.065 114.565 ;
        RECT 75.355 114.395 77.355 114.565 ;
        RECT 78.085 113.875 78.255 123.725 ;
        RECT 78.985 123.035 80.985 123.205 ;
        RECT 81.275 123.035 83.275 123.205 ;
        RECT 78.755 114.780 78.925 122.820 ;
        RECT 81.045 114.780 81.215 122.820 ;
        RECT 83.335 114.780 83.505 122.820 ;
        RECT 78.985 114.395 80.985 114.565 ;
        RECT 81.275 114.395 83.275 114.565 ;
        RECT 84.005 113.875 84.175 123.725 ;
        RECT 84.905 123.035 86.905 123.205 ;
        RECT 87.195 123.035 89.195 123.205 ;
        RECT 84.675 114.780 84.845 122.820 ;
        RECT 86.965 114.780 87.135 122.820 ;
        RECT 89.255 114.780 89.425 122.820 ;
        RECT 84.905 114.395 86.905 114.565 ;
        RECT 87.195 114.395 89.195 114.565 ;
        RECT 89.925 113.875 90.095 123.725 ;
        RECT 90.825 123.035 92.825 123.205 ;
        RECT 93.115 123.035 95.115 123.205 ;
        RECT 90.595 114.780 90.765 122.820 ;
        RECT 92.885 114.780 93.055 122.820 ;
        RECT 95.175 114.780 95.345 122.820 ;
        RECT 90.825 114.395 92.825 114.565 ;
        RECT 93.115 114.395 95.115 114.565 ;
        RECT 95.845 113.875 96.015 123.725 ;
        RECT 96.745 123.035 98.745 123.205 ;
        RECT 99.035 123.035 101.035 123.205 ;
        RECT 96.515 114.780 96.685 122.820 ;
        RECT 98.805 114.780 98.975 122.820 ;
        RECT 101.095 114.780 101.265 122.820 ;
        RECT 96.745 114.395 98.745 114.565 ;
        RECT 99.035 114.395 101.035 114.565 ;
        RECT 101.765 113.875 101.935 123.725 ;
        RECT 102.665 123.035 104.665 123.205 ;
        RECT 104.955 123.035 106.955 123.205 ;
        RECT 102.435 114.780 102.605 122.820 ;
        RECT 104.725 114.780 104.895 122.820 ;
        RECT 107.015 114.780 107.185 122.820 ;
        RECT 102.665 114.395 104.665 114.565 ;
        RECT 104.955 114.395 106.955 114.565 ;
        RECT 107.685 113.875 107.855 123.725 ;
        RECT 108.355 122.820 113.105 123.725 ;
        RECT 108.355 114.780 108.525 122.820 ;
        RECT 110.645 114.780 110.815 122.820 ;
        RECT 112.935 114.780 113.105 122.820 ;
        RECT 108.585 114.395 110.585 114.565 ;
        RECT 110.875 114.395 112.875 114.565 ;
        RECT 113.605 113.875 114.135 123.725 ;
        RECT 71.805 113.705 114.135 113.875 ;
        RECT 71.805 103.855 72.335 113.705 ;
        RECT 73.065 113.015 75.065 113.185 ;
        RECT 75.355 113.015 77.355 113.185 ;
        RECT 72.835 104.760 73.005 112.800 ;
        RECT 75.125 104.760 75.295 112.800 ;
        RECT 77.415 104.760 77.585 112.800 ;
        RECT 72.835 103.855 77.585 104.760 ;
        RECT 78.085 103.855 78.255 113.705 ;
        RECT 78.985 113.015 80.985 113.185 ;
        RECT 81.275 113.015 83.275 113.185 ;
        RECT 78.755 104.760 78.925 112.800 ;
        RECT 81.045 104.760 81.215 112.800 ;
        RECT 83.335 104.760 83.505 112.800 ;
        RECT 78.985 104.375 80.985 104.545 ;
        RECT 81.275 104.375 83.275 104.545 ;
        RECT 84.005 103.855 84.175 113.705 ;
        RECT 84.905 113.015 86.905 113.185 ;
        RECT 87.195 113.015 89.195 113.185 ;
        RECT 84.675 104.760 84.845 112.800 ;
        RECT 86.965 104.760 87.135 112.800 ;
        RECT 89.255 104.760 89.425 112.800 ;
        RECT 84.905 104.375 86.905 104.545 ;
        RECT 87.195 104.375 89.195 104.545 ;
        RECT 89.925 103.855 90.095 113.705 ;
        RECT 90.825 113.015 92.825 113.185 ;
        RECT 93.115 113.015 95.115 113.185 ;
        RECT 90.595 104.760 90.765 112.800 ;
        RECT 92.885 104.760 93.055 112.800 ;
        RECT 95.175 104.760 95.345 112.800 ;
        RECT 90.825 104.375 92.825 104.545 ;
        RECT 93.115 104.375 95.115 104.545 ;
        RECT 95.845 103.855 96.015 113.705 ;
        RECT 96.745 113.015 98.745 113.185 ;
        RECT 99.035 113.015 101.035 113.185 ;
        RECT 96.515 104.760 96.685 112.800 ;
        RECT 98.805 104.760 98.975 112.800 ;
        RECT 101.095 104.760 101.265 112.800 ;
        RECT 96.745 104.375 98.745 104.545 ;
        RECT 99.035 104.375 101.035 104.545 ;
        RECT 101.765 103.855 101.935 113.705 ;
        RECT 102.665 113.015 104.665 113.185 ;
        RECT 104.955 113.015 106.955 113.185 ;
        RECT 102.435 104.760 102.605 112.800 ;
        RECT 104.725 104.760 104.895 112.800 ;
        RECT 107.015 104.760 107.185 112.800 ;
        RECT 102.665 104.375 104.665 104.545 ;
        RECT 104.955 104.375 106.955 104.545 ;
        RECT 107.685 103.855 107.855 113.705 ;
        RECT 108.585 113.015 110.585 113.185 ;
        RECT 110.875 113.015 112.875 113.185 ;
        RECT 108.355 104.760 108.525 112.800 ;
        RECT 110.645 104.760 110.815 112.800 ;
        RECT 112.935 104.760 113.105 112.800 ;
        RECT 108.355 103.855 113.105 104.760 ;
        RECT 113.605 103.855 114.135 113.705 ;
        RECT 71.805 103.325 114.135 103.855 ;
        RECT 115.935 122.945 128.905 123.475 ;
        RECT 115.935 113.485 116.465 122.945 ;
        RECT 117.370 122.275 118.410 122.445 ;
        RECT 116.985 114.215 117.155 122.215 ;
        RECT 118.625 114.215 118.795 122.215 ;
        RECT 117.370 113.985 118.410 114.155 ;
        RECT 119.315 113.485 119.485 122.945 ;
        RECT 120.390 122.275 121.430 122.445 ;
        RECT 120.005 114.215 120.175 122.215 ;
        RECT 121.645 114.215 121.815 122.215 ;
        RECT 120.390 113.985 121.430 114.155 ;
        RECT 122.335 113.485 122.505 122.945 ;
        RECT 123.410 122.275 124.450 122.445 ;
        RECT 123.025 114.215 123.195 122.215 ;
        RECT 124.665 114.215 124.835 122.215 ;
        RECT 123.410 113.985 124.450 114.155 ;
        RECT 125.355 113.485 125.525 122.945 ;
        RECT 126.430 122.275 127.470 122.445 ;
        RECT 126.045 114.215 126.215 122.215 ;
        RECT 127.685 114.215 127.855 122.215 ;
        RECT 126.430 113.985 127.470 114.155 ;
        RECT 128.375 113.485 128.905 122.945 ;
        RECT 115.935 113.315 128.905 113.485 ;
        RECT 115.935 103.855 116.465 113.315 ;
        RECT 117.370 112.645 118.410 112.815 ;
        RECT 116.985 104.585 117.155 112.585 ;
        RECT 118.625 104.585 118.795 112.585 ;
        RECT 117.370 104.355 118.410 104.525 ;
        RECT 119.315 103.855 119.485 113.315 ;
        RECT 120.390 112.645 121.430 112.815 ;
        RECT 120.005 104.585 120.175 112.585 ;
        RECT 121.645 104.585 121.815 112.585 ;
        RECT 120.390 104.355 121.430 104.525 ;
        RECT 122.335 103.855 122.505 113.315 ;
        RECT 123.410 112.645 124.450 112.815 ;
        RECT 123.025 104.585 123.195 112.585 ;
        RECT 124.665 104.585 124.835 112.585 ;
        RECT 123.410 104.355 124.450 104.525 ;
        RECT 125.355 103.855 125.525 113.315 ;
        RECT 126.430 112.645 127.470 112.815 ;
        RECT 126.045 104.585 126.215 112.585 ;
        RECT 127.685 104.585 127.855 112.585 ;
        RECT 126.430 104.355 127.470 104.525 ;
        RECT 128.375 103.855 128.905 113.315 ;
        RECT 115.935 103.325 128.905 103.855 ;
        RECT 135.150 104.785 149.540 108.660 ;
        RECT 10.055 102.145 128.905 102.675 ;
        RECT 10.055 92.295 10.585 102.145 ;
        RECT 11.315 101.455 13.315 101.625 ;
        RECT 13.605 101.455 15.605 101.625 ;
        RECT 15.895 101.455 17.895 101.625 ;
        RECT 18.185 101.455 20.185 101.625 ;
        RECT 20.475 101.455 22.475 101.625 ;
        RECT 22.765 101.455 24.765 101.625 ;
        RECT 25.055 101.455 27.055 101.625 ;
        RECT 27.345 101.455 29.345 101.625 ;
        RECT 11.085 93.200 11.255 101.240 ;
        RECT 13.375 93.200 13.545 101.240 ;
        RECT 15.665 93.200 15.835 101.240 ;
        RECT 17.955 93.200 18.125 101.240 ;
        RECT 20.245 93.200 20.415 101.240 ;
        RECT 22.535 93.200 22.705 101.240 ;
        RECT 24.825 93.200 24.995 101.240 ;
        RECT 27.115 93.200 27.285 101.240 ;
        RECT 29.405 93.200 29.575 101.240 ;
        RECT 11.315 92.815 13.315 92.985 ;
        RECT 13.605 92.815 15.605 92.985 ;
        RECT 15.895 92.815 17.895 92.985 ;
        RECT 18.185 92.815 20.185 92.985 ;
        RECT 20.475 92.815 22.475 92.985 ;
        RECT 22.765 92.815 24.765 92.985 ;
        RECT 25.055 92.815 27.055 92.985 ;
        RECT 27.345 92.815 29.345 92.985 ;
        RECT 30.075 92.295 30.245 102.145 ;
        RECT 30.975 101.455 32.975 101.625 ;
        RECT 33.265 101.455 35.265 101.625 ;
        RECT 35.555 101.455 37.555 101.625 ;
        RECT 37.845 101.455 39.845 101.625 ;
        RECT 40.135 101.455 42.135 101.625 ;
        RECT 42.425 101.455 44.425 101.625 ;
        RECT 44.715 101.455 46.715 101.625 ;
        RECT 47.005 101.455 49.005 101.625 ;
        RECT 30.745 93.200 30.915 101.240 ;
        RECT 33.035 93.200 33.205 101.240 ;
        RECT 35.325 93.200 35.495 101.240 ;
        RECT 37.615 93.200 37.785 101.240 ;
        RECT 39.905 93.200 40.075 101.240 ;
        RECT 42.195 93.200 42.365 101.240 ;
        RECT 44.485 93.200 44.655 101.240 ;
        RECT 46.775 93.200 46.945 101.240 ;
        RECT 49.065 93.200 49.235 101.240 ;
        RECT 30.975 92.815 32.975 92.985 ;
        RECT 33.265 92.815 35.265 92.985 ;
        RECT 35.555 92.815 37.555 92.985 ;
        RECT 37.845 92.815 39.845 92.985 ;
        RECT 40.135 92.815 42.135 92.985 ;
        RECT 42.425 92.815 44.425 92.985 ;
        RECT 44.715 92.815 46.715 92.985 ;
        RECT 47.005 92.815 49.005 92.985 ;
        RECT 49.735 92.295 49.905 102.145 ;
        RECT 50.635 101.455 52.635 101.625 ;
        RECT 52.925 101.455 54.925 101.625 ;
        RECT 55.215 101.455 57.215 101.625 ;
        RECT 57.505 101.455 59.505 101.625 ;
        RECT 59.795 101.455 61.795 101.625 ;
        RECT 62.085 101.455 64.085 101.625 ;
        RECT 64.375 101.455 66.375 101.625 ;
        RECT 66.665 101.455 68.665 101.625 ;
        RECT 50.405 93.200 50.575 101.240 ;
        RECT 52.695 93.200 52.865 101.240 ;
        RECT 54.985 93.200 55.155 101.240 ;
        RECT 57.275 93.200 57.445 101.240 ;
        RECT 59.565 93.200 59.735 101.240 ;
        RECT 61.855 93.200 62.025 101.240 ;
        RECT 64.145 93.200 64.315 101.240 ;
        RECT 66.435 93.200 66.605 101.240 ;
        RECT 68.725 93.200 68.895 101.240 ;
        RECT 50.635 92.815 52.635 92.985 ;
        RECT 52.925 92.815 54.925 92.985 ;
        RECT 55.215 92.815 57.215 92.985 ;
        RECT 57.505 92.815 59.505 92.985 ;
        RECT 59.795 92.815 61.795 92.985 ;
        RECT 62.085 92.815 64.085 92.985 ;
        RECT 64.375 92.815 66.375 92.985 ;
        RECT 66.665 92.815 68.665 92.985 ;
        RECT 69.395 92.295 69.565 102.145 ;
        RECT 70.295 101.455 72.295 101.625 ;
        RECT 72.585 101.455 74.585 101.625 ;
        RECT 74.875 101.455 76.875 101.625 ;
        RECT 77.165 101.455 79.165 101.625 ;
        RECT 79.455 101.455 81.455 101.625 ;
        RECT 81.745 101.455 83.745 101.625 ;
        RECT 84.035 101.455 86.035 101.625 ;
        RECT 86.325 101.455 88.325 101.625 ;
        RECT 70.065 93.200 70.235 101.240 ;
        RECT 72.355 93.200 72.525 101.240 ;
        RECT 74.645 93.200 74.815 101.240 ;
        RECT 76.935 93.200 77.105 101.240 ;
        RECT 79.225 93.200 79.395 101.240 ;
        RECT 81.515 93.200 81.685 101.240 ;
        RECT 83.805 93.200 83.975 101.240 ;
        RECT 86.095 93.200 86.265 101.240 ;
        RECT 88.385 93.200 88.555 101.240 ;
        RECT 70.295 92.815 72.295 92.985 ;
        RECT 72.585 92.815 74.585 92.985 ;
        RECT 74.875 92.815 76.875 92.985 ;
        RECT 77.165 92.815 79.165 92.985 ;
        RECT 79.455 92.815 81.455 92.985 ;
        RECT 81.745 92.815 83.745 92.985 ;
        RECT 84.035 92.815 86.035 92.985 ;
        RECT 86.325 92.815 88.325 92.985 ;
        RECT 89.055 92.295 89.225 102.145 ;
        RECT 89.955 101.455 91.955 101.625 ;
        RECT 92.245 101.455 94.245 101.625 ;
        RECT 94.535 101.455 96.535 101.625 ;
        RECT 96.825 101.455 98.825 101.625 ;
        RECT 99.115 101.455 101.115 101.625 ;
        RECT 101.405 101.455 103.405 101.625 ;
        RECT 103.695 101.455 105.695 101.625 ;
        RECT 105.985 101.455 107.985 101.625 ;
        RECT 89.725 93.200 89.895 101.240 ;
        RECT 92.015 93.200 92.185 101.240 ;
        RECT 94.305 93.200 94.475 101.240 ;
        RECT 96.595 93.200 96.765 101.240 ;
        RECT 98.885 93.200 99.055 101.240 ;
        RECT 101.175 93.200 101.345 101.240 ;
        RECT 103.465 93.200 103.635 101.240 ;
        RECT 105.755 93.200 105.925 101.240 ;
        RECT 108.045 93.200 108.215 101.240 ;
        RECT 89.955 92.815 91.955 92.985 ;
        RECT 92.245 92.815 94.245 92.985 ;
        RECT 94.535 92.815 96.535 92.985 ;
        RECT 96.825 92.815 98.825 92.985 ;
        RECT 99.115 92.815 101.115 92.985 ;
        RECT 101.405 92.815 103.405 92.985 ;
        RECT 103.695 92.815 105.695 92.985 ;
        RECT 105.985 92.815 107.985 92.985 ;
        RECT 108.715 92.295 108.885 102.145 ;
        RECT 109.615 101.455 111.615 101.625 ;
        RECT 111.905 101.455 113.905 101.625 ;
        RECT 114.195 101.455 116.195 101.625 ;
        RECT 116.485 101.455 118.485 101.625 ;
        RECT 118.775 101.455 120.775 101.625 ;
        RECT 121.065 101.455 123.065 101.625 ;
        RECT 123.355 101.455 125.355 101.625 ;
        RECT 125.645 101.455 127.645 101.625 ;
        RECT 109.385 93.200 109.555 101.240 ;
        RECT 111.675 93.200 111.845 101.240 ;
        RECT 113.965 93.200 114.135 101.240 ;
        RECT 116.255 93.200 116.425 101.240 ;
        RECT 118.545 93.200 118.715 101.240 ;
        RECT 120.835 93.200 121.005 101.240 ;
        RECT 123.125 93.200 123.295 101.240 ;
        RECT 125.415 93.200 125.585 101.240 ;
        RECT 127.705 93.200 127.875 101.240 ;
        RECT 109.615 92.815 111.615 92.985 ;
        RECT 111.905 92.815 113.905 92.985 ;
        RECT 114.195 92.815 116.195 92.985 ;
        RECT 116.485 92.815 118.485 92.985 ;
        RECT 118.775 92.815 120.775 92.985 ;
        RECT 121.065 92.815 123.065 92.985 ;
        RECT 123.355 92.815 125.355 92.985 ;
        RECT 125.645 92.815 127.645 92.985 ;
        RECT 128.375 92.295 128.905 102.145 ;
        RECT 10.055 92.125 128.905 92.295 ;
        RECT 10.055 82.275 10.585 92.125 ;
        RECT 11.315 91.435 13.315 91.605 ;
        RECT 13.605 91.435 15.605 91.605 ;
        RECT 15.895 91.435 17.895 91.605 ;
        RECT 18.185 91.435 20.185 91.605 ;
        RECT 20.475 91.435 22.475 91.605 ;
        RECT 22.765 91.435 24.765 91.605 ;
        RECT 25.055 91.435 27.055 91.605 ;
        RECT 27.345 91.435 29.345 91.605 ;
        RECT 11.085 83.180 11.255 91.220 ;
        RECT 13.375 83.180 13.545 91.220 ;
        RECT 15.665 83.180 15.835 91.220 ;
        RECT 17.955 83.180 18.125 91.220 ;
        RECT 20.245 83.180 20.415 91.220 ;
        RECT 22.535 83.180 22.705 91.220 ;
        RECT 24.825 83.180 24.995 91.220 ;
        RECT 27.115 83.180 27.285 91.220 ;
        RECT 29.405 83.180 29.575 91.220 ;
        RECT 11.315 82.795 13.315 82.965 ;
        RECT 13.605 82.795 15.605 82.965 ;
        RECT 15.895 82.795 17.895 82.965 ;
        RECT 18.185 82.795 20.185 82.965 ;
        RECT 20.475 82.795 22.475 82.965 ;
        RECT 22.765 82.795 24.765 82.965 ;
        RECT 25.055 82.795 27.055 82.965 ;
        RECT 27.345 82.795 29.345 82.965 ;
        RECT 30.075 82.275 30.245 92.125 ;
        RECT 30.975 91.435 32.975 91.605 ;
        RECT 33.265 91.435 35.265 91.605 ;
        RECT 35.555 91.435 37.555 91.605 ;
        RECT 37.845 91.435 39.845 91.605 ;
        RECT 40.135 91.435 42.135 91.605 ;
        RECT 42.425 91.435 44.425 91.605 ;
        RECT 44.715 91.435 46.715 91.605 ;
        RECT 47.005 91.435 49.005 91.605 ;
        RECT 30.745 83.180 30.915 91.220 ;
        RECT 33.035 83.180 33.205 91.220 ;
        RECT 35.325 83.180 35.495 91.220 ;
        RECT 37.615 83.180 37.785 91.220 ;
        RECT 39.905 83.180 40.075 91.220 ;
        RECT 42.195 83.180 42.365 91.220 ;
        RECT 44.485 83.180 44.655 91.220 ;
        RECT 46.775 83.180 46.945 91.220 ;
        RECT 49.065 83.180 49.235 91.220 ;
        RECT 30.975 82.795 32.975 82.965 ;
        RECT 33.265 82.795 35.265 82.965 ;
        RECT 35.555 82.795 37.555 82.965 ;
        RECT 37.845 82.795 39.845 82.965 ;
        RECT 40.135 82.795 42.135 82.965 ;
        RECT 42.425 82.795 44.425 82.965 ;
        RECT 44.715 82.795 46.715 82.965 ;
        RECT 47.005 82.795 49.005 82.965 ;
        RECT 49.735 82.275 49.905 92.125 ;
        RECT 50.635 91.435 52.635 91.605 ;
        RECT 52.925 91.435 54.925 91.605 ;
        RECT 55.215 91.435 57.215 91.605 ;
        RECT 57.505 91.435 59.505 91.605 ;
        RECT 59.795 91.435 61.795 91.605 ;
        RECT 62.085 91.435 64.085 91.605 ;
        RECT 64.375 91.435 66.375 91.605 ;
        RECT 66.665 91.435 68.665 91.605 ;
        RECT 50.405 83.180 50.575 91.220 ;
        RECT 52.695 83.180 52.865 91.220 ;
        RECT 54.985 83.180 55.155 91.220 ;
        RECT 57.275 83.180 57.445 91.220 ;
        RECT 59.565 83.180 59.735 91.220 ;
        RECT 61.855 83.180 62.025 91.220 ;
        RECT 64.145 83.180 64.315 91.220 ;
        RECT 66.435 83.180 66.605 91.220 ;
        RECT 68.725 83.180 68.895 91.220 ;
        RECT 50.635 82.795 52.635 82.965 ;
        RECT 52.925 82.795 54.925 82.965 ;
        RECT 55.215 82.795 57.215 82.965 ;
        RECT 57.505 82.795 59.505 82.965 ;
        RECT 59.795 82.795 61.795 82.965 ;
        RECT 62.085 82.795 64.085 82.965 ;
        RECT 64.375 82.795 66.375 82.965 ;
        RECT 66.665 82.795 68.665 82.965 ;
        RECT 69.395 82.275 69.565 92.125 ;
        RECT 70.295 91.435 72.295 91.605 ;
        RECT 72.585 91.435 74.585 91.605 ;
        RECT 74.875 91.435 76.875 91.605 ;
        RECT 77.165 91.435 79.165 91.605 ;
        RECT 79.455 91.435 81.455 91.605 ;
        RECT 81.745 91.435 83.745 91.605 ;
        RECT 84.035 91.435 86.035 91.605 ;
        RECT 86.325 91.435 88.325 91.605 ;
        RECT 70.065 83.180 70.235 91.220 ;
        RECT 72.355 83.180 72.525 91.220 ;
        RECT 74.645 83.180 74.815 91.220 ;
        RECT 76.935 83.180 77.105 91.220 ;
        RECT 79.225 83.180 79.395 91.220 ;
        RECT 81.515 83.180 81.685 91.220 ;
        RECT 83.805 83.180 83.975 91.220 ;
        RECT 86.095 83.180 86.265 91.220 ;
        RECT 88.385 83.180 88.555 91.220 ;
        RECT 70.295 82.795 72.295 82.965 ;
        RECT 72.585 82.795 74.585 82.965 ;
        RECT 74.875 82.795 76.875 82.965 ;
        RECT 77.165 82.795 79.165 82.965 ;
        RECT 79.455 82.795 81.455 82.965 ;
        RECT 81.745 82.795 83.745 82.965 ;
        RECT 84.035 82.795 86.035 82.965 ;
        RECT 86.325 82.795 88.325 82.965 ;
        RECT 89.055 82.275 89.225 92.125 ;
        RECT 89.955 91.435 91.955 91.605 ;
        RECT 92.245 91.435 94.245 91.605 ;
        RECT 94.535 91.435 96.535 91.605 ;
        RECT 96.825 91.435 98.825 91.605 ;
        RECT 99.115 91.435 101.115 91.605 ;
        RECT 101.405 91.435 103.405 91.605 ;
        RECT 103.695 91.435 105.695 91.605 ;
        RECT 105.985 91.435 107.985 91.605 ;
        RECT 89.725 83.180 89.895 91.220 ;
        RECT 92.015 83.180 92.185 91.220 ;
        RECT 94.305 83.180 94.475 91.220 ;
        RECT 96.595 83.180 96.765 91.220 ;
        RECT 98.885 83.180 99.055 91.220 ;
        RECT 101.175 83.180 101.345 91.220 ;
        RECT 103.465 83.180 103.635 91.220 ;
        RECT 105.755 83.180 105.925 91.220 ;
        RECT 108.045 83.180 108.215 91.220 ;
        RECT 89.955 82.795 91.955 82.965 ;
        RECT 92.245 82.795 94.245 82.965 ;
        RECT 94.535 82.795 96.535 82.965 ;
        RECT 96.825 82.795 98.825 82.965 ;
        RECT 99.115 82.795 101.115 82.965 ;
        RECT 101.405 82.795 103.405 82.965 ;
        RECT 103.695 82.795 105.695 82.965 ;
        RECT 105.985 82.795 107.985 82.965 ;
        RECT 108.715 82.275 108.885 92.125 ;
        RECT 109.615 91.435 111.615 91.605 ;
        RECT 111.905 91.435 113.905 91.605 ;
        RECT 114.195 91.435 116.195 91.605 ;
        RECT 116.485 91.435 118.485 91.605 ;
        RECT 118.775 91.435 120.775 91.605 ;
        RECT 121.065 91.435 123.065 91.605 ;
        RECT 123.355 91.435 125.355 91.605 ;
        RECT 125.645 91.435 127.645 91.605 ;
        RECT 109.385 83.180 109.555 91.220 ;
        RECT 111.675 83.180 111.845 91.220 ;
        RECT 113.965 83.180 114.135 91.220 ;
        RECT 116.255 83.180 116.425 91.220 ;
        RECT 118.545 83.180 118.715 91.220 ;
        RECT 120.835 83.180 121.005 91.220 ;
        RECT 123.125 83.180 123.295 91.220 ;
        RECT 125.415 83.180 125.585 91.220 ;
        RECT 127.705 83.180 127.875 91.220 ;
        RECT 109.615 82.795 111.615 82.965 ;
        RECT 111.905 82.795 113.905 82.965 ;
        RECT 114.195 82.795 116.195 82.965 ;
        RECT 116.485 82.795 118.485 82.965 ;
        RECT 118.775 82.795 120.775 82.965 ;
        RECT 121.065 82.795 123.065 82.965 ;
        RECT 123.355 82.795 125.355 82.965 ;
        RECT 125.645 82.795 127.645 82.965 ;
        RECT 128.375 82.275 128.905 92.125 ;
        RECT 10.055 82.105 128.905 82.275 ;
        RECT 10.055 72.255 10.585 82.105 ;
        RECT 11.315 81.415 13.315 81.585 ;
        RECT 13.605 81.415 15.605 81.585 ;
        RECT 15.895 81.415 17.895 81.585 ;
        RECT 18.185 81.415 20.185 81.585 ;
        RECT 20.475 81.415 22.475 81.585 ;
        RECT 22.765 81.415 24.765 81.585 ;
        RECT 25.055 81.415 27.055 81.585 ;
        RECT 27.345 81.415 29.345 81.585 ;
        RECT 11.085 73.160 11.255 81.200 ;
        RECT 13.375 73.160 13.545 81.200 ;
        RECT 15.665 73.160 15.835 81.200 ;
        RECT 17.955 73.160 18.125 81.200 ;
        RECT 20.245 73.160 20.415 81.200 ;
        RECT 22.535 73.160 22.705 81.200 ;
        RECT 24.825 73.160 24.995 81.200 ;
        RECT 27.115 73.160 27.285 81.200 ;
        RECT 29.405 73.160 29.575 81.200 ;
        RECT 11.315 72.775 13.315 72.945 ;
        RECT 13.605 72.775 15.605 72.945 ;
        RECT 15.895 72.775 17.895 72.945 ;
        RECT 18.185 72.775 20.185 72.945 ;
        RECT 20.475 72.775 22.475 72.945 ;
        RECT 22.765 72.775 24.765 72.945 ;
        RECT 25.055 72.775 27.055 72.945 ;
        RECT 27.345 72.775 29.345 72.945 ;
        RECT 30.075 72.255 30.245 82.105 ;
        RECT 30.975 81.415 32.975 81.585 ;
        RECT 33.265 81.415 35.265 81.585 ;
        RECT 35.555 81.415 37.555 81.585 ;
        RECT 37.845 81.415 39.845 81.585 ;
        RECT 40.135 81.415 42.135 81.585 ;
        RECT 42.425 81.415 44.425 81.585 ;
        RECT 44.715 81.415 46.715 81.585 ;
        RECT 47.005 81.415 49.005 81.585 ;
        RECT 30.745 73.160 30.915 81.200 ;
        RECT 33.035 73.160 33.205 81.200 ;
        RECT 35.325 73.160 35.495 81.200 ;
        RECT 37.615 73.160 37.785 81.200 ;
        RECT 39.905 73.160 40.075 81.200 ;
        RECT 42.195 73.160 42.365 81.200 ;
        RECT 44.485 73.160 44.655 81.200 ;
        RECT 46.775 73.160 46.945 81.200 ;
        RECT 49.065 73.160 49.235 81.200 ;
        RECT 30.975 72.775 32.975 72.945 ;
        RECT 33.265 72.775 35.265 72.945 ;
        RECT 35.555 72.775 37.555 72.945 ;
        RECT 37.845 72.775 39.845 72.945 ;
        RECT 40.135 72.775 42.135 72.945 ;
        RECT 42.425 72.775 44.425 72.945 ;
        RECT 44.715 72.775 46.715 72.945 ;
        RECT 47.005 72.775 49.005 72.945 ;
        RECT 49.735 72.255 49.905 82.105 ;
        RECT 50.635 81.415 52.635 81.585 ;
        RECT 52.925 81.415 54.925 81.585 ;
        RECT 55.215 81.415 57.215 81.585 ;
        RECT 57.505 81.415 59.505 81.585 ;
        RECT 59.795 81.415 61.795 81.585 ;
        RECT 62.085 81.415 64.085 81.585 ;
        RECT 64.375 81.415 66.375 81.585 ;
        RECT 66.665 81.415 68.665 81.585 ;
        RECT 50.405 73.160 50.575 81.200 ;
        RECT 52.695 73.160 52.865 81.200 ;
        RECT 54.985 73.160 55.155 81.200 ;
        RECT 57.275 73.160 57.445 81.200 ;
        RECT 59.565 73.160 59.735 81.200 ;
        RECT 61.855 73.160 62.025 81.200 ;
        RECT 64.145 73.160 64.315 81.200 ;
        RECT 66.435 73.160 66.605 81.200 ;
        RECT 68.725 73.160 68.895 81.200 ;
        RECT 50.635 72.775 52.635 72.945 ;
        RECT 52.925 72.775 54.925 72.945 ;
        RECT 55.215 72.775 57.215 72.945 ;
        RECT 57.505 72.775 59.505 72.945 ;
        RECT 59.795 72.775 61.795 72.945 ;
        RECT 62.085 72.775 64.085 72.945 ;
        RECT 64.375 72.775 66.375 72.945 ;
        RECT 66.665 72.775 68.665 72.945 ;
        RECT 69.395 72.255 69.565 82.105 ;
        RECT 70.295 81.415 72.295 81.585 ;
        RECT 72.585 81.415 74.585 81.585 ;
        RECT 74.875 81.415 76.875 81.585 ;
        RECT 77.165 81.415 79.165 81.585 ;
        RECT 79.455 81.415 81.455 81.585 ;
        RECT 81.745 81.415 83.745 81.585 ;
        RECT 84.035 81.415 86.035 81.585 ;
        RECT 86.325 81.415 88.325 81.585 ;
        RECT 70.065 73.160 70.235 81.200 ;
        RECT 72.355 73.160 72.525 81.200 ;
        RECT 74.645 73.160 74.815 81.200 ;
        RECT 76.935 73.160 77.105 81.200 ;
        RECT 79.225 73.160 79.395 81.200 ;
        RECT 81.515 73.160 81.685 81.200 ;
        RECT 83.805 73.160 83.975 81.200 ;
        RECT 86.095 73.160 86.265 81.200 ;
        RECT 88.385 73.160 88.555 81.200 ;
        RECT 70.295 72.775 72.295 72.945 ;
        RECT 72.585 72.775 74.585 72.945 ;
        RECT 74.875 72.775 76.875 72.945 ;
        RECT 77.165 72.775 79.165 72.945 ;
        RECT 79.455 72.775 81.455 72.945 ;
        RECT 81.745 72.775 83.745 72.945 ;
        RECT 84.035 72.775 86.035 72.945 ;
        RECT 86.325 72.775 88.325 72.945 ;
        RECT 89.055 72.255 89.225 82.105 ;
        RECT 89.955 81.415 91.955 81.585 ;
        RECT 92.245 81.415 94.245 81.585 ;
        RECT 94.535 81.415 96.535 81.585 ;
        RECT 96.825 81.415 98.825 81.585 ;
        RECT 99.115 81.415 101.115 81.585 ;
        RECT 101.405 81.415 103.405 81.585 ;
        RECT 103.695 81.415 105.695 81.585 ;
        RECT 105.985 81.415 107.985 81.585 ;
        RECT 89.725 73.160 89.895 81.200 ;
        RECT 92.015 73.160 92.185 81.200 ;
        RECT 94.305 73.160 94.475 81.200 ;
        RECT 96.595 73.160 96.765 81.200 ;
        RECT 98.885 73.160 99.055 81.200 ;
        RECT 101.175 73.160 101.345 81.200 ;
        RECT 103.465 73.160 103.635 81.200 ;
        RECT 105.755 73.160 105.925 81.200 ;
        RECT 108.045 73.160 108.215 81.200 ;
        RECT 89.955 72.775 91.955 72.945 ;
        RECT 92.245 72.775 94.245 72.945 ;
        RECT 94.535 72.775 96.535 72.945 ;
        RECT 96.825 72.775 98.825 72.945 ;
        RECT 99.115 72.775 101.115 72.945 ;
        RECT 101.405 72.775 103.405 72.945 ;
        RECT 103.695 72.775 105.695 72.945 ;
        RECT 105.985 72.775 107.985 72.945 ;
        RECT 108.715 72.255 108.885 82.105 ;
        RECT 109.615 81.415 111.615 81.585 ;
        RECT 111.905 81.415 113.905 81.585 ;
        RECT 114.195 81.415 116.195 81.585 ;
        RECT 116.485 81.415 118.485 81.585 ;
        RECT 118.775 81.415 120.775 81.585 ;
        RECT 121.065 81.415 123.065 81.585 ;
        RECT 123.355 81.415 125.355 81.585 ;
        RECT 125.645 81.415 127.645 81.585 ;
        RECT 109.385 73.160 109.555 81.200 ;
        RECT 111.675 73.160 111.845 81.200 ;
        RECT 113.965 73.160 114.135 81.200 ;
        RECT 116.255 73.160 116.425 81.200 ;
        RECT 118.545 73.160 118.715 81.200 ;
        RECT 120.835 73.160 121.005 81.200 ;
        RECT 123.125 73.160 123.295 81.200 ;
        RECT 125.415 73.160 125.585 81.200 ;
        RECT 127.705 73.160 127.875 81.200 ;
        RECT 109.615 72.775 111.615 72.945 ;
        RECT 111.905 72.775 113.905 72.945 ;
        RECT 114.195 72.775 116.195 72.945 ;
        RECT 116.485 72.775 118.485 72.945 ;
        RECT 118.775 72.775 120.775 72.945 ;
        RECT 121.065 72.775 123.065 72.945 ;
        RECT 123.355 72.775 125.355 72.945 ;
        RECT 125.645 72.775 127.645 72.945 ;
        RECT 128.375 72.255 128.905 82.105 ;
        RECT 10.055 72.085 128.905 72.255 ;
        RECT 10.055 62.235 10.585 72.085 ;
        RECT 11.315 71.395 13.315 71.565 ;
        RECT 13.605 71.395 15.605 71.565 ;
        RECT 15.895 71.395 17.895 71.565 ;
        RECT 18.185 71.395 20.185 71.565 ;
        RECT 20.475 71.395 22.475 71.565 ;
        RECT 22.765 71.395 24.765 71.565 ;
        RECT 25.055 71.395 27.055 71.565 ;
        RECT 27.345 71.395 29.345 71.565 ;
        RECT 11.085 63.140 11.255 71.180 ;
        RECT 13.375 63.140 13.545 71.180 ;
        RECT 15.665 63.140 15.835 71.180 ;
        RECT 17.955 63.140 18.125 71.180 ;
        RECT 20.245 63.140 20.415 71.180 ;
        RECT 22.535 63.140 22.705 71.180 ;
        RECT 24.825 63.140 24.995 71.180 ;
        RECT 27.115 63.140 27.285 71.180 ;
        RECT 29.405 63.140 29.575 71.180 ;
        RECT 11.315 62.755 13.315 62.925 ;
        RECT 13.605 62.755 15.605 62.925 ;
        RECT 15.895 62.755 17.895 62.925 ;
        RECT 18.185 62.755 20.185 62.925 ;
        RECT 20.475 62.755 22.475 62.925 ;
        RECT 22.765 62.755 24.765 62.925 ;
        RECT 25.055 62.755 27.055 62.925 ;
        RECT 27.345 62.755 29.345 62.925 ;
        RECT 30.075 62.235 30.245 72.085 ;
        RECT 30.975 71.395 32.975 71.565 ;
        RECT 33.265 71.395 35.265 71.565 ;
        RECT 35.555 71.395 37.555 71.565 ;
        RECT 37.845 71.395 39.845 71.565 ;
        RECT 40.135 71.395 42.135 71.565 ;
        RECT 42.425 71.395 44.425 71.565 ;
        RECT 44.715 71.395 46.715 71.565 ;
        RECT 47.005 71.395 49.005 71.565 ;
        RECT 30.745 63.140 30.915 71.180 ;
        RECT 33.035 63.140 33.205 71.180 ;
        RECT 35.325 63.140 35.495 71.180 ;
        RECT 37.615 63.140 37.785 71.180 ;
        RECT 39.905 63.140 40.075 71.180 ;
        RECT 42.195 63.140 42.365 71.180 ;
        RECT 44.485 63.140 44.655 71.180 ;
        RECT 46.775 63.140 46.945 71.180 ;
        RECT 49.065 63.140 49.235 71.180 ;
        RECT 30.975 62.755 32.975 62.925 ;
        RECT 33.265 62.755 35.265 62.925 ;
        RECT 35.555 62.755 37.555 62.925 ;
        RECT 37.845 62.755 39.845 62.925 ;
        RECT 40.135 62.755 42.135 62.925 ;
        RECT 42.425 62.755 44.425 62.925 ;
        RECT 44.715 62.755 46.715 62.925 ;
        RECT 47.005 62.755 49.005 62.925 ;
        RECT 49.735 62.235 49.905 72.085 ;
        RECT 50.635 71.395 52.635 71.565 ;
        RECT 52.925 71.395 54.925 71.565 ;
        RECT 55.215 71.395 57.215 71.565 ;
        RECT 57.505 71.395 59.505 71.565 ;
        RECT 59.795 71.395 61.795 71.565 ;
        RECT 62.085 71.395 64.085 71.565 ;
        RECT 64.375 71.395 66.375 71.565 ;
        RECT 66.665 71.395 68.665 71.565 ;
        RECT 50.405 63.140 50.575 71.180 ;
        RECT 52.695 63.140 52.865 71.180 ;
        RECT 54.985 63.140 55.155 71.180 ;
        RECT 57.275 63.140 57.445 71.180 ;
        RECT 59.565 63.140 59.735 71.180 ;
        RECT 61.855 63.140 62.025 71.180 ;
        RECT 64.145 63.140 64.315 71.180 ;
        RECT 66.435 63.140 66.605 71.180 ;
        RECT 68.725 63.140 68.895 71.180 ;
        RECT 50.635 62.755 52.635 62.925 ;
        RECT 52.925 62.755 54.925 62.925 ;
        RECT 55.215 62.755 57.215 62.925 ;
        RECT 57.505 62.755 59.505 62.925 ;
        RECT 59.795 62.755 61.795 62.925 ;
        RECT 62.085 62.755 64.085 62.925 ;
        RECT 64.375 62.755 66.375 62.925 ;
        RECT 66.665 62.755 68.665 62.925 ;
        RECT 69.395 62.235 69.565 72.085 ;
        RECT 70.295 71.395 72.295 71.565 ;
        RECT 72.585 71.395 74.585 71.565 ;
        RECT 74.875 71.395 76.875 71.565 ;
        RECT 77.165 71.395 79.165 71.565 ;
        RECT 79.455 71.395 81.455 71.565 ;
        RECT 81.745 71.395 83.745 71.565 ;
        RECT 84.035 71.395 86.035 71.565 ;
        RECT 86.325 71.395 88.325 71.565 ;
        RECT 70.065 63.140 70.235 71.180 ;
        RECT 72.355 63.140 72.525 71.180 ;
        RECT 74.645 63.140 74.815 71.180 ;
        RECT 76.935 63.140 77.105 71.180 ;
        RECT 79.225 63.140 79.395 71.180 ;
        RECT 81.515 63.140 81.685 71.180 ;
        RECT 83.805 63.140 83.975 71.180 ;
        RECT 86.095 63.140 86.265 71.180 ;
        RECT 88.385 63.140 88.555 71.180 ;
        RECT 70.295 62.755 72.295 62.925 ;
        RECT 72.585 62.755 74.585 62.925 ;
        RECT 74.875 62.755 76.875 62.925 ;
        RECT 77.165 62.755 79.165 62.925 ;
        RECT 79.455 62.755 81.455 62.925 ;
        RECT 81.745 62.755 83.745 62.925 ;
        RECT 84.035 62.755 86.035 62.925 ;
        RECT 86.325 62.755 88.325 62.925 ;
        RECT 89.055 62.235 89.225 72.085 ;
        RECT 89.955 71.395 91.955 71.565 ;
        RECT 92.245 71.395 94.245 71.565 ;
        RECT 94.535 71.395 96.535 71.565 ;
        RECT 96.825 71.395 98.825 71.565 ;
        RECT 99.115 71.395 101.115 71.565 ;
        RECT 101.405 71.395 103.405 71.565 ;
        RECT 103.695 71.395 105.695 71.565 ;
        RECT 105.985 71.395 107.985 71.565 ;
        RECT 89.725 63.140 89.895 71.180 ;
        RECT 92.015 63.140 92.185 71.180 ;
        RECT 94.305 63.140 94.475 71.180 ;
        RECT 96.595 63.140 96.765 71.180 ;
        RECT 98.885 63.140 99.055 71.180 ;
        RECT 101.175 63.140 101.345 71.180 ;
        RECT 103.465 63.140 103.635 71.180 ;
        RECT 105.755 63.140 105.925 71.180 ;
        RECT 108.045 63.140 108.215 71.180 ;
        RECT 89.955 62.755 91.955 62.925 ;
        RECT 92.245 62.755 94.245 62.925 ;
        RECT 94.535 62.755 96.535 62.925 ;
        RECT 96.825 62.755 98.825 62.925 ;
        RECT 99.115 62.755 101.115 62.925 ;
        RECT 101.405 62.755 103.405 62.925 ;
        RECT 103.695 62.755 105.695 62.925 ;
        RECT 105.985 62.755 107.985 62.925 ;
        RECT 108.715 62.235 108.885 72.085 ;
        RECT 109.615 71.395 111.615 71.565 ;
        RECT 111.905 71.395 113.905 71.565 ;
        RECT 114.195 71.395 116.195 71.565 ;
        RECT 116.485 71.395 118.485 71.565 ;
        RECT 118.775 71.395 120.775 71.565 ;
        RECT 121.065 71.395 123.065 71.565 ;
        RECT 123.355 71.395 125.355 71.565 ;
        RECT 125.645 71.395 127.645 71.565 ;
        RECT 109.385 63.140 109.555 71.180 ;
        RECT 111.675 63.140 111.845 71.180 ;
        RECT 113.965 63.140 114.135 71.180 ;
        RECT 116.255 63.140 116.425 71.180 ;
        RECT 118.545 63.140 118.715 71.180 ;
        RECT 120.835 63.140 121.005 71.180 ;
        RECT 123.125 63.140 123.295 71.180 ;
        RECT 125.415 63.140 125.585 71.180 ;
        RECT 127.705 63.140 127.875 71.180 ;
        RECT 109.615 62.755 111.615 62.925 ;
        RECT 111.905 62.755 113.905 62.925 ;
        RECT 114.195 62.755 116.195 62.925 ;
        RECT 116.485 62.755 118.485 62.925 ;
        RECT 118.775 62.755 120.775 62.925 ;
        RECT 121.065 62.755 123.065 62.925 ;
        RECT 123.355 62.755 125.355 62.925 ;
        RECT 125.645 62.755 127.645 62.925 ;
        RECT 128.375 62.235 128.905 72.085 ;
        RECT 10.055 62.065 128.905 62.235 ;
        RECT 10.055 52.215 10.585 62.065 ;
        RECT 11.315 61.375 13.315 61.545 ;
        RECT 13.605 61.375 15.605 61.545 ;
        RECT 15.895 61.375 17.895 61.545 ;
        RECT 18.185 61.375 20.185 61.545 ;
        RECT 20.475 61.375 22.475 61.545 ;
        RECT 22.765 61.375 24.765 61.545 ;
        RECT 25.055 61.375 27.055 61.545 ;
        RECT 27.345 61.375 29.345 61.545 ;
        RECT 11.085 53.120 11.255 61.160 ;
        RECT 13.375 53.120 13.545 61.160 ;
        RECT 15.665 53.120 15.835 61.160 ;
        RECT 17.955 53.120 18.125 61.160 ;
        RECT 20.245 53.120 20.415 61.160 ;
        RECT 22.535 53.120 22.705 61.160 ;
        RECT 24.825 53.120 24.995 61.160 ;
        RECT 27.115 53.120 27.285 61.160 ;
        RECT 29.405 53.120 29.575 61.160 ;
        RECT 11.315 52.735 13.315 52.905 ;
        RECT 13.605 52.735 15.605 52.905 ;
        RECT 15.895 52.735 17.895 52.905 ;
        RECT 18.185 52.735 20.185 52.905 ;
        RECT 20.475 52.735 22.475 52.905 ;
        RECT 22.765 52.735 24.765 52.905 ;
        RECT 25.055 52.735 27.055 52.905 ;
        RECT 27.345 52.735 29.345 52.905 ;
        RECT 30.075 52.215 30.245 62.065 ;
        RECT 30.975 61.375 32.975 61.545 ;
        RECT 33.265 61.375 35.265 61.545 ;
        RECT 35.555 61.375 37.555 61.545 ;
        RECT 37.845 61.375 39.845 61.545 ;
        RECT 40.135 61.375 42.135 61.545 ;
        RECT 42.425 61.375 44.425 61.545 ;
        RECT 44.715 61.375 46.715 61.545 ;
        RECT 47.005 61.375 49.005 61.545 ;
        RECT 30.745 53.120 30.915 61.160 ;
        RECT 33.035 53.120 33.205 61.160 ;
        RECT 35.325 53.120 35.495 61.160 ;
        RECT 37.615 53.120 37.785 61.160 ;
        RECT 39.905 53.120 40.075 61.160 ;
        RECT 42.195 53.120 42.365 61.160 ;
        RECT 44.485 53.120 44.655 61.160 ;
        RECT 46.775 53.120 46.945 61.160 ;
        RECT 49.065 53.120 49.235 61.160 ;
        RECT 30.975 52.735 32.975 52.905 ;
        RECT 33.265 52.735 35.265 52.905 ;
        RECT 35.555 52.735 37.555 52.905 ;
        RECT 37.845 52.735 39.845 52.905 ;
        RECT 40.135 52.735 42.135 52.905 ;
        RECT 42.425 52.735 44.425 52.905 ;
        RECT 44.715 52.735 46.715 52.905 ;
        RECT 47.005 52.735 49.005 52.905 ;
        RECT 49.735 52.215 49.905 62.065 ;
        RECT 50.635 61.375 52.635 61.545 ;
        RECT 52.925 61.375 54.925 61.545 ;
        RECT 55.215 61.375 57.215 61.545 ;
        RECT 57.505 61.375 59.505 61.545 ;
        RECT 59.795 61.375 61.795 61.545 ;
        RECT 62.085 61.375 64.085 61.545 ;
        RECT 64.375 61.375 66.375 61.545 ;
        RECT 66.665 61.375 68.665 61.545 ;
        RECT 50.405 53.120 50.575 61.160 ;
        RECT 52.695 53.120 52.865 61.160 ;
        RECT 54.985 53.120 55.155 61.160 ;
        RECT 57.275 53.120 57.445 61.160 ;
        RECT 59.565 53.120 59.735 61.160 ;
        RECT 61.855 53.120 62.025 61.160 ;
        RECT 64.145 53.120 64.315 61.160 ;
        RECT 66.435 53.120 66.605 61.160 ;
        RECT 68.725 53.120 68.895 61.160 ;
        RECT 50.635 52.735 52.635 52.905 ;
        RECT 52.925 52.735 54.925 52.905 ;
        RECT 55.215 52.735 57.215 52.905 ;
        RECT 57.505 52.735 59.505 52.905 ;
        RECT 59.795 52.735 61.795 52.905 ;
        RECT 62.085 52.735 64.085 52.905 ;
        RECT 64.375 52.735 66.375 52.905 ;
        RECT 66.665 52.735 68.665 52.905 ;
        RECT 69.395 52.215 69.565 62.065 ;
        RECT 70.295 61.375 72.295 61.545 ;
        RECT 72.585 61.375 74.585 61.545 ;
        RECT 74.875 61.375 76.875 61.545 ;
        RECT 77.165 61.375 79.165 61.545 ;
        RECT 79.455 61.375 81.455 61.545 ;
        RECT 81.745 61.375 83.745 61.545 ;
        RECT 84.035 61.375 86.035 61.545 ;
        RECT 86.325 61.375 88.325 61.545 ;
        RECT 70.065 53.120 70.235 61.160 ;
        RECT 72.355 53.120 72.525 61.160 ;
        RECT 74.645 53.120 74.815 61.160 ;
        RECT 76.935 53.120 77.105 61.160 ;
        RECT 79.225 53.120 79.395 61.160 ;
        RECT 81.515 53.120 81.685 61.160 ;
        RECT 83.805 53.120 83.975 61.160 ;
        RECT 86.095 53.120 86.265 61.160 ;
        RECT 88.385 53.120 88.555 61.160 ;
        RECT 70.295 52.735 72.295 52.905 ;
        RECT 72.585 52.735 74.585 52.905 ;
        RECT 74.875 52.735 76.875 52.905 ;
        RECT 77.165 52.735 79.165 52.905 ;
        RECT 79.455 52.735 81.455 52.905 ;
        RECT 81.745 52.735 83.745 52.905 ;
        RECT 84.035 52.735 86.035 52.905 ;
        RECT 86.325 52.735 88.325 52.905 ;
        RECT 89.055 52.215 89.225 62.065 ;
        RECT 89.955 61.375 91.955 61.545 ;
        RECT 92.245 61.375 94.245 61.545 ;
        RECT 94.535 61.375 96.535 61.545 ;
        RECT 96.825 61.375 98.825 61.545 ;
        RECT 99.115 61.375 101.115 61.545 ;
        RECT 101.405 61.375 103.405 61.545 ;
        RECT 103.695 61.375 105.695 61.545 ;
        RECT 105.985 61.375 107.985 61.545 ;
        RECT 89.725 53.120 89.895 61.160 ;
        RECT 92.015 53.120 92.185 61.160 ;
        RECT 94.305 53.120 94.475 61.160 ;
        RECT 96.595 53.120 96.765 61.160 ;
        RECT 98.885 53.120 99.055 61.160 ;
        RECT 101.175 53.120 101.345 61.160 ;
        RECT 103.465 53.120 103.635 61.160 ;
        RECT 105.755 53.120 105.925 61.160 ;
        RECT 108.045 53.120 108.215 61.160 ;
        RECT 89.955 52.735 91.955 52.905 ;
        RECT 92.245 52.735 94.245 52.905 ;
        RECT 94.535 52.735 96.535 52.905 ;
        RECT 96.825 52.735 98.825 52.905 ;
        RECT 99.115 52.735 101.115 52.905 ;
        RECT 101.405 52.735 103.405 52.905 ;
        RECT 103.695 52.735 105.695 52.905 ;
        RECT 105.985 52.735 107.985 52.905 ;
        RECT 108.715 52.215 108.885 62.065 ;
        RECT 109.615 61.375 111.615 61.545 ;
        RECT 111.905 61.375 113.905 61.545 ;
        RECT 114.195 61.375 116.195 61.545 ;
        RECT 116.485 61.375 118.485 61.545 ;
        RECT 118.775 61.375 120.775 61.545 ;
        RECT 121.065 61.375 123.065 61.545 ;
        RECT 123.355 61.375 125.355 61.545 ;
        RECT 125.645 61.375 127.645 61.545 ;
        RECT 109.385 53.120 109.555 61.160 ;
        RECT 111.675 53.120 111.845 61.160 ;
        RECT 113.965 53.120 114.135 61.160 ;
        RECT 116.255 53.120 116.425 61.160 ;
        RECT 118.545 53.120 118.715 61.160 ;
        RECT 120.835 53.120 121.005 61.160 ;
        RECT 123.125 53.120 123.295 61.160 ;
        RECT 125.415 53.120 125.585 61.160 ;
        RECT 127.705 53.120 127.875 61.160 ;
        RECT 109.615 52.735 111.615 52.905 ;
        RECT 111.905 52.735 113.905 52.905 ;
        RECT 114.195 52.735 116.195 52.905 ;
        RECT 116.485 52.735 118.485 52.905 ;
        RECT 118.775 52.735 120.775 52.905 ;
        RECT 121.065 52.735 123.065 52.905 ;
        RECT 123.355 52.735 125.355 52.905 ;
        RECT 125.645 52.735 127.645 52.905 ;
        RECT 128.375 52.215 128.905 62.065 ;
        RECT 10.055 52.045 128.905 52.215 ;
        RECT 10.055 42.195 10.585 52.045 ;
        RECT 11.315 51.355 13.315 51.525 ;
        RECT 13.605 51.355 15.605 51.525 ;
        RECT 15.895 51.355 17.895 51.525 ;
        RECT 18.185 51.355 20.185 51.525 ;
        RECT 20.475 51.355 22.475 51.525 ;
        RECT 22.765 51.355 24.765 51.525 ;
        RECT 25.055 51.355 27.055 51.525 ;
        RECT 27.345 51.355 29.345 51.525 ;
        RECT 11.085 43.100 11.255 51.140 ;
        RECT 13.375 43.100 13.545 51.140 ;
        RECT 15.665 43.100 15.835 51.140 ;
        RECT 17.955 43.100 18.125 51.140 ;
        RECT 20.245 43.100 20.415 51.140 ;
        RECT 22.535 43.100 22.705 51.140 ;
        RECT 24.825 43.100 24.995 51.140 ;
        RECT 27.115 43.100 27.285 51.140 ;
        RECT 29.405 43.100 29.575 51.140 ;
        RECT 11.315 42.715 13.315 42.885 ;
        RECT 13.605 42.715 15.605 42.885 ;
        RECT 15.895 42.715 17.895 42.885 ;
        RECT 18.185 42.715 20.185 42.885 ;
        RECT 20.475 42.715 22.475 42.885 ;
        RECT 22.765 42.715 24.765 42.885 ;
        RECT 25.055 42.715 27.055 42.885 ;
        RECT 27.345 42.715 29.345 42.885 ;
        RECT 30.075 42.195 30.245 52.045 ;
        RECT 30.975 51.355 32.975 51.525 ;
        RECT 33.265 51.355 35.265 51.525 ;
        RECT 35.555 51.355 37.555 51.525 ;
        RECT 37.845 51.355 39.845 51.525 ;
        RECT 40.135 51.355 42.135 51.525 ;
        RECT 42.425 51.355 44.425 51.525 ;
        RECT 44.715 51.355 46.715 51.525 ;
        RECT 47.005 51.355 49.005 51.525 ;
        RECT 30.745 43.100 30.915 51.140 ;
        RECT 33.035 43.100 33.205 51.140 ;
        RECT 35.325 43.100 35.495 51.140 ;
        RECT 37.615 43.100 37.785 51.140 ;
        RECT 39.905 43.100 40.075 51.140 ;
        RECT 42.195 43.100 42.365 51.140 ;
        RECT 44.485 43.100 44.655 51.140 ;
        RECT 46.775 43.100 46.945 51.140 ;
        RECT 49.065 43.100 49.235 51.140 ;
        RECT 30.975 42.715 32.975 42.885 ;
        RECT 33.265 42.715 35.265 42.885 ;
        RECT 35.555 42.715 37.555 42.885 ;
        RECT 37.845 42.715 39.845 42.885 ;
        RECT 40.135 42.715 42.135 42.885 ;
        RECT 42.425 42.715 44.425 42.885 ;
        RECT 44.715 42.715 46.715 42.885 ;
        RECT 47.005 42.715 49.005 42.885 ;
        RECT 49.735 42.195 49.905 52.045 ;
        RECT 50.635 51.355 52.635 51.525 ;
        RECT 52.925 51.355 54.925 51.525 ;
        RECT 55.215 51.355 57.215 51.525 ;
        RECT 57.505 51.355 59.505 51.525 ;
        RECT 59.795 51.355 61.795 51.525 ;
        RECT 62.085 51.355 64.085 51.525 ;
        RECT 64.375 51.355 66.375 51.525 ;
        RECT 66.665 51.355 68.665 51.525 ;
        RECT 50.405 43.100 50.575 51.140 ;
        RECT 52.695 43.100 52.865 51.140 ;
        RECT 54.985 43.100 55.155 51.140 ;
        RECT 57.275 43.100 57.445 51.140 ;
        RECT 59.565 43.100 59.735 51.140 ;
        RECT 61.855 43.100 62.025 51.140 ;
        RECT 64.145 43.100 64.315 51.140 ;
        RECT 66.435 43.100 66.605 51.140 ;
        RECT 68.725 43.100 68.895 51.140 ;
        RECT 50.635 42.715 52.635 42.885 ;
        RECT 52.925 42.715 54.925 42.885 ;
        RECT 55.215 42.715 57.215 42.885 ;
        RECT 57.505 42.715 59.505 42.885 ;
        RECT 59.795 42.715 61.795 42.885 ;
        RECT 62.085 42.715 64.085 42.885 ;
        RECT 64.375 42.715 66.375 42.885 ;
        RECT 66.665 42.715 68.665 42.885 ;
        RECT 69.395 42.195 69.565 52.045 ;
        RECT 70.295 51.355 72.295 51.525 ;
        RECT 72.585 51.355 74.585 51.525 ;
        RECT 74.875 51.355 76.875 51.525 ;
        RECT 77.165 51.355 79.165 51.525 ;
        RECT 79.455 51.355 81.455 51.525 ;
        RECT 81.745 51.355 83.745 51.525 ;
        RECT 84.035 51.355 86.035 51.525 ;
        RECT 86.325 51.355 88.325 51.525 ;
        RECT 70.065 43.100 70.235 51.140 ;
        RECT 72.355 43.100 72.525 51.140 ;
        RECT 74.645 43.100 74.815 51.140 ;
        RECT 76.935 43.100 77.105 51.140 ;
        RECT 79.225 43.100 79.395 51.140 ;
        RECT 81.515 43.100 81.685 51.140 ;
        RECT 83.805 43.100 83.975 51.140 ;
        RECT 86.095 43.100 86.265 51.140 ;
        RECT 88.385 43.100 88.555 51.140 ;
        RECT 70.295 42.715 72.295 42.885 ;
        RECT 72.585 42.715 74.585 42.885 ;
        RECT 74.875 42.715 76.875 42.885 ;
        RECT 77.165 42.715 79.165 42.885 ;
        RECT 79.455 42.715 81.455 42.885 ;
        RECT 81.745 42.715 83.745 42.885 ;
        RECT 84.035 42.715 86.035 42.885 ;
        RECT 86.325 42.715 88.325 42.885 ;
        RECT 89.055 42.195 89.225 52.045 ;
        RECT 89.955 51.355 91.955 51.525 ;
        RECT 92.245 51.355 94.245 51.525 ;
        RECT 94.535 51.355 96.535 51.525 ;
        RECT 96.825 51.355 98.825 51.525 ;
        RECT 99.115 51.355 101.115 51.525 ;
        RECT 101.405 51.355 103.405 51.525 ;
        RECT 103.695 51.355 105.695 51.525 ;
        RECT 105.985 51.355 107.985 51.525 ;
        RECT 89.725 43.100 89.895 51.140 ;
        RECT 92.015 43.100 92.185 51.140 ;
        RECT 94.305 43.100 94.475 51.140 ;
        RECT 96.595 43.100 96.765 51.140 ;
        RECT 98.885 43.100 99.055 51.140 ;
        RECT 101.175 43.100 101.345 51.140 ;
        RECT 103.465 43.100 103.635 51.140 ;
        RECT 105.755 43.100 105.925 51.140 ;
        RECT 108.045 43.100 108.215 51.140 ;
        RECT 89.955 42.715 91.955 42.885 ;
        RECT 92.245 42.715 94.245 42.885 ;
        RECT 94.535 42.715 96.535 42.885 ;
        RECT 96.825 42.715 98.825 42.885 ;
        RECT 99.115 42.715 101.115 42.885 ;
        RECT 101.405 42.715 103.405 42.885 ;
        RECT 103.695 42.715 105.695 42.885 ;
        RECT 105.985 42.715 107.985 42.885 ;
        RECT 108.715 42.195 108.885 52.045 ;
        RECT 109.615 51.355 111.615 51.525 ;
        RECT 111.905 51.355 113.905 51.525 ;
        RECT 114.195 51.355 116.195 51.525 ;
        RECT 116.485 51.355 118.485 51.525 ;
        RECT 118.775 51.355 120.775 51.525 ;
        RECT 121.065 51.355 123.065 51.525 ;
        RECT 123.355 51.355 125.355 51.525 ;
        RECT 125.645 51.355 127.645 51.525 ;
        RECT 109.385 43.100 109.555 51.140 ;
        RECT 111.675 43.100 111.845 51.140 ;
        RECT 113.965 43.100 114.135 51.140 ;
        RECT 116.255 43.100 116.425 51.140 ;
        RECT 118.545 43.100 118.715 51.140 ;
        RECT 120.835 43.100 121.005 51.140 ;
        RECT 123.125 43.100 123.295 51.140 ;
        RECT 125.415 43.100 125.585 51.140 ;
        RECT 127.705 43.100 127.875 51.140 ;
        RECT 109.615 42.715 111.615 42.885 ;
        RECT 111.905 42.715 113.905 42.885 ;
        RECT 114.195 42.715 116.195 42.885 ;
        RECT 116.485 42.715 118.485 42.885 ;
        RECT 118.775 42.715 120.775 42.885 ;
        RECT 121.065 42.715 123.065 42.885 ;
        RECT 123.355 42.715 125.355 42.885 ;
        RECT 125.645 42.715 127.645 42.885 ;
        RECT 128.375 42.195 128.905 52.045 ;
        RECT 10.055 41.665 128.905 42.195 ;
        RECT 10.055 39.070 74.665 39.600 ;
        RECT 10.055 29.310 10.585 39.070 ;
        RECT 11.375 38.380 13.375 38.550 ;
        RECT 13.665 38.380 15.665 38.550 ;
        RECT 15.955 38.380 17.955 38.550 ;
        RECT 18.245 38.380 20.245 38.550 ;
        RECT 11.145 30.170 11.315 38.210 ;
        RECT 13.435 30.170 13.605 38.210 ;
        RECT 15.725 30.170 15.895 38.210 ;
        RECT 18.015 30.170 18.185 38.210 ;
        RECT 20.305 30.170 20.475 38.210 ;
        RECT 11.375 29.830 13.375 30.000 ;
        RECT 13.665 29.830 15.665 30.000 ;
        RECT 15.955 29.830 17.955 30.000 ;
        RECT 18.245 29.830 20.245 30.000 ;
        RECT 21.035 29.310 21.205 39.070 ;
        RECT 21.995 38.380 23.995 38.550 ;
        RECT 24.285 38.380 26.285 38.550 ;
        RECT 26.575 38.380 28.575 38.550 ;
        RECT 28.865 38.380 30.865 38.550 ;
        RECT 21.765 30.170 21.935 38.210 ;
        RECT 24.055 30.170 24.225 38.210 ;
        RECT 26.345 30.170 26.515 38.210 ;
        RECT 28.635 30.170 28.805 38.210 ;
        RECT 30.925 30.170 31.095 38.210 ;
        RECT 21.995 29.830 23.995 30.000 ;
        RECT 24.285 29.830 26.285 30.000 ;
        RECT 26.575 29.830 28.575 30.000 ;
        RECT 28.865 29.830 30.865 30.000 ;
        RECT 31.655 29.310 31.825 39.070 ;
        RECT 32.615 38.380 34.615 38.550 ;
        RECT 34.905 38.380 36.905 38.550 ;
        RECT 37.195 38.380 39.195 38.550 ;
        RECT 39.485 38.380 41.485 38.550 ;
        RECT 32.385 30.170 32.555 38.210 ;
        RECT 34.675 30.170 34.845 38.210 ;
        RECT 36.965 30.170 37.135 38.210 ;
        RECT 39.255 30.170 39.425 38.210 ;
        RECT 41.545 30.170 41.715 38.210 ;
        RECT 32.615 29.830 34.615 30.000 ;
        RECT 34.905 29.830 36.905 30.000 ;
        RECT 37.195 29.830 39.195 30.000 ;
        RECT 39.485 29.830 41.485 30.000 ;
        RECT 42.275 29.310 42.445 39.070 ;
        RECT 43.235 38.380 45.235 38.550 ;
        RECT 45.525 38.380 47.525 38.550 ;
        RECT 47.815 38.380 49.815 38.550 ;
        RECT 50.105 38.380 52.105 38.550 ;
        RECT 43.005 30.170 43.175 38.210 ;
        RECT 45.295 30.170 45.465 38.210 ;
        RECT 47.585 30.170 47.755 38.210 ;
        RECT 49.875 30.170 50.045 38.210 ;
        RECT 52.165 30.170 52.335 38.210 ;
        RECT 43.235 29.830 45.235 30.000 ;
        RECT 45.525 29.830 47.525 30.000 ;
        RECT 47.815 29.830 49.815 30.000 ;
        RECT 50.105 29.830 52.105 30.000 ;
        RECT 52.895 29.310 53.065 39.070 ;
        RECT 53.855 38.380 55.855 38.550 ;
        RECT 56.145 38.380 58.145 38.550 ;
        RECT 58.435 38.380 60.435 38.550 ;
        RECT 60.725 38.380 62.725 38.550 ;
        RECT 53.625 30.170 53.795 38.210 ;
        RECT 55.915 30.170 56.085 38.210 ;
        RECT 58.205 30.170 58.375 38.210 ;
        RECT 60.495 30.170 60.665 38.210 ;
        RECT 62.785 30.170 62.955 38.210 ;
        RECT 53.855 29.830 55.855 30.000 ;
        RECT 56.145 29.830 58.145 30.000 ;
        RECT 58.435 29.830 60.435 30.000 ;
        RECT 60.725 29.830 62.725 30.000 ;
        RECT 63.515 29.310 63.685 39.070 ;
        RECT 64.475 38.380 66.475 38.550 ;
        RECT 66.765 38.380 68.765 38.550 ;
        RECT 69.055 38.380 71.055 38.550 ;
        RECT 71.345 38.380 73.345 38.550 ;
        RECT 64.245 30.170 64.415 38.210 ;
        RECT 66.535 30.170 66.705 38.210 ;
        RECT 68.825 30.170 68.995 38.210 ;
        RECT 71.115 30.170 71.285 38.210 ;
        RECT 73.405 30.170 73.575 38.210 ;
        RECT 64.475 29.830 66.475 30.000 ;
        RECT 66.765 29.830 68.765 30.000 ;
        RECT 69.055 29.830 71.055 30.000 ;
        RECT 71.345 29.830 73.345 30.000 ;
        RECT 74.135 29.310 74.665 39.070 ;
        RECT 10.055 29.140 74.665 29.310 ;
        RECT 10.055 19.380 10.585 29.140 ;
        RECT 11.375 28.450 13.375 28.620 ;
        RECT 13.665 28.450 15.665 28.620 ;
        RECT 15.955 28.450 17.955 28.620 ;
        RECT 18.245 28.450 20.245 28.620 ;
        RECT 11.145 20.240 11.315 28.280 ;
        RECT 13.435 20.240 13.605 28.280 ;
        RECT 15.725 20.240 15.895 28.280 ;
        RECT 18.015 20.240 18.185 28.280 ;
        RECT 20.305 20.240 20.475 28.280 ;
        RECT 11.375 19.900 13.375 20.070 ;
        RECT 13.665 19.900 15.665 20.070 ;
        RECT 15.955 19.900 17.955 20.070 ;
        RECT 18.245 19.900 20.245 20.070 ;
        RECT 21.035 19.380 21.205 29.140 ;
        RECT 21.995 28.450 23.995 28.620 ;
        RECT 24.285 28.450 26.285 28.620 ;
        RECT 26.575 28.450 28.575 28.620 ;
        RECT 28.865 28.450 30.865 28.620 ;
        RECT 21.765 20.240 21.935 28.280 ;
        RECT 24.055 20.240 24.225 28.280 ;
        RECT 26.345 20.240 26.515 28.280 ;
        RECT 28.635 20.240 28.805 28.280 ;
        RECT 30.925 20.240 31.095 28.280 ;
        RECT 21.995 19.900 23.995 20.070 ;
        RECT 24.285 19.900 26.285 20.070 ;
        RECT 26.575 19.900 28.575 20.070 ;
        RECT 28.865 19.900 30.865 20.070 ;
        RECT 31.655 19.380 31.825 29.140 ;
        RECT 32.615 28.450 34.615 28.620 ;
        RECT 34.905 28.450 36.905 28.620 ;
        RECT 37.195 28.450 39.195 28.620 ;
        RECT 39.485 28.450 41.485 28.620 ;
        RECT 32.385 20.240 32.555 28.280 ;
        RECT 34.675 20.240 34.845 28.280 ;
        RECT 36.965 20.240 37.135 28.280 ;
        RECT 39.255 20.240 39.425 28.280 ;
        RECT 41.545 20.240 41.715 28.280 ;
        RECT 32.615 19.900 34.615 20.070 ;
        RECT 34.905 19.900 36.905 20.070 ;
        RECT 37.195 19.900 39.195 20.070 ;
        RECT 39.485 19.900 41.485 20.070 ;
        RECT 42.275 19.380 42.445 29.140 ;
        RECT 43.235 28.450 45.235 28.620 ;
        RECT 45.525 28.450 47.525 28.620 ;
        RECT 47.815 28.450 49.815 28.620 ;
        RECT 50.105 28.450 52.105 28.620 ;
        RECT 43.005 20.240 43.175 28.280 ;
        RECT 45.295 20.240 45.465 28.280 ;
        RECT 47.585 20.240 47.755 28.280 ;
        RECT 49.875 20.240 50.045 28.280 ;
        RECT 52.165 20.240 52.335 28.280 ;
        RECT 43.235 19.900 45.235 20.070 ;
        RECT 45.525 19.900 47.525 20.070 ;
        RECT 47.815 19.900 49.815 20.070 ;
        RECT 50.105 19.900 52.105 20.070 ;
        RECT 52.895 19.380 53.065 29.140 ;
        RECT 53.855 28.450 55.855 28.620 ;
        RECT 56.145 28.450 58.145 28.620 ;
        RECT 58.435 28.450 60.435 28.620 ;
        RECT 60.725 28.450 62.725 28.620 ;
        RECT 53.625 20.240 53.795 28.280 ;
        RECT 55.915 20.240 56.085 28.280 ;
        RECT 58.205 20.240 58.375 28.280 ;
        RECT 60.495 20.240 60.665 28.280 ;
        RECT 62.785 20.240 62.955 28.280 ;
        RECT 53.855 19.900 55.855 20.070 ;
        RECT 56.145 19.900 58.145 20.070 ;
        RECT 58.435 19.900 60.435 20.070 ;
        RECT 60.725 19.900 62.725 20.070 ;
        RECT 63.515 19.380 63.685 29.140 ;
        RECT 64.475 28.450 66.475 28.620 ;
        RECT 66.765 28.450 68.765 28.620 ;
        RECT 69.055 28.450 71.055 28.620 ;
        RECT 71.345 28.450 73.345 28.620 ;
        RECT 64.245 20.240 64.415 28.280 ;
        RECT 66.535 20.240 66.705 28.280 ;
        RECT 68.825 20.240 68.995 28.280 ;
        RECT 71.115 20.240 71.285 28.280 ;
        RECT 73.405 20.240 73.575 28.280 ;
        RECT 64.475 19.900 66.475 20.070 ;
        RECT 66.765 19.900 68.765 20.070 ;
        RECT 69.055 19.900 71.055 20.070 ;
        RECT 71.345 19.900 73.345 20.070 ;
        RECT 74.135 19.380 74.665 29.140 ;
        RECT 10.055 19.210 74.665 19.380 ;
        RECT 10.055 9.450 10.585 19.210 ;
        RECT 11.375 18.520 13.375 18.690 ;
        RECT 13.665 18.520 15.665 18.690 ;
        RECT 15.955 18.520 17.955 18.690 ;
        RECT 18.245 18.520 20.245 18.690 ;
        RECT 11.145 10.310 11.315 18.350 ;
        RECT 13.435 10.310 13.605 18.350 ;
        RECT 15.725 10.310 15.895 18.350 ;
        RECT 18.015 10.310 18.185 18.350 ;
        RECT 20.305 10.310 20.475 18.350 ;
        RECT 11.375 9.970 13.375 10.140 ;
        RECT 13.665 9.970 15.665 10.140 ;
        RECT 15.955 9.970 17.955 10.140 ;
        RECT 18.245 9.970 20.245 10.140 ;
        RECT 21.035 9.450 21.205 19.210 ;
        RECT 21.995 18.520 23.995 18.690 ;
        RECT 24.285 18.520 26.285 18.690 ;
        RECT 26.575 18.520 28.575 18.690 ;
        RECT 28.865 18.520 30.865 18.690 ;
        RECT 21.765 10.310 21.935 18.350 ;
        RECT 24.055 10.310 24.225 18.350 ;
        RECT 26.345 10.310 26.515 18.350 ;
        RECT 28.635 10.310 28.805 18.350 ;
        RECT 30.925 10.310 31.095 18.350 ;
        RECT 21.995 9.970 23.995 10.140 ;
        RECT 24.285 9.970 26.285 10.140 ;
        RECT 26.575 9.970 28.575 10.140 ;
        RECT 28.865 9.970 30.865 10.140 ;
        RECT 31.655 9.450 31.825 19.210 ;
        RECT 32.615 18.520 34.615 18.690 ;
        RECT 34.905 18.520 36.905 18.690 ;
        RECT 37.195 18.520 39.195 18.690 ;
        RECT 39.485 18.520 41.485 18.690 ;
        RECT 32.385 10.310 32.555 18.350 ;
        RECT 34.675 10.310 34.845 18.350 ;
        RECT 36.965 10.310 37.135 18.350 ;
        RECT 39.255 10.310 39.425 18.350 ;
        RECT 41.545 10.310 41.715 18.350 ;
        RECT 32.615 9.970 34.615 10.140 ;
        RECT 34.905 9.970 36.905 10.140 ;
        RECT 37.195 9.970 39.195 10.140 ;
        RECT 39.485 9.970 41.485 10.140 ;
        RECT 42.275 9.450 42.445 19.210 ;
        RECT 43.235 18.520 45.235 18.690 ;
        RECT 45.525 18.520 47.525 18.690 ;
        RECT 47.815 18.520 49.815 18.690 ;
        RECT 50.105 18.520 52.105 18.690 ;
        RECT 43.005 10.310 43.175 18.350 ;
        RECT 45.295 10.310 45.465 18.350 ;
        RECT 47.585 10.310 47.755 18.350 ;
        RECT 49.875 10.310 50.045 18.350 ;
        RECT 52.165 10.310 52.335 18.350 ;
        RECT 43.235 9.970 45.235 10.140 ;
        RECT 45.525 9.970 47.525 10.140 ;
        RECT 47.815 9.970 49.815 10.140 ;
        RECT 50.105 9.970 52.105 10.140 ;
        RECT 52.895 9.450 53.065 19.210 ;
        RECT 53.855 18.520 55.855 18.690 ;
        RECT 56.145 18.520 58.145 18.690 ;
        RECT 58.435 18.520 60.435 18.690 ;
        RECT 60.725 18.520 62.725 18.690 ;
        RECT 53.625 10.310 53.795 18.350 ;
        RECT 55.915 10.310 56.085 18.350 ;
        RECT 58.205 10.310 58.375 18.350 ;
        RECT 60.495 10.310 60.665 18.350 ;
        RECT 62.785 10.310 62.955 18.350 ;
        RECT 53.855 9.970 55.855 10.140 ;
        RECT 56.145 9.970 58.145 10.140 ;
        RECT 58.435 9.970 60.435 10.140 ;
        RECT 60.725 9.970 62.725 10.140 ;
        RECT 63.515 9.450 63.685 19.210 ;
        RECT 64.475 18.520 66.475 18.690 ;
        RECT 66.765 18.520 68.765 18.690 ;
        RECT 69.055 18.520 71.055 18.690 ;
        RECT 71.345 18.520 73.345 18.690 ;
        RECT 64.245 10.310 64.415 18.350 ;
        RECT 66.535 10.310 66.705 18.350 ;
        RECT 68.825 10.310 68.995 18.350 ;
        RECT 71.115 10.310 71.285 18.350 ;
        RECT 73.405 10.310 73.575 18.350 ;
        RECT 64.475 9.970 66.475 10.140 ;
        RECT 66.765 9.970 68.765 10.140 ;
        RECT 69.055 9.970 71.055 10.140 ;
        RECT 71.345 9.970 73.345 10.140 ;
        RECT 74.135 9.450 74.665 19.210 ;
        RECT 10.055 8.920 74.665 9.450 ;
        RECT 79.695 39.070 128.905 39.600 ;
        RECT 79.695 29.310 80.225 39.070 ;
        RECT 80.785 38.210 85.535 39.070 ;
        RECT 80.785 30.170 80.955 38.210 ;
        RECT 83.075 30.170 83.245 38.210 ;
        RECT 85.365 30.170 85.535 38.210 ;
        RECT 81.015 29.830 83.015 30.000 ;
        RECT 83.305 29.830 85.305 30.000 ;
        RECT 86.095 29.310 86.265 39.070 ;
        RECT 87.055 38.380 89.055 38.550 ;
        RECT 89.345 38.380 91.345 38.550 ;
        RECT 86.825 30.170 86.995 38.210 ;
        RECT 89.115 30.170 89.285 38.210 ;
        RECT 91.405 30.170 91.575 38.210 ;
        RECT 87.055 29.830 89.055 30.000 ;
        RECT 89.345 29.830 91.345 30.000 ;
        RECT 92.135 29.310 92.305 39.070 ;
        RECT 93.095 38.380 95.095 38.550 ;
        RECT 95.385 38.380 97.385 38.550 ;
        RECT 92.865 30.170 93.035 38.210 ;
        RECT 95.155 30.170 95.325 38.210 ;
        RECT 97.445 30.170 97.615 38.210 ;
        RECT 93.095 29.830 95.095 30.000 ;
        RECT 95.385 29.830 97.385 30.000 ;
        RECT 98.175 29.310 98.345 39.070 ;
        RECT 99.135 38.380 101.135 38.550 ;
        RECT 101.425 38.380 103.425 38.550 ;
        RECT 98.905 30.170 99.075 38.210 ;
        RECT 101.195 30.170 101.365 38.210 ;
        RECT 103.485 30.170 103.655 38.210 ;
        RECT 99.135 29.830 101.135 30.000 ;
        RECT 101.425 29.830 103.425 30.000 ;
        RECT 104.215 29.310 104.385 39.070 ;
        RECT 105.175 38.380 107.175 38.550 ;
        RECT 107.465 38.380 109.465 38.550 ;
        RECT 104.945 30.170 105.115 38.210 ;
        RECT 107.235 30.170 107.405 38.210 ;
        RECT 109.525 30.170 109.695 38.210 ;
        RECT 105.175 29.830 107.175 30.000 ;
        RECT 107.465 29.830 109.465 30.000 ;
        RECT 110.255 29.310 110.425 39.070 ;
        RECT 111.215 38.380 113.215 38.550 ;
        RECT 113.505 38.380 115.505 38.550 ;
        RECT 110.985 30.170 111.155 38.210 ;
        RECT 113.275 30.170 113.445 38.210 ;
        RECT 115.565 30.170 115.735 38.210 ;
        RECT 111.215 29.830 113.215 30.000 ;
        RECT 113.505 29.830 115.505 30.000 ;
        RECT 116.295 29.310 116.465 39.070 ;
        RECT 117.255 38.380 119.255 38.550 ;
        RECT 119.545 38.380 121.545 38.550 ;
        RECT 117.025 30.170 117.195 38.210 ;
        RECT 119.315 30.170 119.485 38.210 ;
        RECT 121.605 30.170 121.775 38.210 ;
        RECT 117.255 29.830 119.255 30.000 ;
        RECT 119.545 29.830 121.545 30.000 ;
        RECT 122.335 29.310 122.505 39.070 ;
        RECT 123.065 38.210 127.815 39.070 ;
        RECT 123.065 30.170 123.235 38.210 ;
        RECT 125.355 30.170 125.525 38.210 ;
        RECT 127.645 30.170 127.815 38.210 ;
        RECT 123.295 29.830 125.295 30.000 ;
        RECT 125.585 29.830 127.585 30.000 ;
        RECT 128.375 29.310 128.905 39.070 ;
        RECT 79.695 29.140 128.905 29.310 ;
        RECT 79.695 19.380 80.225 29.140 ;
        RECT 81.015 28.450 83.015 28.620 ;
        RECT 83.305 28.450 85.305 28.620 ;
        RECT 80.785 20.240 80.955 28.280 ;
        RECT 83.075 20.240 83.245 28.280 ;
        RECT 85.365 20.240 85.535 28.280 ;
        RECT 80.785 19.380 85.535 20.240 ;
        RECT 86.095 19.380 86.265 29.140 ;
        RECT 87.055 28.450 89.055 28.620 ;
        RECT 89.345 28.450 91.345 28.620 ;
        RECT 86.825 20.240 86.995 28.280 ;
        RECT 89.115 20.240 89.285 28.280 ;
        RECT 91.405 20.240 91.575 28.280 ;
        RECT 87.055 19.900 89.055 20.070 ;
        RECT 89.345 19.900 91.345 20.070 ;
        RECT 92.135 19.380 92.305 29.140 ;
        RECT 93.095 28.450 95.095 28.620 ;
        RECT 95.385 28.450 97.385 28.620 ;
        RECT 92.865 20.240 93.035 28.280 ;
        RECT 95.155 20.240 95.325 28.280 ;
        RECT 97.445 20.240 97.615 28.280 ;
        RECT 93.095 19.900 95.095 20.070 ;
        RECT 95.385 19.900 97.385 20.070 ;
        RECT 98.175 19.380 98.345 29.140 ;
        RECT 99.135 28.450 101.135 28.620 ;
        RECT 101.425 28.450 103.425 28.620 ;
        RECT 98.905 20.240 99.075 28.280 ;
        RECT 101.195 20.240 101.365 28.280 ;
        RECT 103.485 20.240 103.655 28.280 ;
        RECT 99.135 19.900 101.135 20.070 ;
        RECT 101.425 19.900 103.425 20.070 ;
        RECT 104.215 19.380 104.385 29.140 ;
        RECT 105.175 28.450 107.175 28.620 ;
        RECT 107.465 28.450 109.465 28.620 ;
        RECT 104.945 20.240 105.115 28.280 ;
        RECT 107.235 20.240 107.405 28.280 ;
        RECT 109.525 20.240 109.695 28.280 ;
        RECT 105.175 19.900 107.175 20.070 ;
        RECT 107.465 19.900 109.465 20.070 ;
        RECT 110.255 19.380 110.425 29.140 ;
        RECT 111.215 28.450 113.215 28.620 ;
        RECT 113.505 28.450 115.505 28.620 ;
        RECT 110.985 20.240 111.155 28.280 ;
        RECT 113.275 20.240 113.445 28.280 ;
        RECT 115.565 20.240 115.735 28.280 ;
        RECT 111.215 19.900 113.215 20.070 ;
        RECT 113.505 19.900 115.505 20.070 ;
        RECT 116.295 19.380 116.465 29.140 ;
        RECT 117.255 28.450 119.255 28.620 ;
        RECT 119.545 28.450 121.545 28.620 ;
        RECT 117.025 20.240 117.195 28.280 ;
        RECT 119.315 20.240 119.485 28.280 ;
        RECT 121.605 20.240 121.775 28.280 ;
        RECT 117.255 19.900 119.255 20.070 ;
        RECT 119.545 19.900 121.545 20.070 ;
        RECT 122.335 19.380 122.505 29.140 ;
        RECT 123.295 28.450 125.295 28.620 ;
        RECT 125.585 28.450 127.585 28.620 ;
        RECT 123.065 20.240 123.235 28.280 ;
        RECT 125.355 20.240 125.525 28.280 ;
        RECT 127.645 20.240 127.815 28.280 ;
        RECT 123.065 19.380 127.815 20.240 ;
        RECT 128.375 19.380 128.905 29.140 ;
        RECT 79.695 19.210 128.905 19.380 ;
        RECT 79.695 9.450 80.225 19.210 ;
        RECT 81.015 18.520 83.015 18.690 ;
        RECT 83.305 18.520 85.305 18.690 ;
        RECT 80.785 10.310 80.955 18.350 ;
        RECT 83.075 10.310 83.245 18.350 ;
        RECT 85.365 10.310 85.535 18.350 ;
        RECT 80.785 9.450 85.535 10.310 ;
        RECT 86.095 9.450 86.265 19.210 ;
        RECT 87.055 18.520 89.055 18.690 ;
        RECT 89.345 18.520 91.345 18.690 ;
        RECT 86.825 10.310 86.995 18.350 ;
        RECT 89.115 10.310 89.285 18.350 ;
        RECT 91.405 10.310 91.575 18.350 ;
        RECT 86.825 9.450 91.575 10.310 ;
        RECT 92.135 9.450 92.305 19.210 ;
        RECT 93.095 18.520 95.095 18.690 ;
        RECT 95.385 18.520 97.385 18.690 ;
        RECT 92.865 10.310 93.035 18.350 ;
        RECT 95.155 10.310 95.325 18.350 ;
        RECT 97.445 10.310 97.615 18.350 ;
        RECT 92.865 9.450 97.615 10.310 ;
        RECT 98.175 9.450 98.345 19.210 ;
        RECT 99.135 18.520 101.135 18.690 ;
        RECT 101.425 18.520 103.425 18.690 ;
        RECT 98.905 10.310 99.075 18.350 ;
        RECT 101.195 10.310 101.365 18.350 ;
        RECT 103.485 10.310 103.655 18.350 ;
        RECT 98.905 9.450 103.655 10.310 ;
        RECT 104.215 9.450 104.385 19.210 ;
        RECT 105.175 18.520 107.175 18.690 ;
        RECT 107.465 18.520 109.465 18.690 ;
        RECT 104.945 10.310 105.115 18.350 ;
        RECT 107.235 10.310 107.405 18.350 ;
        RECT 109.525 10.310 109.695 18.350 ;
        RECT 104.945 9.450 109.695 10.310 ;
        RECT 110.255 9.450 110.425 19.210 ;
        RECT 111.215 18.520 113.215 18.690 ;
        RECT 113.505 18.520 115.505 18.690 ;
        RECT 110.985 10.310 111.155 18.350 ;
        RECT 113.275 10.310 113.445 18.350 ;
        RECT 115.565 10.310 115.735 18.350 ;
        RECT 110.985 9.450 115.735 10.310 ;
        RECT 116.295 9.450 116.465 19.210 ;
        RECT 117.255 18.520 119.255 18.690 ;
        RECT 119.545 18.520 121.545 18.690 ;
        RECT 117.025 10.310 117.195 18.350 ;
        RECT 119.315 10.310 119.485 18.350 ;
        RECT 121.605 10.310 121.775 18.350 ;
        RECT 117.025 9.450 121.775 10.310 ;
        RECT 122.335 9.450 122.505 19.210 ;
        RECT 123.295 18.520 125.295 18.690 ;
        RECT 125.585 18.520 127.585 18.690 ;
        RECT 123.065 10.310 123.235 18.350 ;
        RECT 125.355 10.310 125.525 18.350 ;
        RECT 127.645 10.310 127.815 18.350 ;
        RECT 123.065 9.450 127.815 10.310 ;
        RECT 128.375 9.450 128.905 19.210 ;
        RECT 135.150 18.895 135.680 104.785 ;
        RECT 136.265 103.615 138.425 104.305 ;
        RECT 136.265 102.445 138.425 103.135 ;
        RECT 136.265 101.275 138.425 101.965 ;
        RECT 136.265 100.105 138.425 100.795 ;
        RECT 136.265 98.935 138.425 99.625 ;
        RECT 136.265 97.765 138.425 98.455 ;
        RECT 136.265 96.595 138.425 97.285 ;
        RECT 136.265 95.425 138.425 96.115 ;
        RECT 136.265 94.255 138.425 94.945 ;
        RECT 136.265 93.085 138.425 93.775 ;
        RECT 136.265 91.915 138.425 92.605 ;
        RECT 136.265 90.745 138.425 91.435 ;
        RECT 136.265 89.575 138.425 90.265 ;
        RECT 136.265 88.405 138.425 89.095 ;
        RECT 136.265 87.235 138.425 87.925 ;
        RECT 136.265 86.065 138.425 86.755 ;
        RECT 136.265 84.895 138.425 85.585 ;
        RECT 136.265 83.725 138.425 84.415 ;
        RECT 136.265 82.555 138.425 83.245 ;
        RECT 136.265 81.385 138.425 82.075 ;
        RECT 136.265 80.215 138.425 80.905 ;
        RECT 136.265 79.045 138.425 79.735 ;
        RECT 136.265 77.875 138.425 78.565 ;
        RECT 136.265 76.705 138.425 77.395 ;
        RECT 136.265 75.535 138.425 76.225 ;
        RECT 136.265 74.365 138.425 75.055 ;
        RECT 136.265 73.195 138.425 73.885 ;
        RECT 136.265 72.025 138.425 72.715 ;
        RECT 136.265 70.855 138.425 71.545 ;
        RECT 136.265 69.685 138.425 70.375 ;
        RECT 136.265 68.515 138.425 69.205 ;
        RECT 136.265 67.345 138.425 68.035 ;
        RECT 136.265 66.175 138.425 66.865 ;
        RECT 136.265 65.005 138.425 65.695 ;
        RECT 136.265 63.835 138.425 64.525 ;
        RECT 136.265 62.665 138.425 63.355 ;
        RECT 136.265 61.495 138.425 62.185 ;
        RECT 136.265 60.325 138.425 61.015 ;
        RECT 136.265 59.155 138.425 59.845 ;
        RECT 136.265 57.985 138.425 58.675 ;
        RECT 136.265 56.815 138.425 57.505 ;
        RECT 136.265 55.645 138.425 56.335 ;
        RECT 136.265 54.475 138.425 55.165 ;
        RECT 136.265 53.305 138.425 53.995 ;
        RECT 136.265 52.135 138.425 52.825 ;
        RECT 136.265 50.965 138.425 51.655 ;
        RECT 136.265 49.795 138.425 50.485 ;
        RECT 136.265 48.625 138.425 49.315 ;
        RECT 136.265 47.455 138.425 48.145 ;
        RECT 136.265 46.285 138.425 46.975 ;
        RECT 136.265 45.115 138.425 45.805 ;
        RECT 136.265 43.945 138.425 44.635 ;
        RECT 136.265 42.775 138.425 43.465 ;
        RECT 136.265 41.605 138.425 42.295 ;
        RECT 136.265 40.435 138.425 41.125 ;
        RECT 136.265 39.265 138.425 39.955 ;
        RECT 136.265 38.095 138.425 38.785 ;
        RECT 136.265 36.925 138.425 37.615 ;
        RECT 136.265 35.755 138.425 36.445 ;
        RECT 136.265 34.585 138.425 35.275 ;
        RECT 136.265 33.415 138.425 34.105 ;
        RECT 136.265 32.245 138.425 32.935 ;
        RECT 136.265 31.075 138.425 31.765 ;
        RECT 136.265 29.905 138.425 30.595 ;
        RECT 136.265 28.735 138.425 29.425 ;
        RECT 136.265 27.565 138.425 28.255 ;
        RECT 136.265 26.395 138.425 27.085 ;
        RECT 136.265 25.225 138.425 25.915 ;
        RECT 136.265 24.055 138.425 24.745 ;
        RECT 136.265 22.885 138.425 23.575 ;
        RECT 136.265 21.715 138.425 22.405 ;
        RECT 136.265 20.545 138.425 21.235 ;
        RECT 136.265 19.375 138.425 20.065 ;
        RECT 139.150 18.895 145.540 104.785 ;
        RECT 146.265 103.615 148.425 104.305 ;
        RECT 146.265 102.445 148.425 103.135 ;
        RECT 146.265 101.275 148.425 101.965 ;
        RECT 146.265 100.105 148.425 100.795 ;
        RECT 146.265 98.935 148.425 99.625 ;
        RECT 146.265 97.765 148.425 98.455 ;
        RECT 146.265 96.595 148.425 97.285 ;
        RECT 146.265 95.425 148.425 96.115 ;
        RECT 146.265 94.255 148.425 94.945 ;
        RECT 146.265 93.085 148.425 93.775 ;
        RECT 146.265 91.915 148.425 92.605 ;
        RECT 146.265 90.745 148.425 91.435 ;
        RECT 146.265 89.575 148.425 90.265 ;
        RECT 146.265 88.405 148.425 89.095 ;
        RECT 146.265 87.235 148.425 87.925 ;
        RECT 146.265 86.065 148.425 86.755 ;
        RECT 146.265 84.895 148.425 85.585 ;
        RECT 146.265 83.725 148.425 84.415 ;
        RECT 146.265 82.555 148.425 83.245 ;
        RECT 146.265 81.385 148.425 82.075 ;
        RECT 146.265 80.215 148.425 80.905 ;
        RECT 146.265 79.045 148.425 79.735 ;
        RECT 146.265 77.875 148.425 78.565 ;
        RECT 146.265 76.705 148.425 77.395 ;
        RECT 146.265 75.535 148.425 76.225 ;
        RECT 146.265 74.365 148.425 75.055 ;
        RECT 146.265 73.195 148.425 73.885 ;
        RECT 146.265 72.025 148.425 72.715 ;
        RECT 146.265 70.855 148.425 71.545 ;
        RECT 146.265 69.685 148.425 70.375 ;
        RECT 146.265 68.515 148.425 69.205 ;
        RECT 146.265 67.345 148.425 68.035 ;
        RECT 146.265 66.175 148.425 66.865 ;
        RECT 146.265 65.005 148.425 65.695 ;
        RECT 146.265 63.835 148.425 64.525 ;
        RECT 146.265 62.665 148.425 63.355 ;
        RECT 146.265 61.495 148.425 62.185 ;
        RECT 146.265 60.325 148.425 61.015 ;
        RECT 146.265 59.155 148.425 59.845 ;
        RECT 146.265 57.985 148.425 58.675 ;
        RECT 146.265 56.815 148.425 57.505 ;
        RECT 146.265 55.645 148.425 56.335 ;
        RECT 146.265 54.475 148.425 55.165 ;
        RECT 146.265 53.305 148.425 53.995 ;
        RECT 146.265 52.135 148.425 52.825 ;
        RECT 146.265 50.965 148.425 51.655 ;
        RECT 146.265 49.795 148.425 50.485 ;
        RECT 146.265 48.625 148.425 49.315 ;
        RECT 146.265 47.455 148.425 48.145 ;
        RECT 146.265 46.285 148.425 46.975 ;
        RECT 146.265 45.115 148.425 45.805 ;
        RECT 146.265 43.945 148.425 44.635 ;
        RECT 146.265 42.775 148.425 43.465 ;
        RECT 146.265 41.605 148.425 42.295 ;
        RECT 146.265 40.435 148.425 41.125 ;
        RECT 146.265 39.265 148.425 39.955 ;
        RECT 146.265 38.095 148.425 38.785 ;
        RECT 146.265 36.925 148.425 37.615 ;
        RECT 146.265 35.755 148.425 36.445 ;
        RECT 146.265 34.585 148.425 35.275 ;
        RECT 146.265 33.415 148.425 34.105 ;
        RECT 146.265 32.245 148.425 32.935 ;
        RECT 146.265 31.075 148.425 31.765 ;
        RECT 146.265 29.905 148.425 30.595 ;
        RECT 146.265 28.735 148.425 29.425 ;
        RECT 146.265 27.565 148.425 28.255 ;
        RECT 146.265 26.395 148.425 27.085 ;
        RECT 146.265 25.225 148.425 25.915 ;
        RECT 146.265 24.055 148.425 24.745 ;
        RECT 146.265 22.885 148.425 23.575 ;
        RECT 146.265 21.715 148.425 22.405 ;
        RECT 146.265 20.545 148.425 21.235 ;
        RECT 146.265 19.375 148.425 20.065 ;
        RECT 149.010 18.895 149.540 104.785 ;
        RECT 135.150 13.490 149.540 18.895 ;
        RECT 79.695 8.920 128.905 9.450 ;
        RECT 155.300 4.700 155.700 180.620 ;
        RECT 162.180 179.815 163.390 180.905 ;
        RECT 164.695 179.815 165.025 180.915 ;
        RECT 165.500 180.585 166.205 180.995 ;
        RECT 166.375 181.625 166.915 181.795 ;
        RECT 167.195 181.625 167.365 182.365 ;
        RECT 167.760 182.000 167.930 182.025 ;
        RECT 167.630 181.625 167.990 182.000 ;
        RECT 166.375 180.925 166.545 181.625 ;
        RECT 166.715 181.125 167.045 181.455 ;
        RECT 167.215 181.125 167.565 181.455 ;
        RECT 166.375 180.755 167.000 180.925 ;
        RECT 167.215 180.585 167.480 181.125 ;
        RECT 167.735 180.970 167.990 181.625 ;
        RECT 168.315 181.715 168.645 182.180 ;
        RECT 168.815 181.895 168.985 182.365 ;
        RECT 169.155 181.715 169.485 182.195 ;
        RECT 168.315 181.545 169.485 181.715 ;
        RECT 168.160 181.165 168.805 181.375 ;
        RECT 168.975 181.165 169.545 181.375 ;
        RECT 169.715 180.995 169.885 182.195 ;
        RECT 170.425 181.795 170.595 182.000 ;
        RECT 165.500 180.415 167.480 180.585 ;
        RECT 165.500 179.985 165.825 180.415 ;
        RECT 165.995 179.815 166.325 180.235 ;
        RECT 167.070 179.815 167.480 180.245 ;
        RECT 167.650 179.985 167.990 180.970 ;
        RECT 168.375 179.815 168.705 180.915 ;
        RECT 169.180 180.585 169.885 180.995 ;
        RECT 170.055 181.625 170.595 181.795 ;
        RECT 170.875 181.625 171.045 182.365 ;
        RECT 171.440 182.000 171.610 182.025 ;
        RECT 171.310 181.625 171.670 182.000 ;
        RECT 170.055 180.925 170.225 181.625 ;
        RECT 170.395 181.125 170.725 181.455 ;
        RECT 170.895 181.125 171.245 181.455 ;
        RECT 170.055 180.755 170.680 180.925 ;
        RECT 170.895 180.585 171.160 181.125 ;
        RECT 171.415 180.970 171.670 181.625 ;
        RECT 171.995 181.715 172.325 182.180 ;
        RECT 172.495 181.895 172.665 182.365 ;
        RECT 172.835 181.715 173.165 182.195 ;
        RECT 171.995 181.545 173.165 181.715 ;
        RECT 171.840 181.165 172.485 181.375 ;
        RECT 172.655 181.165 173.225 181.375 ;
        RECT 173.395 180.995 173.565 182.195 ;
        RECT 174.105 181.795 174.275 182.000 ;
        RECT 169.180 180.415 171.160 180.585 ;
        RECT 169.180 179.985 169.505 180.415 ;
        RECT 169.675 179.815 170.005 180.235 ;
        RECT 170.750 179.815 171.160 180.245 ;
        RECT 171.330 179.985 171.670 180.970 ;
        RECT 172.055 179.815 172.385 180.915 ;
        RECT 172.860 180.585 173.565 180.995 ;
        RECT 173.735 181.625 174.275 181.795 ;
        RECT 174.555 181.625 174.725 182.365 ;
        RECT 174.990 181.625 175.350 182.000 ;
        RECT 173.735 180.925 173.905 181.625 ;
        RECT 174.075 181.125 174.405 181.455 ;
        RECT 174.575 181.125 174.925 181.455 ;
        RECT 173.735 180.755 174.360 180.925 ;
        RECT 174.575 180.585 174.840 181.125 ;
        RECT 175.095 180.970 175.350 181.625 ;
        RECT 175.675 181.715 176.005 182.180 ;
        RECT 176.175 181.895 176.345 182.365 ;
        RECT 176.515 181.715 176.845 182.195 ;
        RECT 175.675 181.545 176.845 181.715 ;
        RECT 175.520 181.165 176.165 181.375 ;
        RECT 176.335 181.165 176.905 181.375 ;
        RECT 177.075 180.995 177.245 182.195 ;
        RECT 177.785 181.795 177.955 182.000 ;
        RECT 172.860 180.415 174.840 180.585 ;
        RECT 172.860 179.985 173.185 180.415 ;
        RECT 173.355 179.815 173.685 180.235 ;
        RECT 174.430 179.815 174.840 180.245 ;
        RECT 175.010 179.985 175.350 180.970 ;
        RECT 175.735 179.815 176.065 180.915 ;
        RECT 176.540 180.585 177.245 180.995 ;
        RECT 177.415 181.625 177.955 181.795 ;
        RECT 178.235 181.625 178.405 182.365 ;
        RECT 178.670 181.625 179.030 182.000 ;
        RECT 177.415 180.925 177.585 181.625 ;
        RECT 177.755 181.125 178.085 181.455 ;
        RECT 178.255 181.125 178.605 181.455 ;
        RECT 177.415 180.755 178.040 180.925 ;
        RECT 178.255 180.585 178.520 181.125 ;
        RECT 178.775 180.970 179.030 181.625 ;
        RECT 176.540 180.415 178.520 180.585 ;
        RECT 176.540 179.985 176.865 180.415 ;
        RECT 177.035 179.815 177.365 180.235 ;
        RECT 178.110 179.815 178.520 180.245 ;
        RECT 178.690 179.985 179.030 180.970 ;
        RECT 179.665 181.625 179.920 182.195 ;
        RECT 180.090 181.965 180.420 182.365 ;
        RECT 180.845 181.830 181.375 182.195 ;
        RECT 181.565 182.025 181.840 182.195 ;
        RECT 181.560 181.855 181.840 182.025 ;
        RECT 180.845 181.795 181.020 181.830 ;
        RECT 180.090 181.625 181.020 181.795 ;
        RECT 179.665 180.955 179.835 181.625 ;
        RECT 180.090 181.455 180.260 181.625 ;
        RECT 180.005 181.125 180.260 181.455 ;
        RECT 180.485 181.125 180.680 181.455 ;
        RECT 179.665 179.985 180.000 180.955 ;
        RECT 180.170 179.815 180.340 180.955 ;
        RECT 180.510 180.155 180.680 181.125 ;
        RECT 180.850 180.495 181.020 181.625 ;
        RECT 181.190 180.835 181.360 181.635 ;
        RECT 181.565 181.035 181.840 181.855 ;
        RECT 182.010 180.835 182.200 182.195 ;
        RECT 182.380 181.830 182.890 182.365 ;
        RECT 183.110 181.555 183.355 182.160 ;
        RECT 183.805 181.625 184.060 182.195 ;
        RECT 184.230 181.965 184.560 182.365 ;
        RECT 184.985 181.830 185.515 182.195 ;
        RECT 185.705 182.025 185.980 182.195 ;
        RECT 185.700 181.855 185.980 182.025 ;
        RECT 184.985 181.795 185.160 181.830 ;
        RECT 184.230 181.625 185.160 181.795 ;
        RECT 182.400 181.385 183.630 181.555 ;
        RECT 181.190 180.665 182.200 180.835 ;
        RECT 182.370 180.820 183.120 181.010 ;
        RECT 180.850 180.325 181.975 180.495 ;
        RECT 182.370 180.155 182.540 180.820 ;
        RECT 183.290 180.575 183.630 181.385 ;
        RECT 180.510 179.985 182.540 180.155 ;
        RECT 182.710 179.815 182.880 180.575 ;
        RECT 183.115 180.165 183.630 180.575 ;
        RECT 183.805 180.955 183.975 181.625 ;
        RECT 184.230 181.455 184.400 181.625 ;
        RECT 184.145 181.125 184.400 181.455 ;
        RECT 184.625 181.125 184.820 181.455 ;
        RECT 183.805 179.985 184.140 180.955 ;
        RECT 184.310 179.815 184.480 180.955 ;
        RECT 184.650 180.155 184.820 181.125 ;
        RECT 184.990 180.495 185.160 181.625 ;
        RECT 185.330 180.835 185.500 181.635 ;
        RECT 185.705 181.035 185.980 181.855 ;
        RECT 186.150 180.835 186.340 182.195 ;
        RECT 186.520 181.830 187.030 182.365 ;
        RECT 187.250 181.555 187.495 182.160 ;
        RECT 187.940 181.640 188.230 182.365 ;
        RECT 188.865 181.625 189.120 182.195 ;
        RECT 189.290 181.965 189.620 182.365 ;
        RECT 190.045 181.830 190.575 182.195 ;
        RECT 190.045 181.795 190.220 181.830 ;
        RECT 189.290 181.625 190.220 181.795 ;
        RECT 190.765 181.685 191.040 182.195 ;
        RECT 186.540 181.385 187.770 181.555 ;
        RECT 185.330 180.665 186.340 180.835 ;
        RECT 186.510 180.820 187.260 181.010 ;
        RECT 184.990 180.325 186.115 180.495 ;
        RECT 186.510 180.155 186.680 180.820 ;
        RECT 187.430 180.575 187.770 181.385 ;
        RECT 184.650 179.985 186.680 180.155 ;
        RECT 186.850 179.815 187.020 180.575 ;
        RECT 187.255 180.165 187.770 180.575 ;
        RECT 187.940 179.815 188.230 180.980 ;
        RECT 188.865 180.955 189.035 181.625 ;
        RECT 189.290 181.455 189.460 181.625 ;
        RECT 189.205 181.125 189.460 181.455 ;
        RECT 189.685 181.125 189.880 181.455 ;
        RECT 188.865 179.985 189.200 180.955 ;
        RECT 189.370 179.815 189.540 180.955 ;
        RECT 189.710 180.155 189.880 181.125 ;
        RECT 190.050 180.495 190.220 181.625 ;
        RECT 190.390 180.835 190.560 181.635 ;
        RECT 190.760 181.515 191.040 181.685 ;
        RECT 190.765 181.035 191.040 181.515 ;
        RECT 191.210 180.835 191.400 182.195 ;
        RECT 191.580 181.830 192.090 182.365 ;
        RECT 192.310 181.555 192.555 182.160 ;
        RECT 193.465 181.625 193.720 182.195 ;
        RECT 193.890 181.965 194.220 182.365 ;
        RECT 194.645 181.830 195.175 182.195 ;
        RECT 194.645 181.795 194.820 181.830 ;
        RECT 193.890 181.625 194.820 181.795 ;
        RECT 191.600 181.385 192.830 181.555 ;
        RECT 190.390 180.665 191.400 180.835 ;
        RECT 191.570 180.820 192.320 181.010 ;
        RECT 190.050 180.325 191.175 180.495 ;
        RECT 191.570 180.155 191.740 180.820 ;
        RECT 192.490 180.575 192.830 181.385 ;
        RECT 189.710 179.985 191.740 180.155 ;
        RECT 191.910 179.815 192.080 180.575 ;
        RECT 192.315 180.165 192.830 180.575 ;
        RECT 193.465 180.955 193.635 181.625 ;
        RECT 193.890 181.455 194.060 181.625 ;
        RECT 193.805 181.125 194.060 181.455 ;
        RECT 194.285 181.125 194.480 181.455 ;
        RECT 193.465 179.985 193.800 180.955 ;
        RECT 193.970 179.815 194.140 180.955 ;
        RECT 194.310 180.155 194.480 181.125 ;
        RECT 194.650 180.495 194.820 181.625 ;
        RECT 194.990 180.835 195.160 181.635 ;
        RECT 195.365 181.345 195.640 182.195 ;
        RECT 195.360 181.175 195.640 181.345 ;
        RECT 195.365 181.035 195.640 181.175 ;
        RECT 195.810 180.835 196.000 182.195 ;
        RECT 196.180 181.830 196.690 182.365 ;
        RECT 196.910 181.555 197.155 182.160 ;
        RECT 198.520 181.690 198.780 182.195 ;
        RECT 198.960 181.985 199.290 182.365 ;
        RECT 199.470 181.815 199.640 182.195 ;
        RECT 196.200 181.385 197.430 181.555 ;
        RECT 194.990 180.665 196.000 180.835 ;
        RECT 196.170 180.820 196.920 181.010 ;
        RECT 194.650 180.325 195.775 180.495 ;
        RECT 196.170 180.155 196.340 180.820 ;
        RECT 197.090 180.575 197.430 181.385 ;
        RECT 194.310 179.985 196.340 180.155 ;
        RECT 196.510 179.815 196.680 180.575 ;
        RECT 196.915 180.165 197.430 180.575 ;
        RECT 198.520 180.890 198.690 181.690 ;
        RECT 198.975 181.645 199.640 181.815 ;
        RECT 199.990 181.815 200.160 182.195 ;
        RECT 200.340 181.985 200.670 182.365 ;
        RECT 199.990 181.645 200.655 181.815 ;
        RECT 200.850 181.690 201.110 182.195 ;
        RECT 198.975 181.390 199.145 181.645 ;
        RECT 198.860 181.060 199.145 181.390 ;
        RECT 199.380 181.095 199.710 181.465 ;
        RECT 199.920 181.095 200.250 181.465 ;
        RECT 200.485 181.390 200.655 181.645 ;
        RECT 198.975 180.915 199.145 181.060 ;
        RECT 200.485 181.060 200.770 181.390 ;
        RECT 200.485 180.915 200.655 181.060 ;
        RECT 198.520 179.985 198.790 180.890 ;
        RECT 198.975 180.745 199.640 180.915 ;
        RECT 198.960 179.815 199.290 180.575 ;
        RECT 199.470 179.985 199.640 180.745 ;
        RECT 199.990 180.745 200.655 180.915 ;
        RECT 200.940 180.890 201.110 181.690 ;
        RECT 201.370 181.815 201.540 182.195 ;
        RECT 201.720 181.985 202.050 182.365 ;
        RECT 201.370 181.645 202.035 181.815 ;
        RECT 202.230 181.690 202.490 182.195 ;
        RECT 201.300 181.095 201.630 181.465 ;
        RECT 201.865 181.390 202.035 181.645 ;
        RECT 201.865 181.060 202.150 181.390 ;
        RECT 201.865 180.915 202.035 181.060 ;
        RECT 199.990 179.985 200.160 180.745 ;
        RECT 200.340 179.815 200.670 180.575 ;
        RECT 200.840 179.985 201.110 180.890 ;
        RECT 201.370 180.745 202.035 180.915 ;
        RECT 202.320 180.890 202.490 181.690 ;
        RECT 202.750 181.815 202.920 182.195 ;
        RECT 203.100 181.985 203.430 182.365 ;
        RECT 202.750 181.645 203.415 181.815 ;
        RECT 203.610 181.690 203.870 182.195 ;
        RECT 202.680 181.095 203.010 181.465 ;
        RECT 203.245 181.390 203.415 181.645 ;
        RECT 203.245 181.060 203.530 181.390 ;
        RECT 203.245 180.915 203.415 181.060 ;
        RECT 201.370 179.985 201.540 180.745 ;
        RECT 201.720 179.815 202.050 180.575 ;
        RECT 202.220 179.985 202.490 180.890 ;
        RECT 202.750 180.745 203.415 180.915 ;
        RECT 203.700 180.890 203.870 181.690 ;
        RECT 204.130 181.815 204.300 182.190 ;
        RECT 204.470 181.985 204.800 182.365 ;
        RECT 204.970 182.025 206.045 182.195 ;
        RECT 204.970 181.815 205.140 182.025 ;
        RECT 204.130 181.645 205.140 181.815 ;
        RECT 205.365 181.685 205.705 181.855 ;
        RECT 205.875 181.690 206.045 182.025 ;
        RECT 205.365 181.515 205.655 181.685 ;
        RECT 204.105 181.345 204.450 181.455 ;
        RECT 204.100 181.175 204.450 181.345 ;
        RECT 202.750 179.985 202.920 180.745 ;
        RECT 203.100 179.815 203.430 180.575 ;
        RECT 203.600 179.985 203.870 180.890 ;
        RECT 204.105 180.835 204.450 181.175 ;
        RECT 204.760 180.835 205.195 181.455 ;
        RECT 205.365 180.995 205.535 181.515 ;
        RECT 206.215 181.345 206.575 182.020 ;
        RECT 206.755 181.645 207.045 182.365 ;
        RECT 207.335 182.025 208.935 182.195 ;
        RECT 207.335 181.655 207.505 182.025 ;
        RECT 208.580 181.985 208.935 182.025 ;
        RECT 209.105 181.905 209.275 182.365 ;
        RECT 207.675 181.605 208.005 181.855 ;
        RECT 207.690 181.530 208.005 181.605 ;
        RECT 208.175 181.735 208.345 181.855 ;
        RECT 209.450 181.735 209.695 182.155 ;
        RECT 209.965 181.985 210.295 182.365 ;
        RECT 210.465 181.795 210.640 182.125 ;
        RECT 210.985 182.035 211.155 182.195 ;
        RECT 210.985 181.865 211.515 182.035 ;
        RECT 211.685 182.025 212.680 182.195 ;
        RECT 211.685 181.865 211.855 182.025 ;
        RECT 208.175 181.565 209.695 181.735 ;
        RECT 206.035 181.165 206.575 181.345 ;
        RECT 206.215 181.055 206.575 181.165 ;
        RECT 205.365 180.825 206.000 180.995 ;
        RECT 206.215 180.825 207.020 181.055 ;
        RECT 204.130 180.485 205.660 180.655 ;
        RECT 204.130 179.985 204.300 180.485 ;
        RECT 205.490 180.325 205.660 180.485 ;
        RECT 205.830 180.495 206.000 180.825 ;
        RECT 205.830 180.325 206.160 180.495 ;
        RECT 204.470 179.815 204.800 180.195 ;
        RECT 204.970 180.155 205.140 180.315 ;
        RECT 206.330 180.155 206.500 180.655 ;
        RECT 204.970 179.985 206.500 180.155 ;
        RECT 206.670 179.985 207.020 180.825 ;
        RECT 207.220 180.455 207.520 181.455 ;
        RECT 207.690 181.005 207.860 181.530 ;
        RECT 208.175 181.525 208.345 181.565 ;
        RECT 208.030 181.345 208.360 181.355 ;
        RECT 208.755 181.345 209.000 181.395 ;
        RECT 208.030 181.185 208.415 181.345 ;
        RECT 208.245 181.175 208.415 181.185 ;
        RECT 208.700 181.175 209.000 181.345 ;
        RECT 207.690 180.835 208.450 181.005 ;
        RECT 207.190 179.815 207.520 180.195 ;
        RECT 207.780 180.155 207.950 180.665 ;
        RECT 208.120 180.325 208.450 180.835 ;
        RECT 208.755 180.775 209.000 181.175 ;
        RECT 209.205 181.345 209.535 181.395 ;
        RECT 209.205 181.175 209.560 181.345 ;
        RECT 209.205 180.775 209.535 181.175 ;
        RECT 210.010 180.775 210.300 181.455 ;
        RECT 210.470 181.345 210.640 181.795 ;
        RECT 210.935 181.515 211.175 181.685 ;
        RECT 210.470 181.175 210.760 181.345 ;
        RECT 208.620 180.365 209.685 180.535 ;
        RECT 208.620 180.155 208.790 180.365 ;
        RECT 207.780 179.985 208.790 180.155 ;
        RECT 209.015 179.815 209.345 180.195 ;
        RECT 209.515 179.985 209.685 180.365 ;
        RECT 210.470 180.315 210.640 181.175 ;
        RECT 209.935 179.815 210.285 180.195 ;
        RECT 210.455 179.985 210.640 180.315 ;
        RECT 210.935 180.315 211.105 181.515 ;
        RECT 211.345 180.695 211.515 181.865 ;
        RECT 212.165 181.685 212.340 181.855 ;
        RECT 211.925 181.525 212.340 181.685 ;
        RECT 212.510 181.735 212.680 182.025 ;
        RECT 212.850 181.905 213.020 182.365 ;
        RECT 212.510 181.565 213.080 181.735 ;
        RECT 211.925 181.515 212.335 181.525 ;
        RECT 212.145 181.175 212.600 181.345 ;
        RECT 212.910 180.785 213.080 181.565 ;
        RECT 211.345 180.465 212.130 180.695 ;
        RECT 211.800 180.325 212.130 180.465 ;
        RECT 212.430 180.615 213.080 180.785 ;
        RECT 210.935 179.985 211.145 180.315 ;
        RECT 211.315 180.155 211.645 180.195 ;
        RECT 212.430 180.155 212.600 180.615 ;
        RECT 211.315 179.985 212.600 180.155 ;
        RECT 212.770 179.815 213.100 180.195 ;
        RECT 213.270 179.985 213.530 182.195 ;
        RECT 213.700 181.640 213.990 182.365 ;
        RECT 214.250 181.815 214.420 182.190 ;
        RECT 214.590 181.985 214.920 182.365 ;
        RECT 215.090 182.025 216.165 182.195 ;
        RECT 215.090 181.815 215.260 182.025 ;
        RECT 214.250 181.645 215.260 181.815 ;
        RECT 215.485 181.685 215.825 181.855 ;
        RECT 215.995 181.690 216.165 182.025 ;
        RECT 215.485 181.515 215.775 181.685 ;
        RECT 214.225 181.345 214.570 181.455 ;
        RECT 214.220 181.175 214.570 181.345 ;
        RECT 213.700 179.815 213.990 180.980 ;
        RECT 214.225 180.835 214.570 181.175 ;
        RECT 214.880 180.835 215.315 181.455 ;
        RECT 215.485 180.995 215.655 181.515 ;
        RECT 216.335 181.345 216.695 182.020 ;
        RECT 216.875 181.645 217.165 182.365 ;
        RECT 217.455 182.025 219.055 182.195 ;
        RECT 217.455 181.655 217.625 182.025 ;
        RECT 218.700 181.985 219.055 182.025 ;
        RECT 219.225 181.905 219.395 182.365 ;
        RECT 217.795 181.605 218.125 181.855 ;
        RECT 217.810 181.530 218.125 181.605 ;
        RECT 218.295 181.735 218.465 181.855 ;
        RECT 219.570 181.735 219.815 182.155 ;
        RECT 220.085 181.985 220.415 182.365 ;
        RECT 220.585 181.795 220.760 182.125 ;
        RECT 221.105 182.035 221.275 182.195 ;
        RECT 221.105 181.865 221.635 182.035 ;
        RECT 221.805 182.025 222.800 182.195 ;
        RECT 221.805 181.865 221.975 182.025 ;
        RECT 218.295 181.565 219.815 181.735 ;
        RECT 216.155 181.165 216.695 181.345 ;
        RECT 216.335 181.055 216.695 181.165 ;
        RECT 215.485 180.825 216.120 180.995 ;
        RECT 216.335 180.825 217.140 181.055 ;
        RECT 214.250 180.485 215.780 180.655 ;
        RECT 214.250 179.985 214.420 180.485 ;
        RECT 215.610 180.325 215.780 180.485 ;
        RECT 215.950 180.495 216.120 180.825 ;
        RECT 215.950 180.325 216.280 180.495 ;
        RECT 214.590 179.815 214.920 180.195 ;
        RECT 215.090 180.155 215.260 180.315 ;
        RECT 216.450 180.155 216.620 180.655 ;
        RECT 215.090 179.985 216.620 180.155 ;
        RECT 216.790 179.985 217.140 180.825 ;
        RECT 217.340 180.455 217.640 181.455 ;
        RECT 217.810 181.005 217.980 181.530 ;
        RECT 218.295 181.525 218.465 181.565 ;
        RECT 218.150 181.345 218.480 181.355 ;
        RECT 218.150 181.185 218.535 181.345 ;
        RECT 218.365 181.175 218.535 181.185 ;
        RECT 218.875 181.005 219.120 181.395 ;
        RECT 217.810 180.835 218.570 181.005 ;
        RECT 218.820 180.835 219.120 181.005 ;
        RECT 217.310 179.815 217.640 180.195 ;
        RECT 217.900 180.155 218.070 180.665 ;
        RECT 218.240 180.325 218.570 180.835 ;
        RECT 218.875 180.775 219.120 180.835 ;
        RECT 219.325 181.005 219.655 181.395 ;
        RECT 219.325 180.835 219.680 181.005 ;
        RECT 219.325 180.775 219.655 180.835 ;
        RECT 220.130 180.775 220.420 181.455 ;
        RECT 220.590 181.345 220.760 181.795 ;
        RECT 221.055 181.515 221.295 181.685 ;
        RECT 220.590 181.175 220.880 181.345 ;
        RECT 218.740 180.365 219.805 180.535 ;
        RECT 218.740 180.155 218.910 180.365 ;
        RECT 217.900 179.985 218.910 180.155 ;
        RECT 219.135 179.815 219.465 180.195 ;
        RECT 219.635 179.985 219.805 180.365 ;
        RECT 220.590 180.315 220.760 181.175 ;
        RECT 220.055 179.815 220.405 180.195 ;
        RECT 220.575 179.985 220.760 180.315 ;
        RECT 221.055 180.315 221.225 181.515 ;
        RECT 221.465 180.695 221.635 181.865 ;
        RECT 222.285 181.685 222.460 181.855 ;
        RECT 222.045 181.525 222.460 181.685 ;
        RECT 222.630 181.735 222.800 182.025 ;
        RECT 222.970 181.905 223.140 182.365 ;
        RECT 222.630 181.565 223.200 181.735 ;
        RECT 222.045 181.515 222.455 181.525 ;
        RECT 222.265 181.175 222.720 181.345 ;
        RECT 223.030 180.785 223.200 181.565 ;
        RECT 221.465 180.465 222.250 180.695 ;
        RECT 221.920 180.325 222.250 180.465 ;
        RECT 222.550 180.615 223.200 180.785 ;
        RECT 221.055 179.985 221.265 180.315 ;
        RECT 221.435 180.155 221.765 180.195 ;
        RECT 222.550 180.155 222.720 180.615 ;
        RECT 221.435 179.985 222.720 180.155 ;
        RECT 222.890 179.815 223.220 180.195 ;
        RECT 223.390 179.985 223.650 182.195 ;
        RECT 223.910 181.815 224.080 182.190 ;
        RECT 224.250 181.985 224.580 182.365 ;
        RECT 224.750 182.025 225.825 182.195 ;
        RECT 224.750 181.815 224.920 182.025 ;
        RECT 223.910 181.645 224.920 181.815 ;
        RECT 225.145 181.685 225.485 181.855 ;
        RECT 225.655 181.690 225.825 182.025 ;
        RECT 225.145 181.515 225.435 181.685 ;
        RECT 223.885 181.345 224.230 181.455 ;
        RECT 223.880 181.175 224.230 181.345 ;
        RECT 223.885 180.835 224.230 181.175 ;
        RECT 224.540 180.835 224.975 181.455 ;
        RECT 225.145 180.995 225.315 181.515 ;
        RECT 225.995 181.345 226.355 182.020 ;
        RECT 226.535 181.645 226.825 182.365 ;
        RECT 227.115 182.025 228.715 182.195 ;
        RECT 227.115 181.655 227.285 182.025 ;
        RECT 228.360 181.985 228.715 182.025 ;
        RECT 228.885 181.905 229.055 182.365 ;
        RECT 227.455 181.605 227.785 181.855 ;
        RECT 227.470 181.530 227.785 181.605 ;
        RECT 227.955 181.735 228.125 181.855 ;
        RECT 229.230 181.735 229.475 182.155 ;
        RECT 229.745 181.985 230.075 182.365 ;
        RECT 230.245 181.795 230.420 182.125 ;
        RECT 230.765 182.035 230.935 182.195 ;
        RECT 230.765 181.865 231.295 182.035 ;
        RECT 231.465 182.025 232.460 182.195 ;
        RECT 231.465 181.865 231.635 182.025 ;
        RECT 227.955 181.565 229.475 181.735 ;
        RECT 225.815 181.165 226.355 181.345 ;
        RECT 225.995 181.055 226.355 181.165 ;
        RECT 225.145 180.825 225.780 180.995 ;
        RECT 225.995 180.825 226.800 181.055 ;
        RECT 223.910 180.485 225.440 180.655 ;
        RECT 223.910 179.985 224.080 180.485 ;
        RECT 225.270 180.325 225.440 180.485 ;
        RECT 225.610 180.495 225.780 180.825 ;
        RECT 225.610 180.325 225.940 180.495 ;
        RECT 224.250 179.815 224.580 180.195 ;
        RECT 224.750 180.155 224.920 180.315 ;
        RECT 226.110 180.155 226.280 180.655 ;
        RECT 224.750 179.985 226.280 180.155 ;
        RECT 226.450 179.985 226.800 180.825 ;
        RECT 227.000 180.455 227.300 181.455 ;
        RECT 227.470 181.005 227.640 181.530 ;
        RECT 227.955 181.525 228.125 181.565 ;
        RECT 227.810 181.345 228.140 181.355 ;
        RECT 227.810 181.185 228.195 181.345 ;
        RECT 228.025 181.175 228.195 181.185 ;
        RECT 227.470 180.835 228.230 181.005 ;
        RECT 226.970 179.815 227.300 180.195 ;
        RECT 227.560 180.155 227.730 180.665 ;
        RECT 227.900 180.325 228.230 180.835 ;
        RECT 228.535 180.775 228.780 181.395 ;
        RECT 228.985 181.005 229.315 181.395 ;
        RECT 228.985 180.835 229.340 181.005 ;
        RECT 228.985 180.775 229.315 180.835 ;
        RECT 229.790 180.775 230.080 181.455 ;
        RECT 230.250 181.345 230.420 181.795 ;
        RECT 230.715 181.515 230.955 181.685 ;
        RECT 230.250 181.175 230.540 181.345 ;
        RECT 228.400 180.365 229.465 180.535 ;
        RECT 228.400 180.155 228.570 180.365 ;
        RECT 227.560 179.985 228.570 180.155 ;
        RECT 228.795 179.815 229.125 180.195 ;
        RECT 229.295 179.985 229.465 180.365 ;
        RECT 230.250 180.315 230.420 181.175 ;
        RECT 229.715 179.815 230.065 180.195 ;
        RECT 230.235 179.985 230.420 180.315 ;
        RECT 230.715 180.315 230.885 181.515 ;
        RECT 231.125 180.695 231.295 181.865 ;
        RECT 231.945 181.685 232.120 181.855 ;
        RECT 231.705 181.525 232.120 181.685 ;
        RECT 232.290 181.735 232.460 182.025 ;
        RECT 232.630 181.905 232.800 182.365 ;
        RECT 232.290 181.565 232.860 181.735 ;
        RECT 231.705 181.515 232.115 181.525 ;
        RECT 231.925 181.175 232.380 181.345 ;
        RECT 232.690 180.785 232.860 181.565 ;
        RECT 231.125 180.465 231.910 180.695 ;
        RECT 231.580 180.325 231.910 180.465 ;
        RECT 232.210 180.615 232.860 180.785 ;
        RECT 230.715 179.985 230.925 180.315 ;
        RECT 231.095 180.155 231.425 180.195 ;
        RECT 232.210 180.155 232.380 180.615 ;
        RECT 231.095 179.985 232.380 180.155 ;
        RECT 232.550 179.815 232.880 180.195 ;
        RECT 233.050 179.985 233.310 182.195 ;
        RECT 233.480 181.690 233.740 182.195 ;
        RECT 233.920 181.985 234.250 182.365 ;
        RECT 234.430 181.815 234.600 182.195 ;
        RECT 233.480 180.890 233.650 181.690 ;
        RECT 233.935 181.645 234.600 181.815 ;
        RECT 233.935 181.390 234.105 181.645 ;
        RECT 234.860 181.615 236.070 182.365 ;
        RECT 233.820 181.060 234.105 181.390 ;
        RECT 234.340 181.095 234.670 181.465 ;
        RECT 233.935 180.915 234.105 181.060 ;
        RECT 233.480 179.985 233.750 180.890 ;
        RECT 233.935 180.745 234.600 180.915 ;
        RECT 233.920 179.815 234.250 180.575 ;
        RECT 234.430 179.985 234.600 180.745 ;
        RECT 234.860 180.905 235.380 181.445 ;
        RECT 235.550 181.075 236.070 181.615 ;
        RECT 234.860 179.815 236.070 180.905 ;
        RECT 162.095 179.645 236.155 179.815 ;
        RECT 162.180 178.555 163.390 179.645 ;
        RECT 162.180 177.845 162.700 178.385 ;
        RECT 162.870 178.015 163.390 178.555 ;
        RECT 163.650 178.715 163.820 179.475 ;
        RECT 164.035 178.885 164.365 179.645 ;
        RECT 163.650 178.545 164.365 178.715 ;
        RECT 164.535 178.570 164.790 179.475 ;
        RECT 163.560 177.995 163.915 178.365 ;
        RECT 164.195 178.335 164.365 178.545 ;
        RECT 164.195 178.005 164.450 178.335 ;
        RECT 162.180 177.095 163.390 177.845 ;
        RECT 164.195 177.815 164.365 178.005 ;
        RECT 164.620 177.840 164.790 178.570 ;
        RECT 164.965 178.495 165.225 179.645 ;
        RECT 165.950 178.715 166.120 179.475 ;
        RECT 166.300 178.885 166.630 179.645 ;
        RECT 165.950 178.545 166.615 178.715 ;
        RECT 166.800 178.570 167.070 179.475 ;
        RECT 167.740 179.185 167.955 179.645 ;
        RECT 168.125 179.015 168.455 179.475 ;
        RECT 166.445 178.400 166.615 178.545 ;
        RECT 165.880 177.995 166.210 178.365 ;
        RECT 166.445 178.070 166.730 178.400 ;
        RECT 163.650 177.645 164.365 177.815 ;
        RECT 163.650 177.265 163.820 177.645 ;
        RECT 164.035 177.095 164.365 177.475 ;
        RECT 164.535 177.265 164.790 177.840 ;
        RECT 164.965 177.095 165.225 177.935 ;
        RECT 166.445 177.815 166.615 178.070 ;
        RECT 165.950 177.645 166.615 177.815 ;
        RECT 166.900 177.770 167.070 178.570 ;
        RECT 165.950 177.265 166.120 177.645 ;
        RECT 166.300 177.095 166.630 177.475 ;
        RECT 166.810 177.265 167.070 177.770 ;
        RECT 167.285 178.845 168.455 179.015 ;
        RECT 168.625 178.845 168.875 179.645 ;
        RECT 167.285 177.555 167.655 178.845 ;
        RECT 169.085 178.675 169.365 178.835 ;
        RECT 168.030 178.505 169.365 178.675 ;
        RECT 169.630 178.715 169.800 179.475 ;
        RECT 169.980 178.885 170.310 179.645 ;
        RECT 169.630 178.545 170.295 178.715 ;
        RECT 170.480 178.570 170.750 179.475 ;
        RECT 168.030 178.335 168.200 178.505 ;
        RECT 170.125 178.400 170.295 178.545 ;
        RECT 167.825 178.085 168.200 178.335 ;
        RECT 168.370 178.085 168.845 178.325 ;
        RECT 169.015 178.085 169.365 178.325 ;
        RECT 168.030 177.915 168.200 178.085 ;
        RECT 169.560 177.995 169.890 178.365 ;
        RECT 170.125 178.070 170.410 178.400 ;
        RECT 168.030 177.745 169.365 177.915 ;
        RECT 170.125 177.815 170.295 178.070 ;
        RECT 167.285 177.265 168.035 177.555 ;
        RECT 168.545 177.095 168.875 177.555 ;
        RECT 169.095 177.535 169.365 177.745 ;
        RECT 169.630 177.645 170.295 177.815 ;
        RECT 170.580 177.770 170.750 178.570 ;
        RECT 171.010 178.715 171.180 179.475 ;
        RECT 171.360 178.885 171.690 179.645 ;
        RECT 171.010 178.545 171.675 178.715 ;
        RECT 171.860 178.570 172.130 179.475 ;
        RECT 171.505 178.400 171.675 178.545 ;
        RECT 170.940 177.995 171.270 178.365 ;
        RECT 171.505 178.070 171.790 178.400 ;
        RECT 171.505 177.815 171.675 178.070 ;
        RECT 169.630 177.265 169.800 177.645 ;
        RECT 169.980 177.095 170.310 177.475 ;
        RECT 170.490 177.265 170.750 177.770 ;
        RECT 171.010 177.645 171.675 177.815 ;
        RECT 171.960 177.770 172.130 178.570 ;
        RECT 172.390 178.715 172.560 179.475 ;
        RECT 172.740 178.885 173.070 179.645 ;
        RECT 172.390 178.545 173.055 178.715 ;
        RECT 173.240 178.570 173.510 179.475 ;
        RECT 172.885 178.400 173.055 178.545 ;
        RECT 172.320 177.995 172.650 178.365 ;
        RECT 172.885 178.070 173.170 178.400 ;
        RECT 172.885 177.815 173.055 178.070 ;
        RECT 171.010 177.265 171.180 177.645 ;
        RECT 171.360 177.095 171.690 177.475 ;
        RECT 171.870 177.265 172.130 177.770 ;
        RECT 172.390 177.645 173.055 177.815 ;
        RECT 173.340 177.770 173.510 178.570 ;
        RECT 173.770 178.715 173.940 179.475 ;
        RECT 174.120 178.885 174.450 179.645 ;
        RECT 173.770 178.545 174.435 178.715 ;
        RECT 174.620 178.570 174.890 179.475 ;
        RECT 174.265 178.400 174.435 178.545 ;
        RECT 173.700 177.995 174.030 178.365 ;
        RECT 174.265 178.070 174.550 178.400 ;
        RECT 174.265 177.815 174.435 178.070 ;
        RECT 172.390 177.265 172.560 177.645 ;
        RECT 172.740 177.095 173.070 177.475 ;
        RECT 173.250 177.265 173.510 177.770 ;
        RECT 173.770 177.645 174.435 177.815 ;
        RECT 174.720 177.770 174.890 178.570 ;
        RECT 175.060 178.480 175.350 179.645 ;
        RECT 176.015 178.845 176.265 179.645 ;
        RECT 176.435 179.015 176.765 179.475 ;
        RECT 176.935 179.185 177.150 179.645 ;
        RECT 176.435 178.845 177.605 179.015 ;
        RECT 175.525 178.675 175.805 178.835 ;
        RECT 175.525 178.505 176.860 178.675 ;
        RECT 176.690 178.335 176.860 178.505 ;
        RECT 175.525 178.085 175.875 178.325 ;
        RECT 176.045 178.085 176.520 178.325 ;
        RECT 176.690 178.085 177.065 178.335 ;
        RECT 176.690 177.915 176.860 178.085 ;
        RECT 173.770 177.265 173.940 177.645 ;
        RECT 174.120 177.095 174.450 177.475 ;
        RECT 174.630 177.265 174.890 177.770 ;
        RECT 175.060 177.095 175.350 177.820 ;
        RECT 175.525 177.745 176.860 177.915 ;
        RECT 175.525 177.535 175.795 177.745 ;
        RECT 177.235 177.555 177.605 178.845 ;
        RECT 178.370 178.715 178.540 179.475 ;
        RECT 178.720 178.885 179.050 179.645 ;
        RECT 178.370 178.545 179.035 178.715 ;
        RECT 179.220 178.570 179.490 179.475 ;
        RECT 178.865 178.400 179.035 178.545 ;
        RECT 178.300 177.995 178.630 178.365 ;
        RECT 178.865 178.070 179.150 178.400 ;
        RECT 178.865 177.815 179.035 178.070 ;
        RECT 176.015 177.095 176.345 177.555 ;
        RECT 176.855 177.265 177.605 177.555 ;
        RECT 178.370 177.645 179.035 177.815 ;
        RECT 179.320 177.770 179.490 178.570 ;
        RECT 179.750 178.715 179.920 179.475 ;
        RECT 180.100 178.885 180.430 179.645 ;
        RECT 179.750 178.545 180.415 178.715 ;
        RECT 180.600 178.570 180.870 179.475 ;
        RECT 180.245 178.400 180.415 178.545 ;
        RECT 179.680 177.995 180.010 178.365 ;
        RECT 180.245 178.070 180.530 178.400 ;
        RECT 180.245 177.815 180.415 178.070 ;
        RECT 178.370 177.265 178.540 177.645 ;
        RECT 178.720 177.095 179.050 177.475 ;
        RECT 179.230 177.265 179.490 177.770 ;
        RECT 179.750 177.645 180.415 177.815 ;
        RECT 180.700 177.770 180.870 178.570 ;
        RECT 181.130 178.715 181.300 179.475 ;
        RECT 181.480 178.885 181.810 179.645 ;
        RECT 181.130 178.545 181.795 178.715 ;
        RECT 181.980 178.570 182.250 179.475 ;
        RECT 181.625 178.400 181.795 178.545 ;
        RECT 181.060 177.995 181.390 178.365 ;
        RECT 181.625 178.070 181.910 178.400 ;
        RECT 181.625 177.815 181.795 178.070 ;
        RECT 179.750 177.265 179.920 177.645 ;
        RECT 180.100 177.095 180.430 177.475 ;
        RECT 180.610 177.265 180.870 177.770 ;
        RECT 181.130 177.645 181.795 177.815 ;
        RECT 182.080 177.770 182.250 178.570 ;
        RECT 181.130 177.265 181.300 177.645 ;
        RECT 181.480 177.095 181.810 177.475 ;
        RECT 181.990 177.265 182.250 177.770 ;
        RECT 182.425 178.505 182.760 179.475 ;
        RECT 182.930 178.505 183.100 179.645 ;
        RECT 183.270 179.305 185.300 179.475 ;
        RECT 182.425 177.835 182.595 178.505 ;
        RECT 183.270 178.335 183.440 179.305 ;
        RECT 182.765 178.005 183.020 178.335 ;
        RECT 183.245 178.005 183.440 178.335 ;
        RECT 183.610 178.965 184.735 179.135 ;
        RECT 182.850 177.835 183.020 178.005 ;
        RECT 183.610 177.835 183.780 178.965 ;
        RECT 182.425 177.265 182.680 177.835 ;
        RECT 182.850 177.665 183.780 177.835 ;
        RECT 183.950 178.625 184.960 178.795 ;
        RECT 183.950 177.825 184.120 178.625 ;
        RECT 183.605 177.630 183.780 177.665 ;
        RECT 182.850 177.095 183.180 177.495 ;
        RECT 183.605 177.265 184.135 177.630 ;
        RECT 184.325 177.605 184.600 178.425 ;
        RECT 184.320 177.435 184.600 177.605 ;
        RECT 184.325 177.265 184.600 177.435 ;
        RECT 184.770 177.265 184.960 178.625 ;
        RECT 185.130 178.640 185.300 179.305 ;
        RECT 185.470 178.885 185.640 179.645 ;
        RECT 185.875 178.885 186.390 179.295 ;
        RECT 185.130 178.450 185.880 178.640 ;
        RECT 186.050 178.075 186.390 178.885 ;
        RECT 186.650 178.715 186.820 179.475 ;
        RECT 187.000 178.885 187.330 179.645 ;
        RECT 186.650 178.545 187.315 178.715 ;
        RECT 187.500 178.570 187.770 179.475 ;
        RECT 187.145 178.400 187.315 178.545 ;
        RECT 185.160 177.905 186.390 178.075 ;
        RECT 186.580 177.995 186.910 178.365 ;
        RECT 187.145 178.070 187.430 178.400 ;
        RECT 185.140 177.095 185.650 177.630 ;
        RECT 185.870 177.300 186.115 177.905 ;
        RECT 187.145 177.815 187.315 178.070 ;
        RECT 186.650 177.645 187.315 177.815 ;
        RECT 187.600 177.770 187.770 178.570 ;
        RECT 187.940 178.480 188.230 179.645 ;
        RECT 188.895 178.845 189.145 179.645 ;
        RECT 189.315 179.015 189.645 179.475 ;
        RECT 189.815 179.185 190.030 179.645 ;
        RECT 189.315 178.845 190.485 179.015 ;
        RECT 191.195 178.845 191.445 179.645 ;
        RECT 191.615 179.015 191.945 179.475 ;
        RECT 192.115 179.185 192.330 179.645 ;
        RECT 191.615 178.845 192.785 179.015 ;
        RECT 188.405 178.675 188.685 178.835 ;
        RECT 188.405 178.505 189.740 178.675 ;
        RECT 189.570 178.335 189.740 178.505 ;
        RECT 188.405 178.085 188.755 178.325 ;
        RECT 188.925 178.085 189.400 178.325 ;
        RECT 189.570 178.085 189.945 178.335 ;
        RECT 189.570 177.915 189.740 178.085 ;
        RECT 186.650 177.265 186.820 177.645 ;
        RECT 187.000 177.095 187.330 177.475 ;
        RECT 187.510 177.265 187.770 177.770 ;
        RECT 187.940 177.095 188.230 177.820 ;
        RECT 188.405 177.745 189.740 177.915 ;
        RECT 188.405 177.535 188.675 177.745 ;
        RECT 190.115 177.555 190.485 178.845 ;
        RECT 190.705 178.675 190.985 178.835 ;
        RECT 190.705 178.505 192.040 178.675 ;
        RECT 191.870 178.335 192.040 178.505 ;
        RECT 190.705 178.085 191.055 178.325 ;
        RECT 191.225 178.085 191.700 178.325 ;
        RECT 191.870 178.085 192.245 178.335 ;
        RECT 191.870 177.915 192.040 178.085 ;
        RECT 188.895 177.095 189.225 177.555 ;
        RECT 189.735 177.265 190.485 177.555 ;
        RECT 190.705 177.745 192.040 177.915 ;
        RECT 190.705 177.535 190.975 177.745 ;
        RECT 192.415 177.555 192.785 178.845 ;
        RECT 191.195 177.095 191.525 177.555 ;
        RECT 192.035 177.265 192.785 177.555 ;
        RECT 193.005 178.505 193.340 179.475 ;
        RECT 193.510 178.505 193.680 179.645 ;
        RECT 193.850 179.305 195.880 179.475 ;
        RECT 193.005 177.835 193.175 178.505 ;
        RECT 193.850 178.335 194.020 179.305 ;
        RECT 193.345 178.005 193.600 178.335 ;
        RECT 193.825 178.005 194.020 178.335 ;
        RECT 194.190 178.965 195.315 179.135 ;
        RECT 193.430 177.835 193.600 178.005 ;
        RECT 194.190 177.835 194.360 178.965 ;
        RECT 193.005 177.265 193.260 177.835 ;
        RECT 193.430 177.665 194.360 177.835 ;
        RECT 194.530 178.625 195.540 178.795 ;
        RECT 194.530 177.825 194.700 178.625 ;
        RECT 194.905 178.285 195.180 178.425 ;
        RECT 194.900 178.115 195.180 178.285 ;
        RECT 194.185 177.630 194.360 177.665 ;
        RECT 193.430 177.095 193.760 177.495 ;
        RECT 194.185 177.265 194.715 177.630 ;
        RECT 194.905 177.265 195.180 178.115 ;
        RECT 195.350 177.265 195.540 178.625 ;
        RECT 195.710 178.640 195.880 179.305 ;
        RECT 196.050 178.885 196.220 179.645 ;
        RECT 196.455 178.885 196.970 179.295 ;
        RECT 195.710 178.450 196.460 178.640 ;
        RECT 196.630 178.075 196.970 178.885 ;
        RECT 198.150 178.715 198.320 179.475 ;
        RECT 198.500 178.885 198.830 179.645 ;
        RECT 198.150 178.545 198.815 178.715 ;
        RECT 199.000 178.570 199.270 179.475 ;
        RECT 198.645 178.400 198.815 178.545 ;
        RECT 195.740 177.905 196.970 178.075 ;
        RECT 198.080 177.995 198.410 178.365 ;
        RECT 198.645 178.070 198.930 178.400 ;
        RECT 195.720 177.095 196.230 177.630 ;
        RECT 196.450 177.300 196.695 177.905 ;
        RECT 198.645 177.815 198.815 178.070 ;
        RECT 198.150 177.645 198.815 177.815 ;
        RECT 199.100 177.770 199.270 178.570 ;
        RECT 199.530 178.715 199.700 179.475 ;
        RECT 199.880 178.885 200.210 179.645 ;
        RECT 199.530 178.545 200.195 178.715 ;
        RECT 200.380 178.570 200.650 179.475 ;
        RECT 200.025 178.400 200.195 178.545 ;
        RECT 199.460 177.995 199.790 178.365 ;
        RECT 200.025 178.070 200.310 178.400 ;
        RECT 200.025 177.815 200.195 178.070 ;
        RECT 198.150 177.265 198.320 177.645 ;
        RECT 198.500 177.095 198.830 177.475 ;
        RECT 199.010 177.265 199.270 177.770 ;
        RECT 199.530 177.645 200.195 177.815 ;
        RECT 200.480 177.770 200.650 178.570 ;
        RECT 200.820 178.480 201.110 179.645 ;
        RECT 201.830 178.715 202.000 179.475 ;
        RECT 202.180 178.885 202.510 179.645 ;
        RECT 201.830 178.545 202.495 178.715 ;
        RECT 202.680 178.570 202.950 179.475 ;
        RECT 202.325 178.400 202.495 178.545 ;
        RECT 201.760 177.995 202.090 178.365 ;
        RECT 202.325 178.070 202.610 178.400 ;
        RECT 199.530 177.265 199.700 177.645 ;
        RECT 199.880 177.095 200.210 177.475 ;
        RECT 200.390 177.265 200.650 177.770 ;
        RECT 200.820 177.095 201.110 177.820 ;
        RECT 202.325 177.815 202.495 178.070 ;
        RECT 201.830 177.645 202.495 177.815 ;
        RECT 202.780 177.770 202.950 178.570 ;
        RECT 201.830 177.265 202.000 177.645 ;
        RECT 202.180 177.095 202.510 177.475 ;
        RECT 202.690 177.265 202.950 177.770 ;
        RECT 204.040 177.265 204.300 179.475 ;
        RECT 204.470 179.265 204.800 179.645 ;
        RECT 204.970 179.305 206.255 179.475 ;
        RECT 204.970 178.845 205.140 179.305 ;
        RECT 205.925 179.265 206.255 179.305 ;
        RECT 206.425 179.145 206.635 179.475 ;
        RECT 204.490 178.675 205.140 178.845 ;
        RECT 205.440 178.995 205.770 179.135 ;
        RECT 205.440 178.765 206.225 178.995 ;
        RECT 204.490 177.895 204.660 178.675 ;
        RECT 204.970 178.115 205.425 178.285 ;
        RECT 205.235 177.935 205.645 177.945 ;
        RECT 204.490 177.725 205.060 177.895 ;
        RECT 204.550 177.095 204.720 177.555 ;
        RECT 204.890 177.435 205.060 177.725 ;
        RECT 205.230 177.775 205.645 177.935 ;
        RECT 205.230 177.605 205.405 177.775 ;
        RECT 206.055 177.595 206.225 178.765 ;
        RECT 206.465 177.945 206.635 179.145 ;
        RECT 206.930 179.145 207.115 179.475 ;
        RECT 207.285 179.265 207.635 179.645 ;
        RECT 206.930 178.285 207.100 179.145 ;
        RECT 207.885 179.095 208.055 179.475 ;
        RECT 208.225 179.265 208.555 179.645 ;
        RECT 208.780 179.305 209.790 179.475 ;
        RECT 208.780 179.095 208.950 179.305 ;
        RECT 207.885 178.925 208.950 179.095 ;
        RECT 206.810 178.115 207.100 178.285 ;
        RECT 206.395 177.775 206.635 177.945 ;
        RECT 206.930 177.665 207.100 178.115 ;
        RECT 207.270 178.005 207.560 178.685 ;
        RECT 208.035 178.065 208.365 178.685 ;
        RECT 208.570 178.285 208.815 178.685 ;
        RECT 209.120 178.625 209.450 179.135 ;
        RECT 209.620 178.795 209.790 179.305 ;
        RECT 210.050 179.265 210.380 179.645 ;
        RECT 209.120 178.455 209.880 178.625 ;
        RECT 208.570 178.115 208.870 178.285 ;
        RECT 209.155 178.275 209.325 178.285 ;
        RECT 209.155 178.115 209.540 178.275 ;
        RECT 208.570 178.065 208.815 178.115 ;
        RECT 209.210 178.105 209.540 178.115 ;
        RECT 209.225 177.895 209.395 177.935 ;
        RECT 209.710 177.930 209.880 178.455 ;
        RECT 210.050 178.005 210.350 179.005 ;
        RECT 210.550 178.635 210.900 179.475 ;
        RECT 211.070 179.305 212.600 179.475 ;
        RECT 211.070 178.805 211.240 179.305 ;
        RECT 212.430 179.145 212.600 179.305 ;
        RECT 212.770 179.265 213.100 179.645 ;
        RECT 211.410 178.965 211.740 179.135 ;
        RECT 211.570 178.635 211.740 178.965 ;
        RECT 211.910 178.975 212.080 179.135 ;
        RECT 213.270 178.975 213.440 179.475 ;
        RECT 211.910 178.805 213.440 178.975 ;
        RECT 210.550 178.405 211.355 178.635 ;
        RECT 211.570 178.465 212.205 178.635 ;
        RECT 210.995 178.295 211.355 178.405 ;
        RECT 210.995 178.115 211.535 178.295 ;
        RECT 207.875 177.725 209.395 177.895 ;
        RECT 205.715 177.435 205.885 177.595 ;
        RECT 204.890 177.265 205.885 177.435 ;
        RECT 206.055 177.425 206.585 177.595 ;
        RECT 206.415 177.265 206.585 177.425 ;
        RECT 206.930 177.335 207.105 177.665 ;
        RECT 207.275 177.095 207.605 177.475 ;
        RECT 207.875 177.305 208.120 177.725 ;
        RECT 209.225 177.605 209.395 177.725 ;
        RECT 209.565 177.855 209.880 177.930 ;
        RECT 209.565 177.605 209.895 177.855 ;
        RECT 208.295 177.095 208.465 177.555 ;
        RECT 208.635 177.435 208.990 177.475 ;
        RECT 210.065 177.435 210.235 177.805 ;
        RECT 208.635 177.265 210.235 177.435 ;
        RECT 210.525 177.095 210.815 177.815 ;
        RECT 210.995 177.440 211.355 178.115 ;
        RECT 212.035 177.945 212.205 178.465 ;
        RECT 212.375 178.005 212.810 178.625 ;
        RECT 213.120 178.455 213.470 178.625 ;
        RECT 213.700 178.480 213.990 179.645 ;
        RECT 214.250 178.715 214.420 179.475 ;
        RECT 214.600 178.885 214.930 179.645 ;
        RECT 214.250 178.545 214.915 178.715 ;
        RECT 215.100 178.570 215.370 179.475 ;
        RECT 213.120 178.005 213.465 178.455 ;
        RECT 214.745 178.400 214.915 178.545 ;
        RECT 214.180 177.995 214.510 178.365 ;
        RECT 214.745 178.070 215.030 178.400 ;
        RECT 211.915 177.775 212.205 177.945 ;
        RECT 211.525 177.435 211.695 177.770 ;
        RECT 211.865 177.605 212.205 177.775 ;
        RECT 212.430 177.645 213.440 177.815 ;
        RECT 212.430 177.435 212.600 177.645 ;
        RECT 211.525 177.265 212.600 177.435 ;
        RECT 212.770 177.095 213.100 177.475 ;
        RECT 213.270 177.270 213.440 177.645 ;
        RECT 213.700 177.095 213.990 177.820 ;
        RECT 214.745 177.815 214.915 178.070 ;
        RECT 214.250 177.645 214.915 177.815 ;
        RECT 215.200 177.770 215.370 178.570 ;
        RECT 215.630 178.715 215.800 179.475 ;
        RECT 215.980 178.885 216.310 179.645 ;
        RECT 215.630 178.545 216.295 178.715 ;
        RECT 216.480 178.570 216.750 179.475 ;
        RECT 217.010 178.975 217.180 179.475 ;
        RECT 217.350 179.265 217.680 179.645 ;
        RECT 217.850 179.305 219.380 179.475 ;
        RECT 217.850 179.145 218.020 179.305 ;
        RECT 218.370 178.975 218.540 179.135 ;
        RECT 217.010 178.805 218.540 178.975 ;
        RECT 218.710 178.965 219.040 179.135 ;
        RECT 218.710 178.635 218.880 178.965 ;
        RECT 219.210 178.805 219.380 179.305 ;
        RECT 219.550 178.635 219.900 179.475 ;
        RECT 220.070 179.265 220.400 179.645 ;
        RECT 220.660 179.305 221.670 179.475 ;
        RECT 216.125 178.400 216.295 178.545 ;
        RECT 215.560 177.995 215.890 178.365 ;
        RECT 216.125 178.070 216.410 178.400 ;
        RECT 216.125 177.815 216.295 178.070 ;
        RECT 214.250 177.265 214.420 177.645 ;
        RECT 214.600 177.095 214.930 177.475 ;
        RECT 215.110 177.265 215.370 177.770 ;
        RECT 215.630 177.645 216.295 177.815 ;
        RECT 216.580 177.770 216.750 178.570 ;
        RECT 216.980 178.455 217.330 178.625 ;
        RECT 216.985 178.005 217.330 178.455 ;
        RECT 217.640 178.005 218.075 178.625 ;
        RECT 218.245 178.465 218.880 178.635 ;
        RECT 218.245 177.945 218.415 178.465 ;
        RECT 219.095 178.405 219.900 178.635 ;
        RECT 219.095 178.295 219.455 178.405 ;
        RECT 218.915 178.115 219.455 178.295 ;
        RECT 215.630 177.265 215.800 177.645 ;
        RECT 215.980 177.095 216.310 177.475 ;
        RECT 216.490 177.265 216.750 177.770 ;
        RECT 217.010 177.645 218.020 177.815 ;
        RECT 217.010 177.270 217.180 177.645 ;
        RECT 217.350 177.095 217.680 177.475 ;
        RECT 217.850 177.435 218.020 177.645 ;
        RECT 218.245 177.775 218.535 177.945 ;
        RECT 218.245 177.605 218.585 177.775 ;
        RECT 218.755 177.435 218.925 177.770 ;
        RECT 219.095 177.440 219.455 178.115 ;
        RECT 220.100 178.005 220.400 179.005 ;
        RECT 220.660 178.795 220.830 179.305 ;
        RECT 221.000 178.625 221.330 179.135 ;
        RECT 221.500 179.095 221.670 179.305 ;
        RECT 221.895 179.265 222.225 179.645 ;
        RECT 222.395 179.095 222.565 179.475 ;
        RECT 222.815 179.265 223.165 179.645 ;
        RECT 223.335 179.145 223.520 179.475 ;
        RECT 221.500 178.925 222.565 179.095 ;
        RECT 221.635 178.625 221.880 178.685 ;
        RECT 220.570 178.455 221.330 178.625 ;
        RECT 221.580 178.455 221.880 178.625 ;
        RECT 220.570 177.930 220.740 178.455 ;
        RECT 221.125 178.275 221.295 178.285 ;
        RECT 220.910 178.115 221.295 178.275 ;
        RECT 220.910 178.105 221.240 178.115 ;
        RECT 221.635 178.065 221.880 178.455 ;
        RECT 222.085 178.625 222.415 178.685 ;
        RECT 222.085 178.455 222.440 178.625 ;
        RECT 222.085 178.065 222.415 178.455 ;
        RECT 222.890 178.005 223.180 178.685 ;
        RECT 223.350 178.285 223.520 179.145 ;
        RECT 223.815 179.145 224.025 179.475 ;
        RECT 224.195 179.305 225.480 179.475 ;
        RECT 224.195 179.265 224.525 179.305 ;
        RECT 223.350 178.115 223.640 178.285 ;
        RECT 220.570 177.855 220.885 177.930 ;
        RECT 217.850 177.265 218.925 177.435 ;
        RECT 219.635 177.095 219.925 177.815 ;
        RECT 220.215 177.435 220.385 177.805 ;
        RECT 220.555 177.605 220.885 177.855 ;
        RECT 221.055 177.895 221.225 177.935 ;
        RECT 221.055 177.725 222.575 177.895 ;
        RECT 221.055 177.605 221.225 177.725 ;
        RECT 221.460 177.435 221.815 177.475 ;
        RECT 220.215 177.265 221.815 177.435 ;
        RECT 221.985 177.095 222.155 177.555 ;
        RECT 222.330 177.305 222.575 177.725 ;
        RECT 223.350 177.665 223.520 178.115 ;
        RECT 223.815 177.945 223.985 179.145 ;
        RECT 224.680 178.995 225.010 179.135 ;
        RECT 224.225 178.765 225.010 178.995 ;
        RECT 225.310 178.845 225.480 179.305 ;
        RECT 225.650 179.265 225.980 179.645 ;
        RECT 223.815 177.775 224.055 177.945 ;
        RECT 222.845 177.095 223.175 177.475 ;
        RECT 223.345 177.335 223.520 177.665 ;
        RECT 224.225 177.595 224.395 178.765 ;
        RECT 225.310 178.675 225.960 178.845 ;
        RECT 225.025 178.115 225.480 178.285 ;
        RECT 224.805 177.935 225.215 177.945 ;
        RECT 224.805 177.775 225.220 177.935 ;
        RECT 225.790 177.895 225.960 178.675 ;
        RECT 225.045 177.605 225.220 177.775 ;
        RECT 225.390 177.725 225.960 177.895 ;
        RECT 223.865 177.425 224.395 177.595 ;
        RECT 224.565 177.435 224.735 177.595 ;
        RECT 225.390 177.435 225.560 177.725 ;
        RECT 223.865 177.265 224.035 177.425 ;
        RECT 224.565 177.265 225.560 177.435 ;
        RECT 225.730 177.095 225.900 177.555 ;
        RECT 226.150 177.265 226.410 179.475 ;
        RECT 226.580 178.480 226.870 179.645 ;
        RECT 227.040 178.570 227.310 179.475 ;
        RECT 227.480 178.885 227.810 179.645 ;
        RECT 227.990 178.715 228.160 179.475 ;
        RECT 226.580 177.095 226.870 177.820 ;
        RECT 227.040 177.770 227.210 178.570 ;
        RECT 227.495 178.545 228.160 178.715 ;
        RECT 228.420 178.570 228.690 179.475 ;
        RECT 228.860 178.885 229.190 179.645 ;
        RECT 229.370 178.715 229.540 179.475 ;
        RECT 227.495 178.400 227.665 178.545 ;
        RECT 227.380 178.070 227.665 178.400 ;
        RECT 227.495 177.815 227.665 178.070 ;
        RECT 227.900 177.995 228.230 178.365 ;
        RECT 227.040 177.265 227.300 177.770 ;
        RECT 227.495 177.645 228.160 177.815 ;
        RECT 227.480 177.095 227.810 177.475 ;
        RECT 227.990 177.265 228.160 177.645 ;
        RECT 228.420 177.770 228.590 178.570 ;
        RECT 228.875 178.545 229.540 178.715 ;
        RECT 229.800 178.570 230.070 179.475 ;
        RECT 230.240 178.885 230.570 179.645 ;
        RECT 230.750 178.715 230.920 179.475 ;
        RECT 228.875 178.400 229.045 178.545 ;
        RECT 228.760 178.070 229.045 178.400 ;
        RECT 228.875 177.815 229.045 178.070 ;
        RECT 229.280 177.995 229.610 178.365 ;
        RECT 228.420 177.265 228.680 177.770 ;
        RECT 228.875 177.645 229.540 177.815 ;
        RECT 228.860 177.095 229.190 177.475 ;
        RECT 229.370 177.265 229.540 177.645 ;
        RECT 229.800 177.770 229.970 178.570 ;
        RECT 230.255 178.545 230.920 178.715 ;
        RECT 231.180 178.570 231.450 179.475 ;
        RECT 231.620 178.885 231.950 179.645 ;
        RECT 232.130 178.715 232.300 179.475 ;
        RECT 230.255 178.400 230.425 178.545 ;
        RECT 230.140 178.070 230.425 178.400 ;
        RECT 230.255 177.815 230.425 178.070 ;
        RECT 230.660 177.995 230.990 178.365 ;
        RECT 229.800 177.265 230.060 177.770 ;
        RECT 230.255 177.645 230.920 177.815 ;
        RECT 230.240 177.095 230.570 177.475 ;
        RECT 230.750 177.265 230.920 177.645 ;
        RECT 231.180 177.770 231.350 178.570 ;
        RECT 231.635 178.545 232.300 178.715 ;
        RECT 232.560 178.570 232.830 179.475 ;
        RECT 233.000 178.885 233.330 179.645 ;
        RECT 233.510 178.715 233.680 179.475 ;
        RECT 231.635 178.400 231.805 178.545 ;
        RECT 231.520 178.070 231.805 178.400 ;
        RECT 231.635 177.815 231.805 178.070 ;
        RECT 232.040 177.995 232.370 178.365 ;
        RECT 231.180 177.265 231.440 177.770 ;
        RECT 231.635 177.645 232.300 177.815 ;
        RECT 231.620 177.095 231.950 177.475 ;
        RECT 232.130 177.265 232.300 177.645 ;
        RECT 232.560 177.770 232.730 178.570 ;
        RECT 233.015 178.545 233.680 178.715 ;
        RECT 234.860 178.555 236.070 179.645 ;
        RECT 233.015 178.400 233.185 178.545 ;
        RECT 232.900 178.070 233.185 178.400 ;
        RECT 233.015 177.815 233.185 178.070 ;
        RECT 233.420 177.995 233.750 178.365 ;
        RECT 234.860 178.015 235.380 178.555 ;
        RECT 235.550 177.845 236.070 178.385 ;
        RECT 232.560 177.265 232.820 177.770 ;
        RECT 233.015 177.645 233.680 177.815 ;
        RECT 233.000 177.095 233.330 177.475 ;
        RECT 233.510 177.265 233.680 177.645 ;
        RECT 234.860 177.095 236.070 177.845 ;
        RECT 162.095 176.925 236.155 177.095 ;
        RECT 162.095 106.340 311.135 106.510 ;
        RECT 162.180 105.590 163.390 106.340 ;
        RECT 162.180 105.050 162.700 105.590 ;
        RECT 163.565 105.500 163.825 106.340 ;
        RECT 164.000 105.595 164.255 106.170 ;
        RECT 164.425 105.960 164.755 106.340 ;
        RECT 164.970 105.790 165.140 106.170 ;
        RECT 164.425 105.620 165.140 105.790 ;
        RECT 162.870 104.880 163.390 105.420 ;
        RECT 162.180 103.790 163.390 104.880 ;
        RECT 163.565 103.790 163.825 104.940 ;
        RECT 164.000 104.865 164.170 105.595 ;
        RECT 164.425 105.430 164.595 105.620 ;
        RECT 165.405 105.500 165.665 106.340 ;
        RECT 165.840 105.595 166.095 106.170 ;
        RECT 166.265 105.960 166.595 106.340 ;
        RECT 166.810 105.790 166.980 106.170 ;
        RECT 166.265 105.620 166.980 105.790 ;
        RECT 164.340 105.100 164.595 105.430 ;
        RECT 164.425 104.890 164.595 105.100 ;
        RECT 164.875 105.070 165.230 105.440 ;
        RECT 164.000 103.960 164.255 104.865 ;
        RECT 164.425 104.720 165.140 104.890 ;
        RECT 164.425 103.790 164.755 104.550 ;
        RECT 164.970 103.960 165.140 104.720 ;
        RECT 165.405 103.790 165.665 104.940 ;
        RECT 165.840 104.865 166.010 105.595 ;
        RECT 166.265 105.430 166.435 105.620 ;
        RECT 167.245 105.500 167.505 106.340 ;
        RECT 167.680 105.595 167.935 106.170 ;
        RECT 168.105 105.960 168.435 106.340 ;
        RECT 168.650 105.790 168.820 106.170 ;
        RECT 168.105 105.620 168.820 105.790 ;
        RECT 166.180 105.100 166.435 105.430 ;
        RECT 166.265 104.890 166.435 105.100 ;
        RECT 166.715 105.070 167.070 105.440 ;
        RECT 165.840 103.960 166.095 104.865 ;
        RECT 166.265 104.720 166.980 104.890 ;
        RECT 166.265 103.790 166.595 104.550 ;
        RECT 166.810 103.960 166.980 104.720 ;
        RECT 167.245 103.790 167.505 104.940 ;
        RECT 167.680 104.865 167.850 105.595 ;
        RECT 168.105 105.430 168.275 105.620 ;
        RECT 169.085 105.500 169.345 106.340 ;
        RECT 169.520 105.595 169.775 106.170 ;
        RECT 169.945 105.960 170.275 106.340 ;
        RECT 170.490 105.790 170.660 106.170 ;
        RECT 169.945 105.620 170.660 105.790 ;
        RECT 168.020 105.100 168.275 105.430 ;
        RECT 168.105 104.890 168.275 105.100 ;
        RECT 168.555 105.070 168.910 105.440 ;
        RECT 167.680 103.960 167.935 104.865 ;
        RECT 168.105 104.720 168.820 104.890 ;
        RECT 168.105 103.790 168.435 104.550 ;
        RECT 168.650 103.960 168.820 104.720 ;
        RECT 169.085 103.790 169.345 104.940 ;
        RECT 169.520 104.865 169.690 105.595 ;
        RECT 169.945 105.430 170.115 105.620 ;
        RECT 170.925 105.600 171.180 106.170 ;
        RECT 171.350 105.940 171.680 106.340 ;
        RECT 172.105 105.805 172.635 106.170 ;
        RECT 172.105 105.770 172.280 105.805 ;
        RECT 171.350 105.600 172.280 105.770 ;
        RECT 169.860 105.100 170.115 105.430 ;
        RECT 169.945 104.890 170.115 105.100 ;
        RECT 170.395 105.070 170.750 105.440 ;
        RECT 170.925 104.930 171.095 105.600 ;
        RECT 171.350 105.430 171.520 105.600 ;
        RECT 171.265 105.100 171.520 105.430 ;
        RECT 171.745 105.100 171.940 105.430 ;
        RECT 169.520 103.960 169.775 104.865 ;
        RECT 169.945 104.720 170.660 104.890 ;
        RECT 169.945 103.790 170.275 104.550 ;
        RECT 170.490 103.960 170.660 104.720 ;
        RECT 170.925 103.960 171.260 104.930 ;
        RECT 171.430 103.790 171.600 104.930 ;
        RECT 171.770 104.130 171.940 105.100 ;
        RECT 172.110 104.470 172.280 105.600 ;
        RECT 172.450 104.810 172.620 105.610 ;
        RECT 172.825 105.320 173.100 106.170 ;
        RECT 172.820 105.150 173.100 105.320 ;
        RECT 172.825 105.010 173.100 105.150 ;
        RECT 173.270 104.810 173.460 106.170 ;
        RECT 173.640 105.805 174.150 106.340 ;
        RECT 174.370 105.530 174.615 106.135 ;
        RECT 175.060 105.615 175.350 106.340 ;
        RECT 175.525 105.600 175.780 106.170 ;
        RECT 175.950 105.940 176.280 106.340 ;
        RECT 176.705 105.805 177.235 106.170 ;
        RECT 176.705 105.770 176.880 105.805 ;
        RECT 175.950 105.600 176.880 105.770 ;
        RECT 173.660 105.360 174.890 105.530 ;
        RECT 172.450 104.640 173.460 104.810 ;
        RECT 173.630 104.795 174.380 104.985 ;
        RECT 172.110 104.300 173.235 104.470 ;
        RECT 173.630 104.130 173.800 104.795 ;
        RECT 174.550 104.550 174.890 105.360 ;
        RECT 171.770 103.960 173.800 104.130 ;
        RECT 173.970 103.790 174.140 104.550 ;
        RECT 174.375 104.140 174.890 104.550 ;
        RECT 175.060 103.790 175.350 104.955 ;
        RECT 175.525 104.930 175.695 105.600 ;
        RECT 175.950 105.430 176.120 105.600 ;
        RECT 175.865 105.100 176.120 105.430 ;
        RECT 176.345 105.100 176.540 105.430 ;
        RECT 175.525 103.960 175.860 104.930 ;
        RECT 176.030 103.790 176.200 104.930 ;
        RECT 176.370 104.130 176.540 105.100 ;
        RECT 176.710 104.470 176.880 105.600 ;
        RECT 177.050 104.810 177.220 105.610 ;
        RECT 177.425 105.320 177.700 106.170 ;
        RECT 177.420 105.150 177.700 105.320 ;
        RECT 177.425 105.010 177.700 105.150 ;
        RECT 177.870 104.810 178.060 106.170 ;
        RECT 178.240 105.805 178.750 106.340 ;
        RECT 178.970 105.530 179.215 106.135 ;
        RECT 180.670 105.790 180.840 106.170 ;
        RECT 181.055 105.960 181.385 106.340 ;
        RECT 180.670 105.620 181.385 105.790 ;
        RECT 178.260 105.360 179.490 105.530 ;
        RECT 177.050 104.640 178.060 104.810 ;
        RECT 178.230 104.795 178.980 104.985 ;
        RECT 176.710 104.300 177.835 104.470 ;
        RECT 178.230 104.130 178.400 104.795 ;
        RECT 179.150 104.550 179.490 105.360 ;
        RECT 180.580 105.070 180.935 105.440 ;
        RECT 181.215 105.430 181.385 105.620 ;
        RECT 181.555 105.595 181.810 106.170 ;
        RECT 181.215 105.100 181.470 105.430 ;
        RECT 181.215 104.890 181.385 105.100 ;
        RECT 176.370 103.960 178.400 104.130 ;
        RECT 178.570 103.790 178.740 104.550 ;
        RECT 178.975 104.140 179.490 104.550 ;
        RECT 180.670 104.720 181.385 104.890 ;
        RECT 181.640 104.865 181.810 105.595 ;
        RECT 181.985 105.500 182.245 106.340 ;
        RECT 182.510 105.790 182.680 106.170 ;
        RECT 182.895 105.960 183.225 106.340 ;
        RECT 182.510 105.620 183.225 105.790 ;
        RECT 182.420 105.070 182.775 105.440 ;
        RECT 183.055 105.430 183.225 105.620 ;
        RECT 183.395 105.595 183.650 106.170 ;
        RECT 183.055 105.100 183.310 105.430 ;
        RECT 180.670 103.960 180.840 104.720 ;
        RECT 181.055 103.790 181.385 104.550 ;
        RECT 181.555 103.960 181.810 104.865 ;
        RECT 181.985 103.790 182.245 104.940 ;
        RECT 183.055 104.890 183.225 105.100 ;
        RECT 182.510 104.720 183.225 104.890 ;
        RECT 183.480 104.865 183.650 105.595 ;
        RECT 183.825 105.500 184.085 106.340 ;
        RECT 184.350 105.790 184.520 106.170 ;
        RECT 184.735 105.960 185.065 106.340 ;
        RECT 184.350 105.620 185.065 105.790 ;
        RECT 184.260 105.070 184.615 105.440 ;
        RECT 184.895 105.430 185.065 105.620 ;
        RECT 185.235 105.595 185.490 106.170 ;
        RECT 184.895 105.100 185.150 105.430 ;
        RECT 182.510 103.960 182.680 104.720 ;
        RECT 182.895 103.790 183.225 104.550 ;
        RECT 183.395 103.960 183.650 104.865 ;
        RECT 183.825 103.790 184.085 104.940 ;
        RECT 184.895 104.890 185.065 105.100 ;
        RECT 184.350 104.720 185.065 104.890 ;
        RECT 185.320 104.865 185.490 105.595 ;
        RECT 185.665 105.500 185.925 106.340 ;
        RECT 186.190 105.790 186.360 106.170 ;
        RECT 186.575 105.960 186.905 106.340 ;
        RECT 186.190 105.620 186.905 105.790 ;
        RECT 186.100 105.070 186.455 105.440 ;
        RECT 186.735 105.430 186.905 105.620 ;
        RECT 187.075 105.595 187.330 106.170 ;
        RECT 186.735 105.100 186.990 105.430 ;
        RECT 184.350 103.960 184.520 104.720 ;
        RECT 184.735 103.790 185.065 104.550 ;
        RECT 185.235 103.960 185.490 104.865 ;
        RECT 185.665 103.790 185.925 104.940 ;
        RECT 186.735 104.890 186.905 105.100 ;
        RECT 186.190 104.720 186.905 104.890 ;
        RECT 187.160 104.865 187.330 105.595 ;
        RECT 187.505 105.500 187.765 106.340 ;
        RECT 187.940 105.615 188.230 106.340 ;
        RECT 188.865 105.600 189.120 106.170 ;
        RECT 189.290 105.940 189.620 106.340 ;
        RECT 190.045 105.805 190.575 106.170 ;
        RECT 190.045 105.770 190.220 105.805 ;
        RECT 189.290 105.600 190.220 105.770 ;
        RECT 186.190 103.960 186.360 104.720 ;
        RECT 186.575 103.790 186.905 104.550 ;
        RECT 187.075 103.960 187.330 104.865 ;
        RECT 187.505 103.790 187.765 104.940 ;
        RECT 187.940 103.790 188.230 104.955 ;
        RECT 188.865 104.930 189.035 105.600 ;
        RECT 189.290 105.430 189.460 105.600 ;
        RECT 189.205 105.100 189.460 105.430 ;
        RECT 189.685 105.100 189.880 105.430 ;
        RECT 188.865 103.960 189.200 104.930 ;
        RECT 189.370 103.790 189.540 104.930 ;
        RECT 189.710 104.130 189.880 105.100 ;
        RECT 190.050 104.470 190.220 105.600 ;
        RECT 190.390 104.810 190.560 105.610 ;
        RECT 190.765 105.320 191.040 106.170 ;
        RECT 190.760 105.150 191.040 105.320 ;
        RECT 190.765 105.010 191.040 105.150 ;
        RECT 191.210 104.810 191.400 106.170 ;
        RECT 191.580 105.805 192.090 106.340 ;
        RECT 192.310 105.530 192.555 106.135 ;
        RECT 193.550 105.790 193.720 106.170 ;
        RECT 193.935 105.960 194.265 106.340 ;
        RECT 193.550 105.620 194.265 105.790 ;
        RECT 191.600 105.360 192.830 105.530 ;
        RECT 190.390 104.640 191.400 104.810 ;
        RECT 191.570 104.795 192.320 104.985 ;
        RECT 190.050 104.300 191.175 104.470 ;
        RECT 191.570 104.130 191.740 104.795 ;
        RECT 192.490 104.550 192.830 105.360 ;
        RECT 193.460 105.070 193.815 105.440 ;
        RECT 194.095 105.430 194.265 105.620 ;
        RECT 194.435 105.595 194.690 106.170 ;
        RECT 194.095 105.100 194.350 105.430 ;
        RECT 194.095 104.890 194.265 105.100 ;
        RECT 189.710 103.960 191.740 104.130 ;
        RECT 191.910 103.790 192.080 104.550 ;
        RECT 192.315 104.140 192.830 104.550 ;
        RECT 193.550 104.720 194.265 104.890 ;
        RECT 194.520 104.865 194.690 105.595 ;
        RECT 194.865 105.500 195.125 106.340 ;
        RECT 195.390 105.790 195.560 106.170 ;
        RECT 195.775 105.960 196.105 106.340 ;
        RECT 195.390 105.620 196.105 105.790 ;
        RECT 195.300 105.070 195.655 105.440 ;
        RECT 195.935 105.430 196.105 105.620 ;
        RECT 196.275 105.595 196.530 106.170 ;
        RECT 195.935 105.100 196.190 105.430 ;
        RECT 193.550 103.960 193.720 104.720 ;
        RECT 193.935 103.790 194.265 104.550 ;
        RECT 194.435 103.960 194.690 104.865 ;
        RECT 194.865 103.790 195.125 104.940 ;
        RECT 195.935 104.890 196.105 105.100 ;
        RECT 195.390 104.720 196.105 104.890 ;
        RECT 196.360 104.865 196.530 105.595 ;
        RECT 196.705 105.500 196.965 106.340 ;
        RECT 197.230 105.790 197.400 106.170 ;
        RECT 197.615 105.960 197.945 106.340 ;
        RECT 197.230 105.620 197.945 105.790 ;
        RECT 197.140 105.070 197.495 105.440 ;
        RECT 197.775 105.430 197.945 105.620 ;
        RECT 198.115 105.595 198.370 106.170 ;
        RECT 197.775 105.100 198.030 105.430 ;
        RECT 195.390 103.960 195.560 104.720 ;
        RECT 195.775 103.790 196.105 104.550 ;
        RECT 196.275 103.960 196.530 104.865 ;
        RECT 196.705 103.790 196.965 104.940 ;
        RECT 197.775 104.890 197.945 105.100 ;
        RECT 197.230 104.720 197.945 104.890 ;
        RECT 198.200 104.865 198.370 105.595 ;
        RECT 198.545 105.500 198.805 106.340 ;
        RECT 199.070 105.790 199.240 106.170 ;
        RECT 199.455 105.960 199.785 106.340 ;
        RECT 199.070 105.620 199.785 105.790 ;
        RECT 198.980 105.070 199.335 105.440 ;
        RECT 199.615 105.430 199.785 105.620 ;
        RECT 199.955 105.595 200.210 106.170 ;
        RECT 199.615 105.100 199.870 105.430 ;
        RECT 197.230 103.960 197.400 104.720 ;
        RECT 197.615 103.790 197.945 104.550 ;
        RECT 198.115 103.960 198.370 104.865 ;
        RECT 198.545 103.790 198.805 104.940 ;
        RECT 199.615 104.890 199.785 105.100 ;
        RECT 199.070 104.720 199.785 104.890 ;
        RECT 200.040 104.865 200.210 105.595 ;
        RECT 200.385 105.500 200.645 106.340 ;
        RECT 200.820 105.615 201.110 106.340 ;
        RECT 201.280 105.590 202.490 106.340 ;
        RECT 202.750 105.790 202.920 106.170 ;
        RECT 203.135 105.960 203.465 106.340 ;
        RECT 202.750 105.620 203.465 105.790 ;
        RECT 201.280 105.050 201.800 105.590 ;
        RECT 199.070 103.960 199.240 104.720 ;
        RECT 199.455 103.790 199.785 104.550 ;
        RECT 199.955 103.960 200.210 104.865 ;
        RECT 200.385 103.790 200.645 104.940 ;
        RECT 200.820 103.790 201.110 104.955 ;
        RECT 201.970 104.880 202.490 105.420 ;
        RECT 202.660 105.070 203.015 105.440 ;
        RECT 203.295 105.430 203.465 105.620 ;
        RECT 203.635 105.595 203.890 106.170 ;
        RECT 203.295 105.100 203.550 105.430 ;
        RECT 203.295 104.890 203.465 105.100 ;
        RECT 201.280 103.790 202.490 104.880 ;
        RECT 202.750 104.720 203.465 104.890 ;
        RECT 203.720 104.865 203.890 105.595 ;
        RECT 204.065 105.500 204.325 106.340 ;
        RECT 204.505 105.500 204.765 106.340 ;
        RECT 204.940 105.595 205.195 106.170 ;
        RECT 205.365 105.960 205.695 106.340 ;
        RECT 205.910 105.790 206.080 106.170 ;
        RECT 205.365 105.620 206.080 105.790 ;
        RECT 202.750 103.960 202.920 104.720 ;
        RECT 203.135 103.790 203.465 104.550 ;
        RECT 203.635 103.960 203.890 104.865 ;
        RECT 204.065 103.790 204.325 104.940 ;
        RECT 204.505 103.790 204.765 104.940 ;
        RECT 204.940 104.865 205.110 105.595 ;
        RECT 205.365 105.430 205.535 105.620 ;
        RECT 206.345 105.600 206.600 106.170 ;
        RECT 206.770 105.940 207.100 106.340 ;
        RECT 207.525 105.805 208.055 106.170 ;
        RECT 207.525 105.770 207.700 105.805 ;
        RECT 206.770 105.600 207.700 105.770 ;
        RECT 205.280 105.100 205.535 105.430 ;
        RECT 205.365 104.890 205.535 105.100 ;
        RECT 205.815 105.070 206.170 105.440 ;
        RECT 206.345 104.930 206.515 105.600 ;
        RECT 206.770 105.430 206.940 105.600 ;
        RECT 206.685 105.100 206.940 105.430 ;
        RECT 207.165 105.100 207.360 105.430 ;
        RECT 204.940 103.960 205.195 104.865 ;
        RECT 205.365 104.720 206.080 104.890 ;
        RECT 205.365 103.790 205.695 104.550 ;
        RECT 205.910 103.960 206.080 104.720 ;
        RECT 206.345 103.960 206.680 104.930 ;
        RECT 206.850 103.790 207.020 104.930 ;
        RECT 207.190 104.130 207.360 105.100 ;
        RECT 207.530 104.470 207.700 105.600 ;
        RECT 207.870 104.810 208.040 105.610 ;
        RECT 208.245 105.320 208.520 106.170 ;
        RECT 208.240 105.150 208.520 105.320 ;
        RECT 208.245 105.010 208.520 105.150 ;
        RECT 208.690 104.810 208.880 106.170 ;
        RECT 209.060 105.805 209.570 106.340 ;
        RECT 209.790 105.530 210.035 106.135 ;
        RECT 210.480 105.590 211.690 106.340 ;
        RECT 209.080 105.360 210.310 105.530 ;
        RECT 207.870 104.640 208.880 104.810 ;
        RECT 209.050 104.795 209.800 104.985 ;
        RECT 207.530 104.300 208.655 104.470 ;
        RECT 209.050 104.130 209.220 104.795 ;
        RECT 209.970 104.550 210.310 105.360 ;
        RECT 210.480 105.050 211.000 105.590 ;
        RECT 211.865 105.500 212.125 106.340 ;
        RECT 212.300 105.595 212.555 106.170 ;
        RECT 212.725 105.960 213.055 106.340 ;
        RECT 213.270 105.790 213.440 106.170 ;
        RECT 212.725 105.620 213.440 105.790 ;
        RECT 211.170 104.880 211.690 105.420 ;
        RECT 207.190 103.960 209.220 104.130 ;
        RECT 209.390 103.790 209.560 104.550 ;
        RECT 209.795 104.140 210.310 104.550 ;
        RECT 210.480 103.790 211.690 104.880 ;
        RECT 211.865 103.790 212.125 104.940 ;
        RECT 212.300 104.865 212.470 105.595 ;
        RECT 212.725 105.430 212.895 105.620 ;
        RECT 213.700 105.615 213.990 106.340 ;
        RECT 214.160 105.590 215.370 106.340 ;
        RECT 212.640 105.100 212.895 105.430 ;
        RECT 212.725 104.890 212.895 105.100 ;
        RECT 213.175 105.070 213.530 105.440 ;
        RECT 214.160 105.050 214.680 105.590 ;
        RECT 215.545 105.500 215.805 106.340 ;
        RECT 215.980 105.595 216.235 106.170 ;
        RECT 216.405 105.960 216.735 106.340 ;
        RECT 216.950 105.790 217.120 106.170 ;
        RECT 216.405 105.620 217.120 105.790 ;
        RECT 217.470 105.790 217.640 106.170 ;
        RECT 217.855 105.960 218.185 106.340 ;
        RECT 217.470 105.620 218.185 105.790 ;
        RECT 212.300 103.960 212.555 104.865 ;
        RECT 212.725 104.720 213.440 104.890 ;
        RECT 212.725 103.790 213.055 104.550 ;
        RECT 213.270 103.960 213.440 104.720 ;
        RECT 213.700 103.790 213.990 104.955 ;
        RECT 214.850 104.880 215.370 105.420 ;
        RECT 214.160 103.790 215.370 104.880 ;
        RECT 215.545 103.790 215.805 104.940 ;
        RECT 215.980 104.865 216.150 105.595 ;
        RECT 216.405 105.430 216.575 105.620 ;
        RECT 216.320 105.100 216.575 105.430 ;
        RECT 216.405 104.890 216.575 105.100 ;
        RECT 216.855 105.070 217.210 105.440 ;
        RECT 217.380 105.070 217.735 105.440 ;
        RECT 218.015 105.430 218.185 105.620 ;
        RECT 218.355 105.595 218.610 106.170 ;
        RECT 218.015 105.100 218.270 105.430 ;
        RECT 218.015 104.890 218.185 105.100 ;
        RECT 215.980 103.960 216.235 104.865 ;
        RECT 216.405 104.720 217.120 104.890 ;
        RECT 216.405 103.790 216.735 104.550 ;
        RECT 216.950 103.960 217.120 104.720 ;
        RECT 217.470 104.720 218.185 104.890 ;
        RECT 218.440 104.865 218.610 105.595 ;
        RECT 218.785 105.500 219.045 106.340 ;
        RECT 219.225 105.600 219.480 106.170 ;
        RECT 219.650 105.940 219.980 106.340 ;
        RECT 220.405 105.805 220.935 106.170 ;
        RECT 220.405 105.770 220.580 105.805 ;
        RECT 219.650 105.600 220.580 105.770 ;
        RECT 221.125 105.660 221.400 106.170 ;
        RECT 217.470 103.960 217.640 104.720 ;
        RECT 217.855 103.790 218.185 104.550 ;
        RECT 218.355 103.960 218.610 104.865 ;
        RECT 218.785 103.790 219.045 104.940 ;
        RECT 219.225 104.930 219.395 105.600 ;
        RECT 219.650 105.430 219.820 105.600 ;
        RECT 219.565 105.100 219.820 105.430 ;
        RECT 220.045 105.100 220.240 105.430 ;
        RECT 219.225 103.960 219.560 104.930 ;
        RECT 219.730 103.790 219.900 104.930 ;
        RECT 220.070 104.130 220.240 105.100 ;
        RECT 220.410 104.470 220.580 105.600 ;
        RECT 220.750 104.810 220.920 105.610 ;
        RECT 221.120 105.490 221.400 105.660 ;
        RECT 221.125 105.010 221.400 105.490 ;
        RECT 221.570 104.810 221.760 106.170 ;
        RECT 221.940 105.805 222.450 106.340 ;
        RECT 222.670 105.530 222.915 106.135 ;
        RECT 223.360 105.590 224.570 106.340 ;
        RECT 221.960 105.360 223.190 105.530 ;
        RECT 220.750 104.640 221.760 104.810 ;
        RECT 221.930 104.795 222.680 104.985 ;
        RECT 220.410 104.300 221.535 104.470 ;
        RECT 221.930 104.130 222.100 104.795 ;
        RECT 222.850 104.550 223.190 105.360 ;
        RECT 223.360 105.050 223.880 105.590 ;
        RECT 224.745 105.500 225.005 106.340 ;
        RECT 225.180 105.595 225.435 106.170 ;
        RECT 225.605 105.960 225.935 106.340 ;
        RECT 226.150 105.790 226.320 106.170 ;
        RECT 225.605 105.620 226.320 105.790 ;
        RECT 224.050 104.880 224.570 105.420 ;
        RECT 220.070 103.960 222.100 104.130 ;
        RECT 222.270 103.790 222.440 104.550 ;
        RECT 222.675 104.140 223.190 104.550 ;
        RECT 223.360 103.790 224.570 104.880 ;
        RECT 224.745 103.790 225.005 104.940 ;
        RECT 225.180 104.865 225.350 105.595 ;
        RECT 225.605 105.430 225.775 105.620 ;
        RECT 226.580 105.615 226.870 106.340 ;
        RECT 227.040 105.600 227.425 106.170 ;
        RECT 227.595 105.880 227.920 106.340 ;
        RECT 228.440 105.710 228.720 106.170 ;
        RECT 225.520 105.100 225.775 105.430 ;
        RECT 225.605 104.890 225.775 105.100 ;
        RECT 226.055 105.070 226.410 105.440 ;
        RECT 225.180 103.960 225.435 104.865 ;
        RECT 225.605 104.720 226.320 104.890 ;
        RECT 225.605 103.790 225.935 104.550 ;
        RECT 226.150 103.960 226.320 104.720 ;
        RECT 226.580 103.790 226.870 104.955 ;
        RECT 227.040 104.930 227.320 105.600 ;
        RECT 227.595 105.540 228.720 105.710 ;
        RECT 227.595 105.430 228.045 105.540 ;
        RECT 227.490 105.100 228.045 105.430 ;
        RECT 228.910 105.370 229.310 106.170 ;
        RECT 229.710 105.880 229.980 106.340 ;
        RECT 230.150 105.710 230.435 106.170 ;
        RECT 227.040 103.960 227.425 104.930 ;
        RECT 227.595 104.640 228.045 105.100 ;
        RECT 228.215 104.810 229.310 105.370 ;
        RECT 227.595 104.420 228.720 104.640 ;
        RECT 227.595 103.790 227.920 104.250 ;
        RECT 228.440 103.960 228.720 104.420 ;
        RECT 228.910 103.960 229.310 104.810 ;
        RECT 229.480 105.540 230.435 105.710 ;
        RECT 229.480 104.640 229.690 105.540 ;
        RECT 231.185 105.500 231.445 106.340 ;
        RECT 231.620 105.595 231.875 106.170 ;
        RECT 232.045 105.960 232.375 106.340 ;
        RECT 232.590 105.790 232.760 106.170 ;
        RECT 232.045 105.620 232.760 105.790 ;
        RECT 229.860 104.810 230.550 105.370 ;
        RECT 229.480 104.420 230.435 104.640 ;
        RECT 229.710 103.790 229.980 104.250 ;
        RECT 230.150 103.960 230.435 104.420 ;
        RECT 231.185 103.790 231.445 104.940 ;
        RECT 231.620 104.865 231.790 105.595 ;
        RECT 232.045 105.430 232.215 105.620 ;
        RECT 233.485 105.500 233.745 106.340 ;
        RECT 233.920 105.595 234.175 106.170 ;
        RECT 234.345 105.960 234.675 106.340 ;
        RECT 234.890 105.790 235.060 106.170 ;
        RECT 234.345 105.620 235.060 105.790 ;
        RECT 231.960 105.100 232.215 105.430 ;
        RECT 232.045 104.890 232.215 105.100 ;
        RECT 232.495 105.070 232.850 105.440 ;
        RECT 231.620 103.960 231.875 104.865 ;
        RECT 232.045 104.720 232.760 104.890 ;
        RECT 232.045 103.790 232.375 104.550 ;
        RECT 232.590 103.960 232.760 104.720 ;
        RECT 233.485 103.790 233.745 104.940 ;
        RECT 233.920 104.865 234.090 105.595 ;
        RECT 234.345 105.430 234.515 105.620 ;
        RECT 235.785 105.500 236.045 106.340 ;
        RECT 236.220 105.595 236.475 106.170 ;
        RECT 236.645 105.960 236.975 106.340 ;
        RECT 237.190 105.790 237.360 106.170 ;
        RECT 236.645 105.620 237.360 105.790 ;
        RECT 234.260 105.100 234.515 105.430 ;
        RECT 234.345 104.890 234.515 105.100 ;
        RECT 234.795 105.070 235.150 105.440 ;
        RECT 233.920 103.960 234.175 104.865 ;
        RECT 234.345 104.720 235.060 104.890 ;
        RECT 234.345 103.790 234.675 104.550 ;
        RECT 234.890 103.960 235.060 104.720 ;
        RECT 235.785 103.790 236.045 104.940 ;
        RECT 236.220 104.865 236.390 105.595 ;
        RECT 236.645 105.430 236.815 105.620 ;
        RECT 237.625 105.500 237.885 106.340 ;
        RECT 238.060 105.595 238.315 106.170 ;
        RECT 238.485 105.960 238.815 106.340 ;
        RECT 239.030 105.790 239.200 106.170 ;
        RECT 238.485 105.620 239.200 105.790 ;
        RECT 236.560 105.100 236.815 105.430 ;
        RECT 236.645 104.890 236.815 105.100 ;
        RECT 237.095 105.070 237.450 105.440 ;
        RECT 236.220 103.960 236.475 104.865 ;
        RECT 236.645 104.720 237.360 104.890 ;
        RECT 236.645 103.790 236.975 104.550 ;
        RECT 237.190 103.960 237.360 104.720 ;
        RECT 237.625 103.790 237.885 104.940 ;
        RECT 238.060 104.865 238.230 105.595 ;
        RECT 238.485 105.430 238.655 105.620 ;
        RECT 239.460 105.615 239.750 106.340 ;
        RECT 240.385 105.600 240.640 106.170 ;
        RECT 240.810 105.940 241.140 106.340 ;
        RECT 241.565 105.805 242.095 106.170 ;
        RECT 242.285 106.000 242.560 106.170 ;
        RECT 242.280 105.830 242.560 106.000 ;
        RECT 241.565 105.770 241.740 105.805 ;
        RECT 240.810 105.600 241.740 105.770 ;
        RECT 238.400 105.100 238.655 105.430 ;
        RECT 238.485 104.890 238.655 105.100 ;
        RECT 238.935 105.070 239.290 105.440 ;
        RECT 238.060 103.960 238.315 104.865 ;
        RECT 238.485 104.720 239.200 104.890 ;
        RECT 238.485 103.790 238.815 104.550 ;
        RECT 239.030 103.960 239.200 104.720 ;
        RECT 239.460 103.790 239.750 104.955 ;
        RECT 240.385 104.930 240.555 105.600 ;
        RECT 240.810 105.430 240.980 105.600 ;
        RECT 240.725 105.100 240.980 105.430 ;
        RECT 241.205 105.100 241.400 105.430 ;
        RECT 240.385 103.960 240.720 104.930 ;
        RECT 240.890 103.790 241.060 104.930 ;
        RECT 241.230 104.130 241.400 105.100 ;
        RECT 241.570 104.470 241.740 105.600 ;
        RECT 241.910 104.810 242.080 105.610 ;
        RECT 242.285 105.010 242.560 105.830 ;
        RECT 242.730 104.810 242.920 106.170 ;
        RECT 243.100 105.805 243.610 106.340 ;
        RECT 243.830 105.530 244.075 106.135 ;
        RECT 244.635 105.710 244.920 106.170 ;
        RECT 245.090 105.880 245.360 106.340 ;
        RECT 244.635 105.540 245.590 105.710 ;
        RECT 243.120 105.360 244.350 105.530 ;
        RECT 241.910 104.640 242.920 104.810 ;
        RECT 243.090 104.795 243.840 104.985 ;
        RECT 241.570 104.300 242.695 104.470 ;
        RECT 243.090 104.130 243.260 104.795 ;
        RECT 244.010 104.550 244.350 105.360 ;
        RECT 244.520 104.810 245.210 105.370 ;
        RECT 245.380 104.640 245.590 105.540 ;
        RECT 241.230 103.960 243.260 104.130 ;
        RECT 243.430 103.790 243.600 104.550 ;
        RECT 243.835 104.140 244.350 104.550 ;
        RECT 244.635 104.420 245.590 104.640 ;
        RECT 245.760 105.370 246.160 106.170 ;
        RECT 246.350 105.710 246.630 106.170 ;
        RECT 247.150 105.880 247.475 106.340 ;
        RECT 246.350 105.540 247.475 105.710 ;
        RECT 247.645 105.600 248.030 106.170 ;
        RECT 247.025 105.430 247.475 105.540 ;
        RECT 245.760 104.810 246.855 105.370 ;
        RECT 247.025 105.100 247.580 105.430 ;
        RECT 244.635 103.960 244.920 104.420 ;
        RECT 245.090 103.790 245.360 104.250 ;
        RECT 245.760 103.960 246.160 104.810 ;
        RECT 247.025 104.640 247.475 105.100 ;
        RECT 247.750 104.930 248.030 105.600 ;
        RECT 246.350 104.420 247.475 104.640 ;
        RECT 246.350 103.960 246.630 104.420 ;
        RECT 247.150 103.790 247.475 104.250 ;
        RECT 247.645 103.960 248.030 104.930 ;
        RECT 248.200 105.600 248.585 106.170 ;
        RECT 248.755 105.880 249.080 106.340 ;
        RECT 249.600 105.710 249.880 106.170 ;
        RECT 248.200 104.930 248.480 105.600 ;
        RECT 248.755 105.540 249.880 105.710 ;
        RECT 248.755 105.430 249.205 105.540 ;
        RECT 248.650 105.100 249.205 105.430 ;
        RECT 250.070 105.370 250.470 106.170 ;
        RECT 250.870 105.880 251.140 106.340 ;
        RECT 251.310 105.710 251.595 106.170 ;
        RECT 248.200 103.960 248.585 104.930 ;
        RECT 248.755 104.640 249.205 105.100 ;
        RECT 249.375 104.810 250.470 105.370 ;
        RECT 248.755 104.420 249.880 104.640 ;
        RECT 248.755 103.790 249.080 104.250 ;
        RECT 249.600 103.960 249.880 104.420 ;
        RECT 250.070 103.960 250.470 104.810 ;
        RECT 250.640 105.540 251.595 105.710 ;
        RECT 252.340 105.615 252.630 106.340 ;
        RECT 253.720 105.600 254.105 106.170 ;
        RECT 254.275 105.880 254.600 106.340 ;
        RECT 255.120 105.710 255.400 106.170 ;
        RECT 250.640 104.640 250.850 105.540 ;
        RECT 251.020 104.810 251.710 105.370 ;
        RECT 250.640 104.420 251.595 104.640 ;
        RECT 250.870 103.790 251.140 104.250 ;
        RECT 251.310 103.960 251.595 104.420 ;
        RECT 252.340 103.790 252.630 104.955 ;
        RECT 253.720 104.930 254.000 105.600 ;
        RECT 254.275 105.540 255.400 105.710 ;
        RECT 254.275 105.430 254.725 105.540 ;
        RECT 254.170 105.100 254.725 105.430 ;
        RECT 255.590 105.370 255.990 106.170 ;
        RECT 256.390 105.880 256.660 106.340 ;
        RECT 256.830 105.710 257.115 106.170 ;
        RECT 253.720 103.960 254.105 104.930 ;
        RECT 254.275 104.640 254.725 105.100 ;
        RECT 254.895 104.810 255.990 105.370 ;
        RECT 254.275 104.420 255.400 104.640 ;
        RECT 254.275 103.790 254.600 104.250 ;
        RECT 255.120 103.960 255.400 104.420 ;
        RECT 255.590 103.960 255.990 104.810 ;
        RECT 256.160 105.540 257.115 105.710 ;
        RECT 257.490 105.790 257.660 106.170 ;
        RECT 257.875 105.960 258.205 106.340 ;
        RECT 257.490 105.620 258.205 105.790 ;
        RECT 256.160 104.640 256.370 105.540 ;
        RECT 256.540 104.810 257.230 105.370 ;
        RECT 257.400 105.070 257.755 105.440 ;
        RECT 258.035 105.430 258.205 105.620 ;
        RECT 258.375 105.595 258.630 106.170 ;
        RECT 258.035 105.100 258.290 105.430 ;
        RECT 258.035 104.890 258.205 105.100 ;
        RECT 257.490 104.720 258.205 104.890 ;
        RECT 258.460 104.865 258.630 105.595 ;
        RECT 258.805 105.500 259.065 106.340 ;
        RECT 259.245 105.500 259.505 106.340 ;
        RECT 259.680 105.595 259.935 106.170 ;
        RECT 260.105 105.960 260.435 106.340 ;
        RECT 260.650 105.790 260.820 106.170 ;
        RECT 260.105 105.620 260.820 105.790 ;
        RECT 256.160 104.420 257.115 104.640 ;
        RECT 256.390 103.790 256.660 104.250 ;
        RECT 256.830 103.960 257.115 104.420 ;
        RECT 257.490 103.960 257.660 104.720 ;
        RECT 257.875 103.790 258.205 104.550 ;
        RECT 258.375 103.960 258.630 104.865 ;
        RECT 258.805 103.790 259.065 104.940 ;
        RECT 259.245 103.790 259.505 104.940 ;
        RECT 259.680 104.865 259.850 105.595 ;
        RECT 260.105 105.430 260.275 105.620 ;
        RECT 261.085 105.500 261.345 106.340 ;
        RECT 261.520 105.595 261.775 106.170 ;
        RECT 261.945 105.960 262.275 106.340 ;
        RECT 262.490 105.790 262.660 106.170 ;
        RECT 261.945 105.620 262.660 105.790 ;
        RECT 260.020 105.100 260.275 105.430 ;
        RECT 260.105 104.890 260.275 105.100 ;
        RECT 260.555 105.070 260.910 105.440 ;
        RECT 259.680 103.960 259.935 104.865 ;
        RECT 260.105 104.720 260.820 104.890 ;
        RECT 260.105 103.790 260.435 104.550 ;
        RECT 260.650 103.960 260.820 104.720 ;
        RECT 261.085 103.790 261.345 104.940 ;
        RECT 261.520 104.865 261.690 105.595 ;
        RECT 261.945 105.430 262.115 105.620 ;
        RECT 262.925 105.500 263.185 106.340 ;
        RECT 263.360 105.595 263.615 106.170 ;
        RECT 263.785 105.960 264.115 106.340 ;
        RECT 264.330 105.790 264.500 106.170 ;
        RECT 263.785 105.620 264.500 105.790 ;
        RECT 261.860 105.100 262.115 105.430 ;
        RECT 261.945 104.890 262.115 105.100 ;
        RECT 262.395 105.070 262.750 105.440 ;
        RECT 261.520 103.960 261.775 104.865 ;
        RECT 261.945 104.720 262.660 104.890 ;
        RECT 261.945 103.790 262.275 104.550 ;
        RECT 262.490 103.960 262.660 104.720 ;
        RECT 262.925 103.790 263.185 104.940 ;
        RECT 263.360 104.865 263.530 105.595 ;
        RECT 263.785 105.430 263.955 105.620 ;
        RECT 265.220 105.615 265.510 106.340 ;
        RECT 265.685 105.500 265.945 106.340 ;
        RECT 266.120 105.595 266.375 106.170 ;
        RECT 266.545 105.960 266.875 106.340 ;
        RECT 267.090 105.790 267.260 106.170 ;
        RECT 266.545 105.620 267.260 105.790 ;
        RECT 263.700 105.100 263.955 105.430 ;
        RECT 263.785 104.890 263.955 105.100 ;
        RECT 264.235 105.070 264.590 105.440 ;
        RECT 263.360 103.960 263.615 104.865 ;
        RECT 263.785 104.720 264.500 104.890 ;
        RECT 263.785 103.790 264.115 104.550 ;
        RECT 264.330 103.960 264.500 104.720 ;
        RECT 265.220 103.790 265.510 104.955 ;
        RECT 265.685 103.790 265.945 104.940 ;
        RECT 266.120 104.865 266.290 105.595 ;
        RECT 266.545 105.430 266.715 105.620 ;
        RECT 267.525 105.500 267.785 106.340 ;
        RECT 267.960 105.595 268.215 106.170 ;
        RECT 268.385 105.960 268.715 106.340 ;
        RECT 268.930 105.790 269.100 106.170 ;
        RECT 268.385 105.620 269.100 105.790 ;
        RECT 269.475 105.710 269.760 106.170 ;
        RECT 269.930 105.880 270.200 106.340 ;
        RECT 266.460 105.100 266.715 105.430 ;
        RECT 266.545 104.890 266.715 105.100 ;
        RECT 266.995 105.070 267.350 105.440 ;
        RECT 266.120 103.960 266.375 104.865 ;
        RECT 266.545 104.720 267.260 104.890 ;
        RECT 266.545 103.790 266.875 104.550 ;
        RECT 267.090 103.960 267.260 104.720 ;
        RECT 267.525 103.790 267.785 104.940 ;
        RECT 267.960 104.865 268.130 105.595 ;
        RECT 268.385 105.430 268.555 105.620 ;
        RECT 269.475 105.540 270.430 105.710 ;
        RECT 268.300 105.100 268.555 105.430 ;
        RECT 268.385 104.890 268.555 105.100 ;
        RECT 268.835 105.070 269.190 105.440 ;
        RECT 267.960 103.960 268.215 104.865 ;
        RECT 268.385 104.720 269.100 104.890 ;
        RECT 269.360 104.810 270.050 105.370 ;
        RECT 268.385 103.790 268.715 104.550 ;
        RECT 268.930 103.960 269.100 104.720 ;
        RECT 270.220 104.640 270.430 105.540 ;
        RECT 269.475 104.420 270.430 104.640 ;
        RECT 270.600 105.370 271.000 106.170 ;
        RECT 271.190 105.710 271.470 106.170 ;
        RECT 271.990 105.880 272.315 106.340 ;
        RECT 271.190 105.540 272.315 105.710 ;
        RECT 272.485 105.600 272.870 106.170 ;
        RECT 271.865 105.430 272.315 105.540 ;
        RECT 270.600 104.810 271.695 105.370 ;
        RECT 271.865 105.100 272.420 105.430 ;
        RECT 269.475 103.960 269.760 104.420 ;
        RECT 269.930 103.790 270.200 104.250 ;
        RECT 270.600 103.960 271.000 104.810 ;
        RECT 271.865 104.640 272.315 105.100 ;
        RECT 272.590 104.930 272.870 105.600 ;
        RECT 273.045 105.500 273.305 106.340 ;
        RECT 273.480 105.595 273.735 106.170 ;
        RECT 273.905 105.960 274.235 106.340 ;
        RECT 274.450 105.790 274.620 106.170 ;
        RECT 273.905 105.620 274.620 105.790 ;
        RECT 274.970 105.790 275.140 106.170 ;
        RECT 275.355 105.960 275.685 106.340 ;
        RECT 274.970 105.620 275.685 105.790 ;
        RECT 271.190 104.420 272.315 104.640 ;
        RECT 271.190 103.960 271.470 104.420 ;
        RECT 271.990 103.790 272.315 104.250 ;
        RECT 272.485 103.960 272.870 104.930 ;
        RECT 273.045 103.790 273.305 104.940 ;
        RECT 273.480 104.865 273.650 105.595 ;
        RECT 273.905 105.430 274.075 105.620 ;
        RECT 273.820 105.100 274.075 105.430 ;
        RECT 273.905 104.890 274.075 105.100 ;
        RECT 274.355 105.070 274.710 105.440 ;
        RECT 274.880 105.070 275.235 105.440 ;
        RECT 275.515 105.430 275.685 105.620 ;
        RECT 275.855 105.595 276.110 106.170 ;
        RECT 275.515 105.100 275.770 105.430 ;
        RECT 275.515 104.890 275.685 105.100 ;
        RECT 273.480 103.960 273.735 104.865 ;
        RECT 273.905 104.720 274.620 104.890 ;
        RECT 273.905 103.790 274.235 104.550 ;
        RECT 274.450 103.960 274.620 104.720 ;
        RECT 274.970 104.720 275.685 104.890 ;
        RECT 275.940 104.865 276.110 105.595 ;
        RECT 276.285 105.500 276.545 106.340 ;
        RECT 276.720 105.590 277.930 106.340 ;
        RECT 278.100 105.615 278.390 106.340 ;
        RECT 276.720 105.050 277.240 105.590 ;
        RECT 278.565 105.500 278.825 106.340 ;
        RECT 279.000 105.595 279.255 106.170 ;
        RECT 279.425 105.960 279.755 106.340 ;
        RECT 279.970 105.790 280.140 106.170 ;
        RECT 279.425 105.620 280.140 105.790 ;
        RECT 274.970 103.960 275.140 104.720 ;
        RECT 275.355 103.790 275.685 104.550 ;
        RECT 275.855 103.960 276.110 104.865 ;
        RECT 276.285 103.790 276.545 104.940 ;
        RECT 277.410 104.880 277.930 105.420 ;
        RECT 276.720 103.790 277.930 104.880 ;
        RECT 278.100 103.790 278.390 104.955 ;
        RECT 278.565 103.790 278.825 104.940 ;
        RECT 279.000 104.865 279.170 105.595 ;
        RECT 279.425 105.430 279.595 105.620 ;
        RECT 280.405 105.500 280.665 106.340 ;
        RECT 280.840 105.595 281.095 106.170 ;
        RECT 281.265 105.960 281.595 106.340 ;
        RECT 281.810 105.790 281.980 106.170 ;
        RECT 281.265 105.620 281.980 105.790 ;
        RECT 279.340 105.100 279.595 105.430 ;
        RECT 279.425 104.890 279.595 105.100 ;
        RECT 279.875 105.070 280.230 105.440 ;
        RECT 279.000 103.960 279.255 104.865 ;
        RECT 279.425 104.720 280.140 104.890 ;
        RECT 279.425 103.790 279.755 104.550 ;
        RECT 279.970 103.960 280.140 104.720 ;
        RECT 280.405 103.790 280.665 104.940 ;
        RECT 280.840 104.865 281.010 105.595 ;
        RECT 281.265 105.430 281.435 105.620 ;
        RECT 282.245 105.500 282.505 106.340 ;
        RECT 282.680 105.595 282.935 106.170 ;
        RECT 283.105 105.960 283.435 106.340 ;
        RECT 283.650 105.790 283.820 106.170 ;
        RECT 283.105 105.620 283.820 105.790 ;
        RECT 281.180 105.100 281.435 105.430 ;
        RECT 281.265 104.890 281.435 105.100 ;
        RECT 281.715 105.070 282.070 105.440 ;
        RECT 280.840 103.960 281.095 104.865 ;
        RECT 281.265 104.720 281.980 104.890 ;
        RECT 281.265 103.790 281.595 104.550 ;
        RECT 281.810 103.960 281.980 104.720 ;
        RECT 282.245 103.790 282.505 104.940 ;
        RECT 282.680 104.865 282.850 105.595 ;
        RECT 283.105 105.430 283.275 105.620 ;
        RECT 284.085 105.500 284.345 106.340 ;
        RECT 284.520 105.595 284.775 106.170 ;
        RECT 284.945 105.960 285.275 106.340 ;
        RECT 285.490 105.790 285.660 106.170 ;
        RECT 284.945 105.620 285.660 105.790 ;
        RECT 283.020 105.100 283.275 105.430 ;
        RECT 283.105 104.890 283.275 105.100 ;
        RECT 283.555 105.070 283.910 105.440 ;
        RECT 282.680 103.960 282.935 104.865 ;
        RECT 283.105 104.720 283.820 104.890 ;
        RECT 283.105 103.790 283.435 104.550 ;
        RECT 283.650 103.960 283.820 104.720 ;
        RECT 284.085 103.790 284.345 104.940 ;
        RECT 284.520 104.865 284.690 105.595 ;
        RECT 284.945 105.430 285.115 105.620 ;
        RECT 285.925 105.500 286.185 106.340 ;
        RECT 286.360 105.595 286.615 106.170 ;
        RECT 286.785 105.960 287.115 106.340 ;
        RECT 287.330 105.790 287.500 106.170 ;
        RECT 286.785 105.620 287.500 105.790 ;
        RECT 284.860 105.100 285.115 105.430 ;
        RECT 284.945 104.890 285.115 105.100 ;
        RECT 285.395 105.070 285.750 105.440 ;
        RECT 284.520 103.960 284.775 104.865 ;
        RECT 284.945 104.720 285.660 104.890 ;
        RECT 284.945 103.790 285.275 104.550 ;
        RECT 285.490 103.960 285.660 104.720 ;
        RECT 285.925 103.790 286.185 104.940 ;
        RECT 286.360 104.865 286.530 105.595 ;
        RECT 286.785 105.430 286.955 105.620 ;
        RECT 287.765 105.500 288.025 106.340 ;
        RECT 288.200 105.595 288.455 106.170 ;
        RECT 288.625 105.960 288.955 106.340 ;
        RECT 289.170 105.790 289.340 106.170 ;
        RECT 288.625 105.620 289.340 105.790 ;
        RECT 286.700 105.100 286.955 105.430 ;
        RECT 286.785 104.890 286.955 105.100 ;
        RECT 287.235 105.070 287.590 105.440 ;
        RECT 286.360 103.960 286.615 104.865 ;
        RECT 286.785 104.720 287.500 104.890 ;
        RECT 286.785 103.790 287.115 104.550 ;
        RECT 287.330 103.960 287.500 104.720 ;
        RECT 287.765 103.790 288.025 104.940 ;
        RECT 288.200 104.865 288.370 105.595 ;
        RECT 288.625 105.430 288.795 105.620 ;
        RECT 289.600 105.590 290.810 106.340 ;
        RECT 290.980 105.615 291.270 106.340 ;
        RECT 288.540 105.100 288.795 105.430 ;
        RECT 288.625 104.890 288.795 105.100 ;
        RECT 289.075 105.070 289.430 105.440 ;
        RECT 289.600 105.050 290.120 105.590 ;
        RECT 291.445 105.500 291.705 106.340 ;
        RECT 291.880 105.595 292.135 106.170 ;
        RECT 292.305 105.960 292.635 106.340 ;
        RECT 292.850 105.790 293.020 106.170 ;
        RECT 292.305 105.620 293.020 105.790 ;
        RECT 288.200 103.960 288.455 104.865 ;
        RECT 288.625 104.720 289.340 104.890 ;
        RECT 290.290 104.880 290.810 105.420 ;
        RECT 288.625 103.790 288.955 104.550 ;
        RECT 289.170 103.960 289.340 104.720 ;
        RECT 289.600 103.790 290.810 104.880 ;
        RECT 290.980 103.790 291.270 104.955 ;
        RECT 291.445 103.790 291.705 104.940 ;
        RECT 291.880 104.865 292.050 105.595 ;
        RECT 292.305 105.430 292.475 105.620 ;
        RECT 293.280 105.590 294.490 106.340 ;
        RECT 294.665 105.790 294.920 106.080 ;
        RECT 295.090 105.960 295.420 106.340 ;
        RECT 294.665 105.620 295.415 105.790 ;
        RECT 292.220 105.100 292.475 105.430 ;
        RECT 292.305 104.890 292.475 105.100 ;
        RECT 292.755 105.070 293.110 105.440 ;
        RECT 293.280 105.050 293.800 105.590 ;
        RECT 291.880 103.960 292.135 104.865 ;
        RECT 292.305 104.720 293.020 104.890 ;
        RECT 293.970 104.880 294.490 105.420 ;
        RECT 292.305 103.790 292.635 104.550 ;
        RECT 292.850 103.960 293.020 104.720 ;
        RECT 293.280 103.790 294.490 104.880 ;
        RECT 294.665 104.800 295.015 105.450 ;
        RECT 295.185 104.630 295.415 105.620 ;
        RECT 294.665 104.460 295.415 104.630 ;
        RECT 294.665 103.960 294.920 104.460 ;
        RECT 295.090 103.790 295.420 104.290 ;
        RECT 295.590 103.960 295.760 106.080 ;
        RECT 296.120 105.980 296.450 106.340 ;
        RECT 296.620 105.950 297.115 106.120 ;
        RECT 297.320 105.950 298.175 106.120 ;
        RECT 295.990 104.760 296.450 105.810 ;
        RECT 295.930 103.975 296.255 104.760 ;
        RECT 296.620 104.590 296.790 105.950 ;
        RECT 296.960 105.040 297.310 105.660 ;
        RECT 297.480 105.440 297.835 105.660 ;
        RECT 297.480 104.850 297.650 105.440 ;
        RECT 298.005 105.240 298.175 105.950 ;
        RECT 299.050 105.880 299.380 106.340 ;
        RECT 299.590 105.980 299.940 106.150 ;
        RECT 298.380 105.410 299.170 105.660 ;
        RECT 299.590 105.590 299.850 105.980 ;
        RECT 300.160 105.890 301.110 106.170 ;
        RECT 301.280 105.900 301.470 106.340 ;
        RECT 301.640 105.960 302.710 106.130 ;
        RECT 299.340 105.240 299.510 105.420 ;
        RECT 296.620 104.420 297.015 104.590 ;
        RECT 297.185 104.460 297.650 104.850 ;
        RECT 297.820 105.070 299.510 105.240 ;
        RECT 296.845 104.290 297.015 104.420 ;
        RECT 297.820 104.290 297.990 105.070 ;
        RECT 299.680 104.900 299.850 105.590 ;
        RECT 298.350 104.730 299.850 104.900 ;
        RECT 300.040 104.930 300.250 105.720 ;
        RECT 300.420 105.100 300.770 105.720 ;
        RECT 300.940 105.110 301.110 105.890 ;
        RECT 301.640 105.730 301.810 105.960 ;
        RECT 301.280 105.560 301.810 105.730 ;
        RECT 301.280 105.280 301.500 105.560 ;
        RECT 301.980 105.390 302.220 105.790 ;
        RECT 300.940 104.940 301.345 105.110 ;
        RECT 301.680 105.020 302.220 105.390 ;
        RECT 302.390 105.605 302.710 105.960 ;
        RECT 302.955 105.880 303.260 106.340 ;
        RECT 303.430 105.630 303.685 106.160 ;
        RECT 302.390 105.430 302.715 105.605 ;
        RECT 302.390 105.130 303.305 105.430 ;
        RECT 302.565 105.100 303.305 105.130 ;
        RECT 300.040 104.770 300.715 104.930 ;
        RECT 301.175 104.850 301.345 104.940 ;
        RECT 300.040 104.760 301.005 104.770 ;
        RECT 299.680 104.590 299.850 104.730 ;
        RECT 296.425 103.790 296.675 104.250 ;
        RECT 296.845 103.960 297.095 104.290 ;
        RECT 297.310 103.960 297.990 104.290 ;
        RECT 298.160 104.390 299.235 104.560 ;
        RECT 299.680 104.420 300.240 104.590 ;
        RECT 300.545 104.470 301.005 104.760 ;
        RECT 301.175 104.680 302.395 104.850 ;
        RECT 298.160 104.050 298.330 104.390 ;
        RECT 298.565 103.790 298.895 104.220 ;
        RECT 299.065 104.050 299.235 104.390 ;
        RECT 299.530 103.790 299.900 104.250 ;
        RECT 300.070 103.960 300.240 104.420 ;
        RECT 301.175 104.300 301.345 104.680 ;
        RECT 302.565 104.510 302.735 105.100 ;
        RECT 303.475 104.980 303.685 105.630 ;
        RECT 303.860 105.615 304.150 106.340 ;
        RECT 304.410 105.790 304.580 106.170 ;
        RECT 304.795 105.960 305.125 106.340 ;
        RECT 304.410 105.620 305.125 105.790 ;
        RECT 304.320 105.070 304.675 105.440 ;
        RECT 304.955 105.430 305.125 105.620 ;
        RECT 305.295 105.595 305.550 106.170 ;
        RECT 304.955 105.100 305.210 105.430 ;
        RECT 300.475 103.960 301.345 104.300 ;
        RECT 301.935 104.340 302.735 104.510 ;
        RECT 301.515 103.790 301.765 104.250 ;
        RECT 301.935 104.050 302.105 104.340 ;
        RECT 302.285 103.790 302.615 104.170 ;
        RECT 302.955 103.790 303.260 104.930 ;
        RECT 303.430 104.100 303.685 104.980 ;
        RECT 303.860 103.790 304.150 104.955 ;
        RECT 304.955 104.890 305.125 105.100 ;
        RECT 304.410 104.720 305.125 104.890 ;
        RECT 305.380 104.865 305.550 105.595 ;
        RECT 305.725 105.500 305.985 106.340 ;
        RECT 306.250 105.790 306.420 106.170 ;
        RECT 306.635 105.960 306.965 106.340 ;
        RECT 306.250 105.620 306.965 105.790 ;
        RECT 306.160 105.070 306.515 105.440 ;
        RECT 306.795 105.430 306.965 105.620 ;
        RECT 307.135 105.595 307.390 106.170 ;
        RECT 306.795 105.100 307.050 105.430 ;
        RECT 304.410 103.960 304.580 104.720 ;
        RECT 304.795 103.790 305.125 104.550 ;
        RECT 305.295 103.960 305.550 104.865 ;
        RECT 305.725 103.790 305.985 104.940 ;
        RECT 306.795 104.890 306.965 105.100 ;
        RECT 306.250 104.720 306.965 104.890 ;
        RECT 307.220 104.865 307.390 105.595 ;
        RECT 307.565 105.500 307.825 106.340 ;
        RECT 308.090 105.790 308.260 106.170 ;
        RECT 308.475 105.960 308.805 106.340 ;
        RECT 308.090 105.620 308.805 105.790 ;
        RECT 308.000 105.070 308.355 105.440 ;
        RECT 308.635 105.430 308.805 105.620 ;
        RECT 308.975 105.595 309.230 106.170 ;
        RECT 308.635 105.100 308.890 105.430 ;
        RECT 306.250 103.960 306.420 104.720 ;
        RECT 306.635 103.790 306.965 104.550 ;
        RECT 307.135 103.960 307.390 104.865 ;
        RECT 307.565 103.790 307.825 104.940 ;
        RECT 308.635 104.890 308.805 105.100 ;
        RECT 308.090 104.720 308.805 104.890 ;
        RECT 309.060 104.865 309.230 105.595 ;
        RECT 309.405 105.500 309.665 106.340 ;
        RECT 309.840 105.590 311.050 106.340 ;
        RECT 308.090 103.960 308.260 104.720 ;
        RECT 308.475 103.790 308.805 104.550 ;
        RECT 308.975 103.960 309.230 104.865 ;
        RECT 309.405 103.790 309.665 104.940 ;
        RECT 309.840 104.880 310.360 105.420 ;
        RECT 310.530 105.050 311.050 105.590 ;
        RECT 309.840 103.790 311.050 104.880 ;
        RECT 162.095 103.620 311.135 103.790 ;
        RECT 162.180 102.530 163.390 103.620 ;
        RECT 162.180 101.820 162.700 102.360 ;
        RECT 162.870 101.990 163.390 102.530 ;
        RECT 164.025 102.470 164.285 103.620 ;
        RECT 164.460 102.545 164.715 103.450 ;
        RECT 164.885 102.860 165.215 103.620 ;
        RECT 165.430 102.690 165.600 103.450 ;
        RECT 165.865 102.950 166.120 103.450 ;
        RECT 166.290 103.120 166.620 103.620 ;
        RECT 165.865 102.780 166.615 102.950 ;
        RECT 162.180 101.070 163.390 101.820 ;
        RECT 164.025 101.070 164.285 101.910 ;
        RECT 164.460 101.815 164.630 102.545 ;
        RECT 164.885 102.520 165.600 102.690 ;
        RECT 164.885 102.310 165.055 102.520 ;
        RECT 164.800 101.980 165.055 102.310 ;
        RECT 164.460 101.240 164.715 101.815 ;
        RECT 164.885 101.790 165.055 101.980 ;
        RECT 165.335 101.970 165.690 102.340 ;
        RECT 165.865 101.960 166.215 102.610 ;
        RECT 166.385 101.790 166.615 102.780 ;
        RECT 164.885 101.620 165.600 101.790 ;
        RECT 164.885 101.070 165.215 101.450 ;
        RECT 165.430 101.240 165.600 101.620 ;
        RECT 165.865 101.620 166.615 101.790 ;
        RECT 165.865 101.330 166.120 101.620 ;
        RECT 166.290 101.070 166.620 101.450 ;
        RECT 166.790 101.330 166.960 103.450 ;
        RECT 167.130 102.650 167.455 103.435 ;
        RECT 167.625 103.160 167.875 103.620 ;
        RECT 168.045 103.120 168.295 103.450 ;
        RECT 168.510 103.120 169.190 103.450 ;
        RECT 168.045 102.990 168.215 103.120 ;
        RECT 167.820 102.820 168.215 102.990 ;
        RECT 167.190 101.600 167.650 102.650 ;
        RECT 167.820 101.460 167.990 102.820 ;
        RECT 168.385 102.560 168.850 102.950 ;
        RECT 168.160 101.750 168.510 102.370 ;
        RECT 168.680 101.970 168.850 102.560 ;
        RECT 169.020 102.340 169.190 103.120 ;
        RECT 169.360 103.020 169.530 103.360 ;
        RECT 169.765 103.190 170.095 103.620 ;
        RECT 170.265 103.020 170.435 103.360 ;
        RECT 170.730 103.160 171.100 103.620 ;
        RECT 169.360 102.850 170.435 103.020 ;
        RECT 171.270 102.990 171.440 103.450 ;
        RECT 171.675 103.110 172.545 103.450 ;
        RECT 172.715 103.160 172.965 103.620 ;
        RECT 170.880 102.820 171.440 102.990 ;
        RECT 170.880 102.680 171.050 102.820 ;
        RECT 169.550 102.510 171.050 102.680 ;
        RECT 171.745 102.650 172.205 102.940 ;
        RECT 169.020 102.170 170.710 102.340 ;
        RECT 168.680 101.750 169.035 101.970 ;
        RECT 169.205 101.460 169.375 102.170 ;
        RECT 169.580 101.750 170.370 102.000 ;
        RECT 170.540 101.990 170.710 102.170 ;
        RECT 170.880 101.820 171.050 102.510 ;
        RECT 167.320 101.070 167.650 101.430 ;
        RECT 167.820 101.290 168.315 101.460 ;
        RECT 168.520 101.290 169.375 101.460 ;
        RECT 170.250 101.070 170.580 101.530 ;
        RECT 170.790 101.430 171.050 101.820 ;
        RECT 171.240 102.640 172.205 102.650 ;
        RECT 172.375 102.730 172.545 103.110 ;
        RECT 173.135 103.070 173.305 103.360 ;
        RECT 173.485 103.240 173.815 103.620 ;
        RECT 173.135 102.900 173.935 103.070 ;
        RECT 171.240 102.480 171.915 102.640 ;
        RECT 172.375 102.560 173.595 102.730 ;
        RECT 171.240 101.690 171.450 102.480 ;
        RECT 172.375 102.470 172.545 102.560 ;
        RECT 171.620 101.690 171.970 102.310 ;
        RECT 172.140 102.300 172.545 102.470 ;
        RECT 172.140 101.520 172.310 102.300 ;
        RECT 172.480 101.850 172.700 102.130 ;
        RECT 172.880 102.020 173.420 102.390 ;
        RECT 173.765 102.310 173.935 102.900 ;
        RECT 174.155 102.480 174.460 103.620 ;
        RECT 174.630 102.430 174.885 103.310 ;
        RECT 175.060 102.455 175.350 103.620 ;
        RECT 175.520 102.530 176.730 103.620 ;
        RECT 176.905 102.950 177.160 103.450 ;
        RECT 177.330 103.120 177.660 103.620 ;
        RECT 176.905 102.780 177.655 102.950 ;
        RECT 173.765 102.280 174.505 102.310 ;
        RECT 172.480 101.680 173.010 101.850 ;
        RECT 170.790 101.260 171.140 101.430 ;
        RECT 171.360 101.240 172.310 101.520 ;
        RECT 172.480 101.070 172.670 101.510 ;
        RECT 172.840 101.450 173.010 101.680 ;
        RECT 173.180 101.620 173.420 102.020 ;
        RECT 173.590 101.980 174.505 102.280 ;
        RECT 173.590 101.805 173.915 101.980 ;
        RECT 173.590 101.450 173.910 101.805 ;
        RECT 174.675 101.780 174.885 102.430 ;
        RECT 175.520 101.820 176.040 102.360 ;
        RECT 176.210 101.990 176.730 102.530 ;
        RECT 176.905 101.960 177.255 102.610 ;
        RECT 172.840 101.280 173.910 101.450 ;
        RECT 174.155 101.070 174.460 101.530 ;
        RECT 174.630 101.250 174.885 101.780 ;
        RECT 175.060 101.070 175.350 101.795 ;
        RECT 175.520 101.070 176.730 101.820 ;
        RECT 177.425 101.790 177.655 102.780 ;
        RECT 176.905 101.620 177.655 101.790 ;
        RECT 176.905 101.330 177.160 101.620 ;
        RECT 177.330 101.070 177.660 101.450 ;
        RECT 177.830 101.330 178.000 103.450 ;
        RECT 178.170 102.650 178.495 103.435 ;
        RECT 178.665 103.160 178.915 103.620 ;
        RECT 179.085 103.120 179.335 103.450 ;
        RECT 179.550 103.120 180.230 103.450 ;
        RECT 179.085 102.990 179.255 103.120 ;
        RECT 178.860 102.820 179.255 102.990 ;
        RECT 178.230 101.600 178.690 102.650 ;
        RECT 178.860 101.460 179.030 102.820 ;
        RECT 179.425 102.560 179.890 102.950 ;
        RECT 179.200 101.750 179.550 102.370 ;
        RECT 179.720 101.970 179.890 102.560 ;
        RECT 180.060 102.340 180.230 103.120 ;
        RECT 180.400 103.020 180.570 103.360 ;
        RECT 180.805 103.190 181.135 103.620 ;
        RECT 181.305 103.020 181.475 103.360 ;
        RECT 181.770 103.160 182.140 103.620 ;
        RECT 180.400 102.850 181.475 103.020 ;
        RECT 182.310 102.990 182.480 103.450 ;
        RECT 182.715 103.110 183.585 103.450 ;
        RECT 183.755 103.160 184.005 103.620 ;
        RECT 181.920 102.820 182.480 102.990 ;
        RECT 181.920 102.680 182.090 102.820 ;
        RECT 180.590 102.510 182.090 102.680 ;
        RECT 182.785 102.650 183.245 102.940 ;
        RECT 180.060 102.170 181.750 102.340 ;
        RECT 179.720 101.750 180.075 101.970 ;
        RECT 180.245 101.460 180.415 102.170 ;
        RECT 180.620 101.750 181.410 102.000 ;
        RECT 181.580 101.990 181.750 102.170 ;
        RECT 181.920 101.820 182.090 102.510 ;
        RECT 178.360 101.070 178.690 101.430 ;
        RECT 178.860 101.290 179.355 101.460 ;
        RECT 179.560 101.290 180.415 101.460 ;
        RECT 181.290 101.070 181.620 101.530 ;
        RECT 181.830 101.430 182.090 101.820 ;
        RECT 182.280 102.640 183.245 102.650 ;
        RECT 183.415 102.730 183.585 103.110 ;
        RECT 184.175 103.070 184.345 103.360 ;
        RECT 184.525 103.240 184.855 103.620 ;
        RECT 184.175 102.900 184.975 103.070 ;
        RECT 182.280 102.480 182.955 102.640 ;
        RECT 183.415 102.560 184.635 102.730 ;
        RECT 182.280 101.690 182.490 102.480 ;
        RECT 183.415 102.470 183.585 102.560 ;
        RECT 182.660 101.690 183.010 102.310 ;
        RECT 183.180 102.300 183.585 102.470 ;
        RECT 183.180 101.520 183.350 102.300 ;
        RECT 183.520 101.850 183.740 102.130 ;
        RECT 183.920 102.020 184.460 102.390 ;
        RECT 184.805 102.310 184.975 102.900 ;
        RECT 185.195 102.480 185.500 103.620 ;
        RECT 185.670 102.430 185.925 103.310 ;
        RECT 186.105 102.950 186.360 103.450 ;
        RECT 186.530 103.120 186.860 103.620 ;
        RECT 186.105 102.780 186.855 102.950 ;
        RECT 184.805 102.280 185.545 102.310 ;
        RECT 183.520 101.680 184.050 101.850 ;
        RECT 181.830 101.260 182.180 101.430 ;
        RECT 182.400 101.240 183.350 101.520 ;
        RECT 183.520 101.070 183.710 101.510 ;
        RECT 183.880 101.450 184.050 101.680 ;
        RECT 184.220 101.620 184.460 102.020 ;
        RECT 184.630 101.980 185.545 102.280 ;
        RECT 184.630 101.805 184.955 101.980 ;
        RECT 184.630 101.450 184.950 101.805 ;
        RECT 185.715 101.780 185.925 102.430 ;
        RECT 186.105 101.960 186.455 102.610 ;
        RECT 186.625 101.790 186.855 102.780 ;
        RECT 183.880 101.280 184.950 101.450 ;
        RECT 185.195 101.070 185.500 101.530 ;
        RECT 185.670 101.250 185.925 101.780 ;
        RECT 186.105 101.620 186.855 101.790 ;
        RECT 186.105 101.330 186.360 101.620 ;
        RECT 186.530 101.070 186.860 101.450 ;
        RECT 187.030 101.330 187.200 103.450 ;
        RECT 187.370 102.650 187.695 103.435 ;
        RECT 187.865 103.160 188.115 103.620 ;
        RECT 188.285 103.120 188.535 103.450 ;
        RECT 188.750 103.120 189.430 103.450 ;
        RECT 188.285 102.990 188.455 103.120 ;
        RECT 188.060 102.820 188.455 102.990 ;
        RECT 187.430 101.600 187.890 102.650 ;
        RECT 188.060 101.460 188.230 102.820 ;
        RECT 188.625 102.560 189.090 102.950 ;
        RECT 188.400 101.750 188.750 102.370 ;
        RECT 188.920 101.970 189.090 102.560 ;
        RECT 189.260 102.340 189.430 103.120 ;
        RECT 189.600 103.020 189.770 103.360 ;
        RECT 190.005 103.190 190.335 103.620 ;
        RECT 190.505 103.020 190.675 103.360 ;
        RECT 190.970 103.160 191.340 103.620 ;
        RECT 189.600 102.850 190.675 103.020 ;
        RECT 191.510 102.990 191.680 103.450 ;
        RECT 191.915 103.110 192.785 103.450 ;
        RECT 192.955 103.160 193.205 103.620 ;
        RECT 191.120 102.820 191.680 102.990 ;
        RECT 191.120 102.680 191.290 102.820 ;
        RECT 189.790 102.510 191.290 102.680 ;
        RECT 191.985 102.650 192.445 102.940 ;
        RECT 189.260 102.170 190.950 102.340 ;
        RECT 188.920 101.750 189.275 101.970 ;
        RECT 189.445 101.460 189.615 102.170 ;
        RECT 189.820 101.750 190.610 102.000 ;
        RECT 190.780 101.990 190.950 102.170 ;
        RECT 191.120 101.820 191.290 102.510 ;
        RECT 187.560 101.070 187.890 101.430 ;
        RECT 188.060 101.290 188.555 101.460 ;
        RECT 188.760 101.290 189.615 101.460 ;
        RECT 190.490 101.070 190.820 101.530 ;
        RECT 191.030 101.430 191.290 101.820 ;
        RECT 191.480 102.640 192.445 102.650 ;
        RECT 192.615 102.730 192.785 103.110 ;
        RECT 193.375 103.070 193.545 103.360 ;
        RECT 193.725 103.240 194.055 103.620 ;
        RECT 193.375 102.900 194.175 103.070 ;
        RECT 191.480 102.480 192.155 102.640 ;
        RECT 192.615 102.560 193.835 102.730 ;
        RECT 191.480 101.690 191.690 102.480 ;
        RECT 192.615 102.470 192.785 102.560 ;
        RECT 191.860 101.690 192.210 102.310 ;
        RECT 192.380 102.300 192.785 102.470 ;
        RECT 192.380 101.520 192.550 102.300 ;
        RECT 192.720 101.850 192.940 102.130 ;
        RECT 193.120 102.020 193.660 102.390 ;
        RECT 194.005 102.310 194.175 102.900 ;
        RECT 194.395 102.480 194.700 103.620 ;
        RECT 194.870 102.430 195.125 103.310 ;
        RECT 194.005 102.280 194.745 102.310 ;
        RECT 192.720 101.680 193.250 101.850 ;
        RECT 191.030 101.260 191.380 101.430 ;
        RECT 191.600 101.240 192.550 101.520 ;
        RECT 192.720 101.070 192.910 101.510 ;
        RECT 193.080 101.450 193.250 101.680 ;
        RECT 193.420 101.620 193.660 102.020 ;
        RECT 193.830 101.980 194.745 102.280 ;
        RECT 193.830 101.805 194.155 101.980 ;
        RECT 193.830 101.450 194.150 101.805 ;
        RECT 194.915 101.780 195.125 102.430 ;
        RECT 193.080 101.280 194.150 101.450 ;
        RECT 194.395 101.070 194.700 101.530 ;
        RECT 194.870 101.250 195.125 101.780 ;
        RECT 195.305 102.480 195.640 103.450 ;
        RECT 195.810 102.480 195.980 103.620 ;
        RECT 196.150 103.280 198.180 103.450 ;
        RECT 195.305 101.810 195.475 102.480 ;
        RECT 196.150 102.310 196.320 103.280 ;
        RECT 195.645 101.980 195.900 102.310 ;
        RECT 196.125 101.980 196.320 102.310 ;
        RECT 196.490 102.940 197.615 103.110 ;
        RECT 195.730 101.810 195.900 101.980 ;
        RECT 196.490 101.810 196.660 102.940 ;
        RECT 195.305 101.240 195.560 101.810 ;
        RECT 195.730 101.640 196.660 101.810 ;
        RECT 196.830 102.600 197.840 102.770 ;
        RECT 196.830 101.800 197.000 102.600 ;
        RECT 197.205 102.260 197.480 102.400 ;
        RECT 197.200 102.090 197.480 102.260 ;
        RECT 196.485 101.605 196.660 101.640 ;
        RECT 195.730 101.070 196.060 101.470 ;
        RECT 196.485 101.240 197.015 101.605 ;
        RECT 197.205 101.240 197.480 102.090 ;
        RECT 197.650 101.240 197.840 102.600 ;
        RECT 198.010 102.615 198.180 103.280 ;
        RECT 198.350 102.860 198.520 103.620 ;
        RECT 198.755 102.860 199.270 103.270 ;
        RECT 198.010 102.425 198.760 102.615 ;
        RECT 198.930 102.050 199.270 102.860 ;
        RECT 199.440 102.530 200.650 103.620 ;
        RECT 198.040 101.880 199.270 102.050 ;
        RECT 198.020 101.070 198.530 101.605 ;
        RECT 198.750 101.275 198.995 101.880 ;
        RECT 199.440 101.820 199.960 102.360 ;
        RECT 200.130 101.990 200.650 102.530 ;
        RECT 200.820 102.455 201.110 103.620 ;
        RECT 201.370 102.690 201.540 103.450 ;
        RECT 201.755 102.860 202.085 103.620 ;
        RECT 201.370 102.520 202.085 102.690 ;
        RECT 202.255 102.545 202.510 103.450 ;
        RECT 201.280 101.970 201.635 102.340 ;
        RECT 201.915 102.310 202.085 102.520 ;
        RECT 201.915 101.980 202.170 102.310 ;
        RECT 199.440 101.070 200.650 101.820 ;
        RECT 200.820 101.070 201.110 101.795 ;
        RECT 201.915 101.790 202.085 101.980 ;
        RECT 202.340 101.815 202.510 102.545 ;
        RECT 202.685 102.470 202.945 103.620 ;
        RECT 203.125 102.950 203.380 103.450 ;
        RECT 203.550 103.120 203.880 103.620 ;
        RECT 203.125 102.780 203.875 102.950 ;
        RECT 203.125 101.960 203.475 102.610 ;
        RECT 201.370 101.620 202.085 101.790 ;
        RECT 201.370 101.240 201.540 101.620 ;
        RECT 201.755 101.070 202.085 101.450 ;
        RECT 202.255 101.240 202.510 101.815 ;
        RECT 202.685 101.070 202.945 101.910 ;
        RECT 203.645 101.790 203.875 102.780 ;
        RECT 203.125 101.620 203.875 101.790 ;
        RECT 203.125 101.330 203.380 101.620 ;
        RECT 203.550 101.070 203.880 101.450 ;
        RECT 204.050 101.330 204.220 103.450 ;
        RECT 204.390 102.650 204.715 103.435 ;
        RECT 204.885 103.160 205.135 103.620 ;
        RECT 205.305 103.120 205.555 103.450 ;
        RECT 205.770 103.120 206.450 103.450 ;
        RECT 205.305 102.990 205.475 103.120 ;
        RECT 205.080 102.820 205.475 102.990 ;
        RECT 204.450 101.600 204.910 102.650 ;
        RECT 205.080 101.460 205.250 102.820 ;
        RECT 205.645 102.560 206.110 102.950 ;
        RECT 205.420 101.750 205.770 102.370 ;
        RECT 205.940 101.970 206.110 102.560 ;
        RECT 206.280 102.340 206.450 103.120 ;
        RECT 206.620 103.020 206.790 103.360 ;
        RECT 207.025 103.190 207.355 103.620 ;
        RECT 207.525 103.020 207.695 103.360 ;
        RECT 207.990 103.160 208.360 103.620 ;
        RECT 206.620 102.850 207.695 103.020 ;
        RECT 208.530 102.990 208.700 103.450 ;
        RECT 208.935 103.110 209.805 103.450 ;
        RECT 209.975 103.160 210.225 103.620 ;
        RECT 208.140 102.820 208.700 102.990 ;
        RECT 208.140 102.680 208.310 102.820 ;
        RECT 206.810 102.510 208.310 102.680 ;
        RECT 209.005 102.650 209.465 102.940 ;
        RECT 206.280 102.170 207.970 102.340 ;
        RECT 205.940 101.750 206.295 101.970 ;
        RECT 206.465 101.460 206.635 102.170 ;
        RECT 206.840 101.750 207.630 102.000 ;
        RECT 207.800 101.990 207.970 102.170 ;
        RECT 208.140 101.820 208.310 102.510 ;
        RECT 204.580 101.070 204.910 101.430 ;
        RECT 205.080 101.290 205.575 101.460 ;
        RECT 205.780 101.290 206.635 101.460 ;
        RECT 207.510 101.070 207.840 101.530 ;
        RECT 208.050 101.430 208.310 101.820 ;
        RECT 208.500 102.640 209.465 102.650 ;
        RECT 209.635 102.730 209.805 103.110 ;
        RECT 210.395 103.070 210.565 103.360 ;
        RECT 210.745 103.240 211.075 103.620 ;
        RECT 210.395 102.900 211.195 103.070 ;
        RECT 208.500 102.480 209.175 102.640 ;
        RECT 209.635 102.560 210.855 102.730 ;
        RECT 208.500 101.690 208.710 102.480 ;
        RECT 209.635 102.470 209.805 102.560 ;
        RECT 208.880 101.690 209.230 102.310 ;
        RECT 209.400 102.300 209.805 102.470 ;
        RECT 209.400 101.520 209.570 102.300 ;
        RECT 209.740 101.850 209.960 102.130 ;
        RECT 210.140 102.020 210.680 102.390 ;
        RECT 211.025 102.310 211.195 102.900 ;
        RECT 211.415 102.480 211.720 103.620 ;
        RECT 211.890 102.430 212.145 103.310 ;
        RECT 211.025 102.280 211.765 102.310 ;
        RECT 209.740 101.680 210.270 101.850 ;
        RECT 208.050 101.260 208.400 101.430 ;
        RECT 208.620 101.240 209.570 101.520 ;
        RECT 209.740 101.070 209.930 101.510 ;
        RECT 210.100 101.450 210.270 101.680 ;
        RECT 210.440 101.620 210.680 102.020 ;
        RECT 210.850 101.980 211.765 102.280 ;
        RECT 210.850 101.805 211.175 101.980 ;
        RECT 210.850 101.450 211.170 101.805 ;
        RECT 211.935 101.780 212.145 102.430 ;
        RECT 210.100 101.280 211.170 101.450 ;
        RECT 211.415 101.070 211.720 101.530 ;
        RECT 211.890 101.250 212.145 101.780 ;
        RECT 212.325 102.480 212.660 103.450 ;
        RECT 212.830 102.480 213.000 103.620 ;
        RECT 213.170 103.280 215.200 103.450 ;
        RECT 212.325 101.810 212.495 102.480 ;
        RECT 213.170 102.310 213.340 103.280 ;
        RECT 212.665 101.980 212.920 102.310 ;
        RECT 213.145 101.980 213.340 102.310 ;
        RECT 213.510 102.940 214.635 103.110 ;
        RECT 212.750 101.810 212.920 101.980 ;
        RECT 213.510 101.810 213.680 102.940 ;
        RECT 212.325 101.240 212.580 101.810 ;
        RECT 212.750 101.640 213.680 101.810 ;
        RECT 213.850 102.600 214.860 102.770 ;
        RECT 213.850 101.800 214.020 102.600 ;
        RECT 213.505 101.605 213.680 101.640 ;
        RECT 212.750 101.070 213.080 101.470 ;
        RECT 213.505 101.240 214.035 101.605 ;
        RECT 214.225 101.580 214.500 102.400 ;
        RECT 214.220 101.410 214.500 101.580 ;
        RECT 214.225 101.240 214.500 101.410 ;
        RECT 214.670 101.240 214.860 102.600 ;
        RECT 215.030 102.615 215.200 103.280 ;
        RECT 215.370 102.860 215.540 103.620 ;
        RECT 215.775 102.860 216.290 103.270 ;
        RECT 215.030 102.425 215.780 102.615 ;
        RECT 215.950 102.050 216.290 102.860 ;
        RECT 217.385 102.950 217.640 103.450 ;
        RECT 217.810 103.120 218.140 103.620 ;
        RECT 217.385 102.780 218.135 102.950 ;
        RECT 215.060 101.880 216.290 102.050 ;
        RECT 217.385 101.960 217.735 102.610 ;
        RECT 215.040 101.070 215.550 101.605 ;
        RECT 215.770 101.275 216.015 101.880 ;
        RECT 217.905 101.790 218.135 102.780 ;
        RECT 217.385 101.620 218.135 101.790 ;
        RECT 217.385 101.330 217.640 101.620 ;
        RECT 217.810 101.070 218.140 101.450 ;
        RECT 218.310 101.330 218.480 103.450 ;
        RECT 218.650 102.650 218.975 103.435 ;
        RECT 219.145 103.160 219.395 103.620 ;
        RECT 219.565 103.120 219.815 103.450 ;
        RECT 220.030 103.120 220.710 103.450 ;
        RECT 219.565 102.990 219.735 103.120 ;
        RECT 219.340 102.820 219.735 102.990 ;
        RECT 218.710 101.600 219.170 102.650 ;
        RECT 219.340 101.460 219.510 102.820 ;
        RECT 219.905 102.560 220.370 102.950 ;
        RECT 219.680 101.750 220.030 102.370 ;
        RECT 220.200 101.970 220.370 102.560 ;
        RECT 220.540 102.340 220.710 103.120 ;
        RECT 220.880 103.020 221.050 103.360 ;
        RECT 221.285 103.190 221.615 103.620 ;
        RECT 221.785 103.020 221.955 103.360 ;
        RECT 222.250 103.160 222.620 103.620 ;
        RECT 220.880 102.850 221.955 103.020 ;
        RECT 222.790 102.990 222.960 103.450 ;
        RECT 223.195 103.110 224.065 103.450 ;
        RECT 224.235 103.160 224.485 103.620 ;
        RECT 222.400 102.820 222.960 102.990 ;
        RECT 222.400 102.680 222.570 102.820 ;
        RECT 221.070 102.510 222.570 102.680 ;
        RECT 223.265 102.650 223.725 102.940 ;
        RECT 220.540 102.170 222.230 102.340 ;
        RECT 220.200 101.750 220.555 101.970 ;
        RECT 220.725 101.460 220.895 102.170 ;
        RECT 221.100 101.750 221.890 102.000 ;
        RECT 222.060 101.990 222.230 102.170 ;
        RECT 222.400 101.820 222.570 102.510 ;
        RECT 218.840 101.070 219.170 101.430 ;
        RECT 219.340 101.290 219.835 101.460 ;
        RECT 220.040 101.290 220.895 101.460 ;
        RECT 221.770 101.070 222.100 101.530 ;
        RECT 222.310 101.430 222.570 101.820 ;
        RECT 222.760 102.640 223.725 102.650 ;
        RECT 223.895 102.730 224.065 103.110 ;
        RECT 224.655 103.070 224.825 103.360 ;
        RECT 225.005 103.240 225.335 103.620 ;
        RECT 224.655 102.900 225.455 103.070 ;
        RECT 222.760 102.480 223.435 102.640 ;
        RECT 223.895 102.560 225.115 102.730 ;
        RECT 222.760 101.690 222.970 102.480 ;
        RECT 223.895 102.470 224.065 102.560 ;
        RECT 223.140 101.690 223.490 102.310 ;
        RECT 223.660 102.300 224.065 102.470 ;
        RECT 223.660 101.520 223.830 102.300 ;
        RECT 224.000 101.850 224.220 102.130 ;
        RECT 224.400 102.020 224.940 102.390 ;
        RECT 225.285 102.310 225.455 102.900 ;
        RECT 225.675 102.480 225.980 103.620 ;
        RECT 226.150 102.430 226.405 103.310 ;
        RECT 226.580 102.455 226.870 103.620 ;
        RECT 227.045 102.480 227.380 103.450 ;
        RECT 227.550 102.480 227.720 103.620 ;
        RECT 227.890 103.280 229.920 103.450 ;
        RECT 225.285 102.280 226.025 102.310 ;
        RECT 224.000 101.680 224.530 101.850 ;
        RECT 222.310 101.260 222.660 101.430 ;
        RECT 222.880 101.240 223.830 101.520 ;
        RECT 224.000 101.070 224.190 101.510 ;
        RECT 224.360 101.450 224.530 101.680 ;
        RECT 224.700 101.620 224.940 102.020 ;
        RECT 225.110 101.980 226.025 102.280 ;
        RECT 225.110 101.805 225.435 101.980 ;
        RECT 225.110 101.450 225.430 101.805 ;
        RECT 226.195 101.780 226.405 102.430 ;
        RECT 227.045 101.810 227.215 102.480 ;
        RECT 227.890 102.310 228.060 103.280 ;
        RECT 227.385 101.980 227.640 102.310 ;
        RECT 227.865 101.980 228.060 102.310 ;
        RECT 228.230 102.940 229.355 103.110 ;
        RECT 227.470 101.810 227.640 101.980 ;
        RECT 228.230 101.810 228.400 102.940 ;
        RECT 224.360 101.280 225.430 101.450 ;
        RECT 225.675 101.070 225.980 101.530 ;
        RECT 226.150 101.250 226.405 101.780 ;
        RECT 226.580 101.070 226.870 101.795 ;
        RECT 227.045 101.240 227.300 101.810 ;
        RECT 227.470 101.640 228.400 101.810 ;
        RECT 228.570 102.600 229.580 102.770 ;
        RECT 228.570 101.800 228.740 102.600 ;
        RECT 228.225 101.605 228.400 101.640 ;
        RECT 227.470 101.070 227.800 101.470 ;
        RECT 228.225 101.240 228.755 101.605 ;
        RECT 228.945 101.580 229.220 102.400 ;
        RECT 228.940 101.410 229.220 101.580 ;
        RECT 228.945 101.240 229.220 101.410 ;
        RECT 229.390 101.240 229.580 102.600 ;
        RECT 229.750 102.615 229.920 103.280 ;
        RECT 230.090 102.860 230.260 103.620 ;
        RECT 230.495 102.860 231.010 103.270 ;
        RECT 229.750 102.425 230.500 102.615 ;
        RECT 230.670 102.050 231.010 102.860 ;
        RECT 231.185 102.470 231.445 103.620 ;
        RECT 231.620 102.545 231.875 103.450 ;
        RECT 232.045 102.860 232.375 103.620 ;
        RECT 232.590 102.690 232.760 103.450 ;
        RECT 229.780 101.880 231.010 102.050 ;
        RECT 229.760 101.070 230.270 101.605 ;
        RECT 230.490 101.275 230.735 101.880 ;
        RECT 231.185 101.070 231.445 101.910 ;
        RECT 231.620 101.815 231.790 102.545 ;
        RECT 232.045 102.520 232.760 102.690 ;
        RECT 233.020 102.530 236.530 103.620 ;
        RECT 236.705 102.950 236.960 103.450 ;
        RECT 237.130 103.120 237.460 103.620 ;
        RECT 236.705 102.780 237.455 102.950 ;
        RECT 232.045 102.310 232.215 102.520 ;
        RECT 231.960 101.980 232.215 102.310 ;
        RECT 231.620 101.240 231.875 101.815 ;
        RECT 232.045 101.790 232.215 101.980 ;
        RECT 232.495 101.970 232.850 102.340 ;
        RECT 233.020 101.840 234.670 102.360 ;
        RECT 234.840 102.010 236.530 102.530 ;
        RECT 236.705 101.960 237.055 102.610 ;
        RECT 232.045 101.620 232.760 101.790 ;
        RECT 232.045 101.070 232.375 101.450 ;
        RECT 232.590 101.240 232.760 101.620 ;
        RECT 233.020 101.070 236.530 101.840 ;
        RECT 237.225 101.790 237.455 102.780 ;
        RECT 236.705 101.620 237.455 101.790 ;
        RECT 236.705 101.330 236.960 101.620 ;
        RECT 237.130 101.070 237.460 101.450 ;
        RECT 237.630 101.330 237.800 103.450 ;
        RECT 237.970 102.650 238.295 103.435 ;
        RECT 238.465 103.160 238.715 103.620 ;
        RECT 238.885 103.120 239.135 103.450 ;
        RECT 239.350 103.120 240.030 103.450 ;
        RECT 238.885 102.990 239.055 103.120 ;
        RECT 238.660 102.820 239.055 102.990 ;
        RECT 238.030 101.600 238.490 102.650 ;
        RECT 238.660 101.460 238.830 102.820 ;
        RECT 239.225 102.560 239.690 102.950 ;
        RECT 239.000 101.750 239.350 102.370 ;
        RECT 239.520 101.970 239.690 102.560 ;
        RECT 239.860 102.340 240.030 103.120 ;
        RECT 240.200 103.020 240.370 103.360 ;
        RECT 240.605 103.190 240.935 103.620 ;
        RECT 241.105 103.020 241.275 103.360 ;
        RECT 241.570 103.160 241.940 103.620 ;
        RECT 240.200 102.850 241.275 103.020 ;
        RECT 242.110 102.990 242.280 103.450 ;
        RECT 242.515 103.110 243.385 103.450 ;
        RECT 243.555 103.160 243.805 103.620 ;
        RECT 241.720 102.820 242.280 102.990 ;
        RECT 241.720 102.680 241.890 102.820 ;
        RECT 240.390 102.510 241.890 102.680 ;
        RECT 242.585 102.650 243.045 102.940 ;
        RECT 239.860 102.170 241.550 102.340 ;
        RECT 239.520 101.750 239.875 101.970 ;
        RECT 240.045 101.460 240.215 102.170 ;
        RECT 240.420 101.750 241.210 102.000 ;
        RECT 241.380 101.990 241.550 102.170 ;
        RECT 241.720 101.820 241.890 102.510 ;
        RECT 238.160 101.070 238.490 101.430 ;
        RECT 238.660 101.290 239.155 101.460 ;
        RECT 239.360 101.290 240.215 101.460 ;
        RECT 241.090 101.070 241.420 101.530 ;
        RECT 241.630 101.430 241.890 101.820 ;
        RECT 242.080 102.640 243.045 102.650 ;
        RECT 243.215 102.730 243.385 103.110 ;
        RECT 243.975 103.070 244.145 103.360 ;
        RECT 244.325 103.240 244.655 103.620 ;
        RECT 243.975 102.900 244.775 103.070 ;
        RECT 242.080 102.480 242.755 102.640 ;
        RECT 243.215 102.560 244.435 102.730 ;
        RECT 242.080 101.690 242.290 102.480 ;
        RECT 243.215 102.470 243.385 102.560 ;
        RECT 242.460 101.690 242.810 102.310 ;
        RECT 242.980 102.300 243.385 102.470 ;
        RECT 242.980 101.520 243.150 102.300 ;
        RECT 243.320 101.850 243.540 102.130 ;
        RECT 243.720 102.020 244.260 102.390 ;
        RECT 244.605 102.310 244.775 102.900 ;
        RECT 244.995 102.480 245.300 103.620 ;
        RECT 245.470 102.430 245.725 103.310 ;
        RECT 244.605 102.280 245.345 102.310 ;
        RECT 243.320 101.680 243.850 101.850 ;
        RECT 241.630 101.260 241.980 101.430 ;
        RECT 242.200 101.240 243.150 101.520 ;
        RECT 243.320 101.070 243.510 101.510 ;
        RECT 243.680 101.450 243.850 101.680 ;
        RECT 244.020 101.620 244.260 102.020 ;
        RECT 244.430 101.980 245.345 102.280 ;
        RECT 244.430 101.805 244.755 101.980 ;
        RECT 244.430 101.450 244.750 101.805 ;
        RECT 245.515 101.780 245.725 102.430 ;
        RECT 243.680 101.280 244.750 101.450 ;
        RECT 244.995 101.070 245.300 101.530 ;
        RECT 245.470 101.250 245.725 101.780 ;
        RECT 245.905 102.480 246.240 103.450 ;
        RECT 246.410 102.480 246.580 103.620 ;
        RECT 246.750 103.280 248.780 103.450 ;
        RECT 245.905 101.810 246.075 102.480 ;
        RECT 246.750 102.310 246.920 103.280 ;
        RECT 246.245 101.980 246.500 102.310 ;
        RECT 246.725 101.980 246.920 102.310 ;
        RECT 247.090 102.940 248.215 103.110 ;
        RECT 246.330 101.810 246.500 101.980 ;
        RECT 247.090 101.810 247.260 102.940 ;
        RECT 245.905 101.240 246.160 101.810 ;
        RECT 246.330 101.640 247.260 101.810 ;
        RECT 247.430 102.600 248.440 102.770 ;
        RECT 247.430 101.800 247.600 102.600 ;
        RECT 247.085 101.605 247.260 101.640 ;
        RECT 246.330 101.070 246.660 101.470 ;
        RECT 247.085 101.240 247.615 101.605 ;
        RECT 247.805 101.580 248.080 102.400 ;
        RECT 247.800 101.410 248.080 101.580 ;
        RECT 247.805 101.240 248.080 101.410 ;
        RECT 248.250 101.240 248.440 102.600 ;
        RECT 248.610 102.615 248.780 103.280 ;
        RECT 248.950 102.860 249.120 103.620 ;
        RECT 249.355 102.860 249.870 103.270 ;
        RECT 248.610 102.425 249.360 102.615 ;
        RECT 249.530 102.050 249.870 102.860 ;
        RECT 250.045 102.470 250.305 103.620 ;
        RECT 250.480 102.545 250.735 103.450 ;
        RECT 250.905 102.860 251.235 103.620 ;
        RECT 251.450 102.690 251.620 103.450 ;
        RECT 248.640 101.880 249.870 102.050 ;
        RECT 248.620 101.070 249.130 101.605 ;
        RECT 249.350 101.275 249.595 101.880 ;
        RECT 250.045 101.070 250.305 101.910 ;
        RECT 250.480 101.815 250.650 102.545 ;
        RECT 250.905 102.520 251.620 102.690 ;
        RECT 250.905 102.310 251.075 102.520 ;
        RECT 252.340 102.455 252.630 103.620 ;
        RECT 252.805 102.950 253.060 103.450 ;
        RECT 253.230 103.120 253.560 103.620 ;
        RECT 252.805 102.780 253.555 102.950 ;
        RECT 250.820 101.980 251.075 102.310 ;
        RECT 250.480 101.240 250.735 101.815 ;
        RECT 250.905 101.790 251.075 101.980 ;
        RECT 251.355 101.970 251.710 102.340 ;
        RECT 252.805 101.960 253.155 102.610 ;
        RECT 250.905 101.620 251.620 101.790 ;
        RECT 250.905 101.070 251.235 101.450 ;
        RECT 251.450 101.240 251.620 101.620 ;
        RECT 252.340 101.070 252.630 101.795 ;
        RECT 253.325 101.790 253.555 102.780 ;
        RECT 252.805 101.620 253.555 101.790 ;
        RECT 252.805 101.330 253.060 101.620 ;
        RECT 253.230 101.070 253.560 101.450 ;
        RECT 253.730 101.330 253.900 103.450 ;
        RECT 254.070 102.650 254.395 103.435 ;
        RECT 254.565 103.160 254.815 103.620 ;
        RECT 254.985 103.120 255.235 103.450 ;
        RECT 255.450 103.120 256.130 103.450 ;
        RECT 254.985 102.990 255.155 103.120 ;
        RECT 254.760 102.820 255.155 102.990 ;
        RECT 254.130 101.600 254.590 102.650 ;
        RECT 254.760 101.460 254.930 102.820 ;
        RECT 255.325 102.560 255.790 102.950 ;
        RECT 255.100 101.750 255.450 102.370 ;
        RECT 255.620 101.970 255.790 102.560 ;
        RECT 255.960 102.340 256.130 103.120 ;
        RECT 256.300 103.020 256.470 103.360 ;
        RECT 256.705 103.190 257.035 103.620 ;
        RECT 257.205 103.020 257.375 103.360 ;
        RECT 257.670 103.160 258.040 103.620 ;
        RECT 256.300 102.850 257.375 103.020 ;
        RECT 258.210 102.990 258.380 103.450 ;
        RECT 258.615 103.110 259.485 103.450 ;
        RECT 259.655 103.160 259.905 103.620 ;
        RECT 257.820 102.820 258.380 102.990 ;
        RECT 257.820 102.680 257.990 102.820 ;
        RECT 256.490 102.510 257.990 102.680 ;
        RECT 258.685 102.650 259.145 102.940 ;
        RECT 255.960 102.170 257.650 102.340 ;
        RECT 255.620 101.750 255.975 101.970 ;
        RECT 256.145 101.460 256.315 102.170 ;
        RECT 256.520 101.750 257.310 102.000 ;
        RECT 257.480 101.990 257.650 102.170 ;
        RECT 257.820 101.820 257.990 102.510 ;
        RECT 254.260 101.070 254.590 101.430 ;
        RECT 254.760 101.290 255.255 101.460 ;
        RECT 255.460 101.290 256.315 101.460 ;
        RECT 257.190 101.070 257.520 101.530 ;
        RECT 257.730 101.430 257.990 101.820 ;
        RECT 258.180 102.640 259.145 102.650 ;
        RECT 259.315 102.730 259.485 103.110 ;
        RECT 260.075 103.070 260.245 103.360 ;
        RECT 260.425 103.240 260.755 103.620 ;
        RECT 260.075 102.900 260.875 103.070 ;
        RECT 258.180 102.480 258.855 102.640 ;
        RECT 259.315 102.560 260.535 102.730 ;
        RECT 258.180 101.690 258.390 102.480 ;
        RECT 259.315 102.470 259.485 102.560 ;
        RECT 258.560 101.690 258.910 102.310 ;
        RECT 259.080 102.300 259.485 102.470 ;
        RECT 259.080 101.520 259.250 102.300 ;
        RECT 259.420 101.850 259.640 102.130 ;
        RECT 259.820 102.020 260.360 102.390 ;
        RECT 260.705 102.310 260.875 102.900 ;
        RECT 261.095 102.480 261.400 103.620 ;
        RECT 261.570 102.430 261.825 103.310 ;
        RECT 262.005 102.950 262.260 103.450 ;
        RECT 262.430 103.120 262.760 103.620 ;
        RECT 262.005 102.780 262.755 102.950 ;
        RECT 260.705 102.280 261.445 102.310 ;
        RECT 259.420 101.680 259.950 101.850 ;
        RECT 257.730 101.260 258.080 101.430 ;
        RECT 258.300 101.240 259.250 101.520 ;
        RECT 259.420 101.070 259.610 101.510 ;
        RECT 259.780 101.450 259.950 101.680 ;
        RECT 260.120 101.620 260.360 102.020 ;
        RECT 260.530 101.980 261.445 102.280 ;
        RECT 260.530 101.805 260.855 101.980 ;
        RECT 260.530 101.450 260.850 101.805 ;
        RECT 261.615 101.780 261.825 102.430 ;
        RECT 262.005 101.960 262.355 102.610 ;
        RECT 262.525 101.790 262.755 102.780 ;
        RECT 259.780 101.280 260.850 101.450 ;
        RECT 261.095 101.070 261.400 101.530 ;
        RECT 261.570 101.250 261.825 101.780 ;
        RECT 262.005 101.620 262.755 101.790 ;
        RECT 262.005 101.330 262.260 101.620 ;
        RECT 262.430 101.070 262.760 101.450 ;
        RECT 262.930 101.330 263.100 103.450 ;
        RECT 263.270 102.650 263.595 103.435 ;
        RECT 263.765 103.160 264.015 103.620 ;
        RECT 264.185 103.120 264.435 103.450 ;
        RECT 264.650 103.120 265.330 103.450 ;
        RECT 264.185 102.990 264.355 103.120 ;
        RECT 263.960 102.820 264.355 102.990 ;
        RECT 263.330 101.600 263.790 102.650 ;
        RECT 263.960 101.460 264.130 102.820 ;
        RECT 264.525 102.560 264.990 102.950 ;
        RECT 264.300 101.750 264.650 102.370 ;
        RECT 264.820 101.970 264.990 102.560 ;
        RECT 265.160 102.340 265.330 103.120 ;
        RECT 265.500 103.020 265.670 103.360 ;
        RECT 265.905 103.190 266.235 103.620 ;
        RECT 266.405 103.020 266.575 103.360 ;
        RECT 266.870 103.160 267.240 103.620 ;
        RECT 265.500 102.850 266.575 103.020 ;
        RECT 267.410 102.990 267.580 103.450 ;
        RECT 267.815 103.110 268.685 103.450 ;
        RECT 268.855 103.160 269.105 103.620 ;
        RECT 267.020 102.820 267.580 102.990 ;
        RECT 267.020 102.680 267.190 102.820 ;
        RECT 265.690 102.510 267.190 102.680 ;
        RECT 267.885 102.650 268.345 102.940 ;
        RECT 265.160 102.170 266.850 102.340 ;
        RECT 264.820 101.750 265.175 101.970 ;
        RECT 265.345 101.460 265.515 102.170 ;
        RECT 265.720 101.750 266.510 102.000 ;
        RECT 266.680 101.990 266.850 102.170 ;
        RECT 267.020 101.820 267.190 102.510 ;
        RECT 263.460 101.070 263.790 101.430 ;
        RECT 263.960 101.290 264.455 101.460 ;
        RECT 264.660 101.290 265.515 101.460 ;
        RECT 266.390 101.070 266.720 101.530 ;
        RECT 266.930 101.430 267.190 101.820 ;
        RECT 267.380 102.640 268.345 102.650 ;
        RECT 268.515 102.730 268.685 103.110 ;
        RECT 269.275 103.070 269.445 103.360 ;
        RECT 269.625 103.240 269.955 103.620 ;
        RECT 269.275 102.900 270.075 103.070 ;
        RECT 267.380 102.480 268.055 102.640 ;
        RECT 268.515 102.560 269.735 102.730 ;
        RECT 267.380 101.690 267.590 102.480 ;
        RECT 268.515 102.470 268.685 102.560 ;
        RECT 267.760 101.690 268.110 102.310 ;
        RECT 268.280 102.300 268.685 102.470 ;
        RECT 268.280 101.520 268.450 102.300 ;
        RECT 268.620 101.850 268.840 102.130 ;
        RECT 269.020 102.020 269.560 102.390 ;
        RECT 269.905 102.310 270.075 102.900 ;
        RECT 270.295 102.480 270.600 103.620 ;
        RECT 270.770 102.430 271.025 103.310 ;
        RECT 269.905 102.280 270.645 102.310 ;
        RECT 268.620 101.680 269.150 101.850 ;
        RECT 266.930 101.260 267.280 101.430 ;
        RECT 267.500 101.240 268.450 101.520 ;
        RECT 268.620 101.070 268.810 101.510 ;
        RECT 268.980 101.450 269.150 101.680 ;
        RECT 269.320 101.620 269.560 102.020 ;
        RECT 269.730 101.980 270.645 102.280 ;
        RECT 269.730 101.805 270.055 101.980 ;
        RECT 269.730 101.450 270.050 101.805 ;
        RECT 270.815 101.780 271.025 102.430 ;
        RECT 271.200 102.860 271.715 103.270 ;
        RECT 271.950 102.860 272.120 103.620 ;
        RECT 272.290 103.280 274.320 103.450 ;
        RECT 271.200 102.050 271.540 102.860 ;
        RECT 272.290 102.615 272.460 103.280 ;
        RECT 272.855 102.940 273.980 103.110 ;
        RECT 271.710 102.425 272.460 102.615 ;
        RECT 272.630 102.600 273.640 102.770 ;
        RECT 271.200 101.880 272.430 102.050 ;
        RECT 268.980 101.280 270.050 101.450 ;
        RECT 270.295 101.070 270.600 101.530 ;
        RECT 270.770 101.250 271.025 101.780 ;
        RECT 271.475 101.275 271.720 101.880 ;
        RECT 271.940 101.070 272.450 101.605 ;
        RECT 272.630 101.240 272.820 102.600 ;
        RECT 272.990 102.260 273.265 102.400 ;
        RECT 272.990 102.090 273.270 102.260 ;
        RECT 272.990 101.240 273.265 102.090 ;
        RECT 273.470 101.800 273.640 102.600 ;
        RECT 273.810 101.810 273.980 102.940 ;
        RECT 274.150 102.310 274.320 103.280 ;
        RECT 274.490 102.480 274.660 103.620 ;
        RECT 274.830 102.480 275.165 103.450 ;
        RECT 274.150 101.980 274.345 102.310 ;
        RECT 274.570 101.980 274.825 102.310 ;
        RECT 274.570 101.810 274.740 101.980 ;
        RECT 274.995 101.810 275.165 102.480 ;
        RECT 275.345 102.470 275.605 103.620 ;
        RECT 275.780 102.545 276.035 103.450 ;
        RECT 276.205 102.860 276.535 103.620 ;
        RECT 276.750 102.690 276.920 103.450 ;
        RECT 273.810 101.640 274.740 101.810 ;
        RECT 273.810 101.605 273.985 101.640 ;
        RECT 273.455 101.240 273.985 101.605 ;
        RECT 274.410 101.070 274.740 101.470 ;
        RECT 274.910 101.240 275.165 101.810 ;
        RECT 275.345 101.070 275.605 101.910 ;
        RECT 275.780 101.815 275.950 102.545 ;
        RECT 276.205 102.520 276.920 102.690 ;
        RECT 276.205 102.310 276.375 102.520 ;
        RECT 278.100 102.455 278.390 103.620 ;
        RECT 278.565 102.430 278.820 103.310 ;
        RECT 278.990 102.480 279.295 103.620 ;
        RECT 279.635 103.240 279.965 103.620 ;
        RECT 280.145 103.070 280.315 103.360 ;
        RECT 280.485 103.160 280.735 103.620 ;
        RECT 279.515 102.900 280.315 103.070 ;
        RECT 280.905 103.110 281.775 103.450 ;
        RECT 276.120 101.980 276.375 102.310 ;
        RECT 275.780 101.240 276.035 101.815 ;
        RECT 276.205 101.790 276.375 101.980 ;
        RECT 276.655 101.970 277.010 102.340 ;
        RECT 276.205 101.620 276.920 101.790 ;
        RECT 276.205 101.070 276.535 101.450 ;
        RECT 276.750 101.240 276.920 101.620 ;
        RECT 278.100 101.070 278.390 101.795 ;
        RECT 278.565 101.780 278.775 102.430 ;
        RECT 279.515 102.310 279.685 102.900 ;
        RECT 280.905 102.730 281.075 103.110 ;
        RECT 282.010 102.990 282.180 103.450 ;
        RECT 282.350 103.160 282.720 103.620 ;
        RECT 283.015 103.020 283.185 103.360 ;
        RECT 283.355 103.190 283.685 103.620 ;
        RECT 283.920 103.020 284.090 103.360 ;
        RECT 279.855 102.560 281.075 102.730 ;
        RECT 281.245 102.650 281.705 102.940 ;
        RECT 282.010 102.820 282.570 102.990 ;
        RECT 283.015 102.850 284.090 103.020 ;
        RECT 284.260 103.120 284.940 103.450 ;
        RECT 285.155 103.120 285.405 103.450 ;
        RECT 285.575 103.160 285.825 103.620 ;
        RECT 282.400 102.680 282.570 102.820 ;
        RECT 281.245 102.640 282.210 102.650 ;
        RECT 280.905 102.470 281.075 102.560 ;
        RECT 281.535 102.480 282.210 102.640 ;
        RECT 278.945 102.280 279.685 102.310 ;
        RECT 278.945 101.980 279.860 102.280 ;
        RECT 279.535 101.805 279.860 101.980 ;
        RECT 278.565 101.250 278.820 101.780 ;
        RECT 278.990 101.070 279.295 101.530 ;
        RECT 279.540 101.450 279.860 101.805 ;
        RECT 280.030 102.020 280.570 102.390 ;
        RECT 280.905 102.300 281.310 102.470 ;
        RECT 280.030 101.620 280.270 102.020 ;
        RECT 280.750 101.850 280.970 102.130 ;
        RECT 280.440 101.680 280.970 101.850 ;
        RECT 280.440 101.450 280.610 101.680 ;
        RECT 281.140 101.520 281.310 102.300 ;
        RECT 281.480 101.690 281.830 102.310 ;
        RECT 282.000 101.690 282.210 102.480 ;
        RECT 282.400 102.510 283.900 102.680 ;
        RECT 282.400 101.820 282.570 102.510 ;
        RECT 284.260 102.340 284.430 103.120 ;
        RECT 285.235 102.990 285.405 103.120 ;
        RECT 282.740 102.170 284.430 102.340 ;
        RECT 284.600 102.560 285.065 102.950 ;
        RECT 285.235 102.820 285.630 102.990 ;
        RECT 282.740 101.990 282.910 102.170 ;
        RECT 279.540 101.280 280.610 101.450 ;
        RECT 280.780 101.070 280.970 101.510 ;
        RECT 281.140 101.240 282.090 101.520 ;
        RECT 282.400 101.430 282.660 101.820 ;
        RECT 283.080 101.750 283.870 102.000 ;
        RECT 282.310 101.260 282.660 101.430 ;
        RECT 282.870 101.070 283.200 101.530 ;
        RECT 284.075 101.460 284.245 102.170 ;
        RECT 284.600 101.970 284.770 102.560 ;
        RECT 284.415 101.750 284.770 101.970 ;
        RECT 284.940 101.750 285.290 102.370 ;
        RECT 285.460 101.460 285.630 102.820 ;
        RECT 285.995 102.650 286.320 103.435 ;
        RECT 285.800 101.600 286.260 102.650 ;
        RECT 284.075 101.290 284.930 101.460 ;
        RECT 285.135 101.290 285.630 101.460 ;
        RECT 285.800 101.070 286.130 101.430 ;
        RECT 286.490 101.330 286.660 103.450 ;
        RECT 286.830 103.120 287.160 103.620 ;
        RECT 287.330 102.950 287.585 103.450 ;
        RECT 286.835 102.780 287.585 102.950 ;
        RECT 288.685 102.950 288.940 103.450 ;
        RECT 289.110 103.120 289.440 103.620 ;
        RECT 288.685 102.780 289.435 102.950 ;
        RECT 286.835 101.790 287.065 102.780 ;
        RECT 287.235 101.960 287.585 102.610 ;
        RECT 288.685 101.960 289.035 102.610 ;
        RECT 289.205 101.790 289.435 102.780 ;
        RECT 286.835 101.620 287.585 101.790 ;
        RECT 286.830 101.070 287.160 101.450 ;
        RECT 287.330 101.330 287.585 101.620 ;
        RECT 288.685 101.620 289.435 101.790 ;
        RECT 288.685 101.330 288.940 101.620 ;
        RECT 289.110 101.070 289.440 101.450 ;
        RECT 289.610 101.330 289.780 103.450 ;
        RECT 289.950 102.650 290.275 103.435 ;
        RECT 290.445 103.160 290.695 103.620 ;
        RECT 290.865 103.120 291.115 103.450 ;
        RECT 291.330 103.120 292.010 103.450 ;
        RECT 290.865 102.990 291.035 103.120 ;
        RECT 290.640 102.820 291.035 102.990 ;
        RECT 290.010 101.600 290.470 102.650 ;
        RECT 290.640 101.460 290.810 102.820 ;
        RECT 291.205 102.560 291.670 102.950 ;
        RECT 290.980 101.750 291.330 102.370 ;
        RECT 291.500 101.970 291.670 102.560 ;
        RECT 291.840 102.340 292.010 103.120 ;
        RECT 292.180 103.020 292.350 103.360 ;
        RECT 292.585 103.190 292.915 103.620 ;
        RECT 293.085 103.020 293.255 103.360 ;
        RECT 293.550 103.160 293.920 103.620 ;
        RECT 292.180 102.850 293.255 103.020 ;
        RECT 294.090 102.990 294.260 103.450 ;
        RECT 294.495 103.110 295.365 103.450 ;
        RECT 295.535 103.160 295.785 103.620 ;
        RECT 293.700 102.820 294.260 102.990 ;
        RECT 293.700 102.680 293.870 102.820 ;
        RECT 292.370 102.510 293.870 102.680 ;
        RECT 294.565 102.650 295.025 102.940 ;
        RECT 291.840 102.170 293.530 102.340 ;
        RECT 291.500 101.750 291.855 101.970 ;
        RECT 292.025 101.460 292.195 102.170 ;
        RECT 292.400 101.750 293.190 102.000 ;
        RECT 293.360 101.990 293.530 102.170 ;
        RECT 293.700 101.820 293.870 102.510 ;
        RECT 290.140 101.070 290.470 101.430 ;
        RECT 290.640 101.290 291.135 101.460 ;
        RECT 291.340 101.290 292.195 101.460 ;
        RECT 293.070 101.070 293.400 101.530 ;
        RECT 293.610 101.430 293.870 101.820 ;
        RECT 294.060 102.640 295.025 102.650 ;
        RECT 295.195 102.730 295.365 103.110 ;
        RECT 295.955 103.070 296.125 103.360 ;
        RECT 296.305 103.240 296.635 103.620 ;
        RECT 295.955 102.900 296.755 103.070 ;
        RECT 294.060 102.480 294.735 102.640 ;
        RECT 295.195 102.560 296.415 102.730 ;
        RECT 294.060 101.690 294.270 102.480 ;
        RECT 295.195 102.470 295.365 102.560 ;
        RECT 294.440 101.690 294.790 102.310 ;
        RECT 294.960 102.300 295.365 102.470 ;
        RECT 294.960 101.520 295.130 102.300 ;
        RECT 295.300 101.850 295.520 102.130 ;
        RECT 295.700 102.020 296.240 102.390 ;
        RECT 296.585 102.310 296.755 102.900 ;
        RECT 296.975 102.480 297.280 103.620 ;
        RECT 297.450 102.430 297.705 103.310 ;
        RECT 296.585 102.280 297.325 102.310 ;
        RECT 295.300 101.680 295.830 101.850 ;
        RECT 293.610 101.260 293.960 101.430 ;
        RECT 294.180 101.240 295.130 101.520 ;
        RECT 295.300 101.070 295.490 101.510 ;
        RECT 295.660 101.450 295.830 101.680 ;
        RECT 296.000 101.620 296.240 102.020 ;
        RECT 296.410 101.980 297.325 102.280 ;
        RECT 296.410 101.805 296.735 101.980 ;
        RECT 296.410 101.450 296.730 101.805 ;
        RECT 297.495 101.780 297.705 102.430 ;
        RECT 295.660 101.280 296.730 101.450 ;
        RECT 296.975 101.070 297.280 101.530 ;
        RECT 297.450 101.250 297.705 101.780 ;
        RECT 297.885 102.480 298.220 103.450 ;
        RECT 298.390 102.480 298.560 103.620 ;
        RECT 298.730 103.280 300.760 103.450 ;
        RECT 297.885 101.810 298.055 102.480 ;
        RECT 298.730 102.310 298.900 103.280 ;
        RECT 298.225 101.980 298.480 102.310 ;
        RECT 298.705 101.980 298.900 102.310 ;
        RECT 299.070 102.940 300.195 103.110 ;
        RECT 298.310 101.810 298.480 101.980 ;
        RECT 299.070 101.810 299.240 102.940 ;
        RECT 297.885 101.240 298.140 101.810 ;
        RECT 298.310 101.640 299.240 101.810 ;
        RECT 299.410 102.600 300.420 102.770 ;
        RECT 299.410 101.800 299.580 102.600 ;
        RECT 299.785 101.920 300.060 102.400 ;
        RECT 299.780 101.750 300.060 101.920 ;
        RECT 299.065 101.605 299.240 101.640 ;
        RECT 298.310 101.070 298.640 101.470 ;
        RECT 299.065 101.240 299.595 101.605 ;
        RECT 299.785 101.240 300.060 101.750 ;
        RECT 300.230 101.240 300.420 102.600 ;
        RECT 300.590 102.615 300.760 103.280 ;
        RECT 300.930 102.860 301.100 103.620 ;
        RECT 301.335 102.860 301.850 103.270 ;
        RECT 300.590 102.425 301.340 102.615 ;
        RECT 301.510 102.050 301.850 102.860 ;
        RECT 302.110 102.690 302.280 103.450 ;
        RECT 302.495 102.860 302.825 103.620 ;
        RECT 302.110 102.520 302.825 102.690 ;
        RECT 302.995 102.545 303.250 103.450 ;
        RECT 300.620 101.880 301.850 102.050 ;
        RECT 302.020 101.970 302.375 102.340 ;
        RECT 302.655 102.310 302.825 102.520 ;
        RECT 302.655 101.980 302.910 102.310 ;
        RECT 300.600 101.070 301.110 101.605 ;
        RECT 301.330 101.275 301.575 101.880 ;
        RECT 302.655 101.790 302.825 101.980 ;
        RECT 303.080 101.815 303.250 102.545 ;
        RECT 303.425 102.470 303.685 103.620 ;
        RECT 303.860 102.455 304.150 103.620 ;
        RECT 304.325 102.480 304.660 103.450 ;
        RECT 304.830 102.480 305.000 103.620 ;
        RECT 305.170 103.280 307.200 103.450 ;
        RECT 302.110 101.620 302.825 101.790 ;
        RECT 302.110 101.240 302.280 101.620 ;
        RECT 302.495 101.070 302.825 101.450 ;
        RECT 302.995 101.240 303.250 101.815 ;
        RECT 303.425 101.070 303.685 101.910 ;
        RECT 304.325 101.810 304.495 102.480 ;
        RECT 305.170 102.310 305.340 103.280 ;
        RECT 304.665 101.980 304.920 102.310 ;
        RECT 305.145 101.980 305.340 102.310 ;
        RECT 305.510 102.940 306.635 103.110 ;
        RECT 304.750 101.810 304.920 101.980 ;
        RECT 305.510 101.810 305.680 102.940 ;
        RECT 303.860 101.070 304.150 101.795 ;
        RECT 304.325 101.240 304.580 101.810 ;
        RECT 304.750 101.640 305.680 101.810 ;
        RECT 305.850 102.600 306.860 102.770 ;
        RECT 305.850 101.800 306.020 102.600 ;
        RECT 306.225 102.260 306.500 102.400 ;
        RECT 306.220 102.090 306.500 102.260 ;
        RECT 305.505 101.605 305.680 101.640 ;
        RECT 304.750 101.070 305.080 101.470 ;
        RECT 305.505 101.240 306.035 101.605 ;
        RECT 306.225 101.240 306.500 102.090 ;
        RECT 306.670 101.240 306.860 102.600 ;
        RECT 307.030 102.615 307.200 103.280 ;
        RECT 307.370 102.860 307.540 103.620 ;
        RECT 307.775 102.860 308.290 103.270 ;
        RECT 307.030 102.425 307.780 102.615 ;
        RECT 307.950 102.050 308.290 102.860 ;
        RECT 308.460 102.530 309.670 103.620 ;
        RECT 307.060 101.880 308.290 102.050 ;
        RECT 307.040 101.070 307.550 101.605 ;
        RECT 307.770 101.275 308.015 101.880 ;
        RECT 308.460 101.820 308.980 102.360 ;
        RECT 309.150 101.990 309.670 102.530 ;
        RECT 309.840 102.530 311.050 103.620 ;
        RECT 309.840 101.990 310.360 102.530 ;
        RECT 310.530 101.820 311.050 102.360 ;
        RECT 308.460 101.070 309.670 101.820 ;
        RECT 309.840 101.070 311.050 101.820 ;
        RECT 162.095 100.900 311.135 101.070 ;
        RECT 162.180 100.150 163.390 100.900 ;
        RECT 162.180 99.610 162.700 100.150 ;
        RECT 163.565 100.060 163.825 100.900 ;
        RECT 164.000 100.155 164.255 100.730 ;
        RECT 164.425 100.520 164.755 100.900 ;
        RECT 164.970 100.350 165.140 100.730 ;
        RECT 164.425 100.180 165.140 100.350 ;
        RECT 165.490 100.350 165.660 100.730 ;
        RECT 165.875 100.520 166.205 100.900 ;
        RECT 165.490 100.180 166.205 100.350 ;
        RECT 162.870 99.440 163.390 99.980 ;
        RECT 162.180 98.350 163.390 99.440 ;
        RECT 163.565 98.350 163.825 99.500 ;
        RECT 164.000 99.425 164.170 100.155 ;
        RECT 164.425 99.990 164.595 100.180 ;
        RECT 164.340 99.660 164.595 99.990 ;
        RECT 164.425 99.450 164.595 99.660 ;
        RECT 164.875 99.630 165.230 100.000 ;
        RECT 165.400 99.630 165.755 100.000 ;
        RECT 166.035 99.990 166.205 100.180 ;
        RECT 166.375 100.155 166.630 100.730 ;
        RECT 166.035 99.660 166.290 99.990 ;
        RECT 166.035 99.450 166.205 99.660 ;
        RECT 164.000 98.520 164.255 99.425 ;
        RECT 164.425 99.280 165.140 99.450 ;
        RECT 164.425 98.350 164.755 99.110 ;
        RECT 164.970 98.520 165.140 99.280 ;
        RECT 165.490 99.280 166.205 99.450 ;
        RECT 166.460 99.425 166.630 100.155 ;
        RECT 166.805 100.060 167.065 100.900 ;
        RECT 167.245 100.350 167.500 100.640 ;
        RECT 167.670 100.520 168.000 100.900 ;
        RECT 167.245 100.180 167.995 100.350 ;
        RECT 165.490 98.520 165.660 99.280 ;
        RECT 165.875 98.350 166.205 99.110 ;
        RECT 166.375 98.520 166.630 99.425 ;
        RECT 166.805 98.350 167.065 99.500 ;
        RECT 167.245 99.360 167.595 100.010 ;
        RECT 167.765 99.190 167.995 100.180 ;
        RECT 167.245 99.020 167.995 99.190 ;
        RECT 167.245 98.520 167.500 99.020 ;
        RECT 167.670 98.350 168.000 98.850 ;
        RECT 168.170 98.520 168.340 100.640 ;
        RECT 168.700 100.540 169.030 100.900 ;
        RECT 169.200 100.510 169.695 100.680 ;
        RECT 169.900 100.510 170.755 100.680 ;
        RECT 168.570 99.320 169.030 100.370 ;
        RECT 168.510 98.535 168.835 99.320 ;
        RECT 169.200 99.150 169.370 100.510 ;
        RECT 169.540 99.600 169.890 100.220 ;
        RECT 170.060 100.000 170.415 100.220 ;
        RECT 170.060 99.410 170.230 100.000 ;
        RECT 170.585 99.800 170.755 100.510 ;
        RECT 171.630 100.440 171.960 100.900 ;
        RECT 172.170 100.540 172.520 100.710 ;
        RECT 170.960 99.970 171.750 100.220 ;
        RECT 172.170 100.150 172.430 100.540 ;
        RECT 172.740 100.450 173.690 100.730 ;
        RECT 173.860 100.460 174.050 100.900 ;
        RECT 174.220 100.520 175.290 100.690 ;
        RECT 171.920 99.800 172.090 99.980 ;
        RECT 169.200 98.980 169.595 99.150 ;
        RECT 169.765 99.020 170.230 99.410 ;
        RECT 170.400 99.630 172.090 99.800 ;
        RECT 169.425 98.850 169.595 98.980 ;
        RECT 170.400 98.850 170.570 99.630 ;
        RECT 172.260 99.460 172.430 100.150 ;
        RECT 170.930 99.290 172.430 99.460 ;
        RECT 172.620 99.490 172.830 100.280 ;
        RECT 173.000 99.660 173.350 100.280 ;
        RECT 173.520 99.670 173.690 100.450 ;
        RECT 174.220 100.290 174.390 100.520 ;
        RECT 173.860 100.120 174.390 100.290 ;
        RECT 173.860 99.840 174.080 100.120 ;
        RECT 174.560 99.950 174.800 100.350 ;
        RECT 173.520 99.500 173.925 99.670 ;
        RECT 174.260 99.580 174.800 99.950 ;
        RECT 174.970 100.165 175.290 100.520 ;
        RECT 175.535 100.440 175.840 100.900 ;
        RECT 176.010 100.190 176.265 100.720 ;
        RECT 174.970 99.990 175.295 100.165 ;
        RECT 174.970 99.690 175.885 99.990 ;
        RECT 175.145 99.660 175.885 99.690 ;
        RECT 172.620 99.330 173.295 99.490 ;
        RECT 173.755 99.410 173.925 99.500 ;
        RECT 172.620 99.320 173.585 99.330 ;
        RECT 172.260 99.150 172.430 99.290 ;
        RECT 169.005 98.350 169.255 98.810 ;
        RECT 169.425 98.520 169.675 98.850 ;
        RECT 169.890 98.520 170.570 98.850 ;
        RECT 170.740 98.950 171.815 99.120 ;
        RECT 172.260 98.980 172.820 99.150 ;
        RECT 173.125 99.030 173.585 99.320 ;
        RECT 173.755 99.240 174.975 99.410 ;
        RECT 170.740 98.610 170.910 98.950 ;
        RECT 171.145 98.350 171.475 98.780 ;
        RECT 171.645 98.610 171.815 98.950 ;
        RECT 172.110 98.350 172.480 98.810 ;
        RECT 172.650 98.520 172.820 98.980 ;
        RECT 173.755 98.860 173.925 99.240 ;
        RECT 175.145 99.070 175.315 99.660 ;
        RECT 176.055 99.540 176.265 100.190 ;
        RECT 173.055 98.520 173.925 98.860 ;
        RECT 174.515 98.900 175.315 99.070 ;
        RECT 174.095 98.350 174.345 98.810 ;
        RECT 174.515 98.610 174.685 98.900 ;
        RECT 174.865 98.350 175.195 98.730 ;
        RECT 175.535 98.350 175.840 99.490 ;
        RECT 176.010 98.660 176.265 99.540 ;
        RECT 176.445 100.160 176.700 100.730 ;
        RECT 176.870 100.500 177.200 100.900 ;
        RECT 177.625 100.365 178.155 100.730 ;
        RECT 177.625 100.330 177.800 100.365 ;
        RECT 176.870 100.160 177.800 100.330 ;
        RECT 176.445 99.490 176.615 100.160 ;
        RECT 176.870 99.990 177.040 100.160 ;
        RECT 176.785 99.660 177.040 99.990 ;
        RECT 177.265 99.660 177.460 99.990 ;
        RECT 176.445 98.520 176.780 99.490 ;
        RECT 176.950 98.350 177.120 99.490 ;
        RECT 177.290 98.690 177.460 99.660 ;
        RECT 177.630 99.030 177.800 100.160 ;
        RECT 177.970 99.370 178.140 100.170 ;
        RECT 178.345 99.880 178.620 100.730 ;
        RECT 178.340 99.710 178.620 99.880 ;
        RECT 178.345 99.570 178.620 99.710 ;
        RECT 178.790 99.370 178.980 100.730 ;
        RECT 179.160 100.365 179.670 100.900 ;
        RECT 179.890 100.090 180.135 100.695 ;
        RECT 179.180 99.920 180.410 100.090 ;
        RECT 180.585 100.060 180.845 100.900 ;
        RECT 181.020 100.155 181.275 100.730 ;
        RECT 181.445 100.520 181.775 100.900 ;
        RECT 181.990 100.350 182.160 100.730 ;
        RECT 181.445 100.180 182.160 100.350 ;
        RECT 177.970 99.200 178.980 99.370 ;
        RECT 179.150 99.355 179.900 99.545 ;
        RECT 177.630 98.860 178.755 99.030 ;
        RECT 179.150 98.690 179.320 99.355 ;
        RECT 180.070 99.110 180.410 99.920 ;
        RECT 177.290 98.520 179.320 98.690 ;
        RECT 179.490 98.350 179.660 99.110 ;
        RECT 179.895 98.700 180.410 99.110 ;
        RECT 180.585 98.350 180.845 99.500 ;
        RECT 181.020 99.425 181.190 100.155 ;
        RECT 181.445 99.990 181.615 100.180 ;
        RECT 182.885 100.060 183.145 100.900 ;
        RECT 183.320 100.155 183.575 100.730 ;
        RECT 183.745 100.520 184.075 100.900 ;
        RECT 184.290 100.350 184.460 100.730 ;
        RECT 183.745 100.180 184.460 100.350 ;
        RECT 181.360 99.660 181.615 99.990 ;
        RECT 181.445 99.450 181.615 99.660 ;
        RECT 181.895 99.630 182.250 100.000 ;
        RECT 181.020 98.520 181.275 99.425 ;
        RECT 181.445 99.280 182.160 99.450 ;
        RECT 181.445 98.350 181.775 99.110 ;
        RECT 181.990 98.520 182.160 99.280 ;
        RECT 182.885 98.350 183.145 99.500 ;
        RECT 183.320 99.425 183.490 100.155 ;
        RECT 183.745 99.990 183.915 100.180 ;
        RECT 185.185 100.060 185.445 100.900 ;
        RECT 185.620 100.155 185.875 100.730 ;
        RECT 186.045 100.520 186.375 100.900 ;
        RECT 186.590 100.350 186.760 100.730 ;
        RECT 186.045 100.180 186.760 100.350 ;
        RECT 183.660 99.660 183.915 99.990 ;
        RECT 183.745 99.450 183.915 99.660 ;
        RECT 184.195 99.630 184.550 100.000 ;
        RECT 183.320 98.520 183.575 99.425 ;
        RECT 183.745 99.280 184.460 99.450 ;
        RECT 183.745 98.350 184.075 99.110 ;
        RECT 184.290 98.520 184.460 99.280 ;
        RECT 185.185 98.350 185.445 99.500 ;
        RECT 185.620 99.425 185.790 100.155 ;
        RECT 186.045 99.990 186.215 100.180 ;
        RECT 187.940 100.175 188.230 100.900 ;
        RECT 188.405 100.350 188.660 100.640 ;
        RECT 188.830 100.520 189.160 100.900 ;
        RECT 188.405 100.180 189.155 100.350 ;
        RECT 185.960 99.660 186.215 99.990 ;
        RECT 186.045 99.450 186.215 99.660 ;
        RECT 186.495 99.630 186.850 100.000 ;
        RECT 185.620 98.520 185.875 99.425 ;
        RECT 186.045 99.280 186.760 99.450 ;
        RECT 186.045 98.350 186.375 99.110 ;
        RECT 186.590 98.520 186.760 99.280 ;
        RECT 187.940 98.350 188.230 99.515 ;
        RECT 188.405 99.360 188.755 100.010 ;
        RECT 188.925 99.190 189.155 100.180 ;
        RECT 188.405 99.020 189.155 99.190 ;
        RECT 188.405 98.520 188.660 99.020 ;
        RECT 188.830 98.350 189.160 98.850 ;
        RECT 189.330 98.520 189.500 100.640 ;
        RECT 189.860 100.540 190.190 100.900 ;
        RECT 190.360 100.510 190.855 100.680 ;
        RECT 191.060 100.510 191.915 100.680 ;
        RECT 189.730 99.320 190.190 100.370 ;
        RECT 189.670 98.535 189.995 99.320 ;
        RECT 190.360 99.150 190.530 100.510 ;
        RECT 190.700 99.600 191.050 100.220 ;
        RECT 191.220 100.000 191.575 100.220 ;
        RECT 191.220 99.410 191.390 100.000 ;
        RECT 191.745 99.800 191.915 100.510 ;
        RECT 192.790 100.440 193.120 100.900 ;
        RECT 193.330 100.540 193.680 100.710 ;
        RECT 192.120 99.970 192.910 100.220 ;
        RECT 193.330 100.150 193.590 100.540 ;
        RECT 193.900 100.450 194.850 100.730 ;
        RECT 195.020 100.460 195.210 100.900 ;
        RECT 195.380 100.520 196.450 100.690 ;
        RECT 193.080 99.800 193.250 99.980 ;
        RECT 190.360 98.980 190.755 99.150 ;
        RECT 190.925 99.020 191.390 99.410 ;
        RECT 191.560 99.630 193.250 99.800 ;
        RECT 190.585 98.850 190.755 98.980 ;
        RECT 191.560 98.850 191.730 99.630 ;
        RECT 193.420 99.460 193.590 100.150 ;
        RECT 192.090 99.290 193.590 99.460 ;
        RECT 193.780 99.490 193.990 100.280 ;
        RECT 194.160 99.660 194.510 100.280 ;
        RECT 194.680 99.670 194.850 100.450 ;
        RECT 195.380 100.290 195.550 100.520 ;
        RECT 195.020 100.120 195.550 100.290 ;
        RECT 195.020 99.840 195.240 100.120 ;
        RECT 195.720 99.950 195.960 100.350 ;
        RECT 194.680 99.500 195.085 99.670 ;
        RECT 195.420 99.580 195.960 99.950 ;
        RECT 196.130 100.165 196.450 100.520 ;
        RECT 196.695 100.440 197.000 100.900 ;
        RECT 197.170 100.190 197.425 100.720 ;
        RECT 196.130 99.990 196.455 100.165 ;
        RECT 196.130 99.690 197.045 99.990 ;
        RECT 196.305 99.660 197.045 99.690 ;
        RECT 193.780 99.330 194.455 99.490 ;
        RECT 194.915 99.410 195.085 99.500 ;
        RECT 193.780 99.320 194.745 99.330 ;
        RECT 193.420 99.150 193.590 99.290 ;
        RECT 190.165 98.350 190.415 98.810 ;
        RECT 190.585 98.520 190.835 98.850 ;
        RECT 191.050 98.520 191.730 98.850 ;
        RECT 191.900 98.950 192.975 99.120 ;
        RECT 193.420 98.980 193.980 99.150 ;
        RECT 194.285 99.030 194.745 99.320 ;
        RECT 194.915 99.240 196.135 99.410 ;
        RECT 191.900 98.610 192.070 98.950 ;
        RECT 192.305 98.350 192.635 98.780 ;
        RECT 192.805 98.610 192.975 98.950 ;
        RECT 193.270 98.350 193.640 98.810 ;
        RECT 193.810 98.520 193.980 98.980 ;
        RECT 194.915 98.860 195.085 99.240 ;
        RECT 196.305 99.070 196.475 99.660 ;
        RECT 197.215 99.540 197.425 100.190 ;
        RECT 197.600 100.130 201.110 100.900 ;
        RECT 201.280 100.150 202.490 100.900 ;
        RECT 202.665 100.190 202.920 100.720 ;
        RECT 203.090 100.440 203.395 100.900 ;
        RECT 203.640 100.520 204.710 100.690 ;
        RECT 197.600 99.610 199.250 100.130 ;
        RECT 194.215 98.520 195.085 98.860 ;
        RECT 195.675 98.900 196.475 99.070 ;
        RECT 195.255 98.350 195.505 98.810 ;
        RECT 195.675 98.610 195.845 98.900 ;
        RECT 196.025 98.350 196.355 98.730 ;
        RECT 196.695 98.350 197.000 99.490 ;
        RECT 197.170 98.660 197.425 99.540 ;
        RECT 199.420 99.440 201.110 99.960 ;
        RECT 201.280 99.610 201.800 100.150 ;
        RECT 201.970 99.440 202.490 99.980 ;
        RECT 197.600 98.350 201.110 99.440 ;
        RECT 201.280 98.350 202.490 99.440 ;
        RECT 202.665 99.540 202.875 100.190 ;
        RECT 203.640 100.165 203.960 100.520 ;
        RECT 203.635 99.990 203.960 100.165 ;
        RECT 203.045 99.690 203.960 99.990 ;
        RECT 204.130 99.950 204.370 100.350 ;
        RECT 204.540 100.290 204.710 100.520 ;
        RECT 204.880 100.460 205.070 100.900 ;
        RECT 205.240 100.450 206.190 100.730 ;
        RECT 206.410 100.540 206.760 100.710 ;
        RECT 204.540 100.120 205.070 100.290 ;
        RECT 203.045 99.660 203.785 99.690 ;
        RECT 202.665 98.660 202.920 99.540 ;
        RECT 203.090 98.350 203.395 99.490 ;
        RECT 203.615 99.070 203.785 99.660 ;
        RECT 204.130 99.580 204.670 99.950 ;
        RECT 204.850 99.840 205.070 100.120 ;
        RECT 205.240 99.670 205.410 100.450 ;
        RECT 205.005 99.500 205.410 99.670 ;
        RECT 205.580 99.660 205.930 100.280 ;
        RECT 205.005 99.410 205.175 99.500 ;
        RECT 206.100 99.490 206.310 100.280 ;
        RECT 203.955 99.240 205.175 99.410 ;
        RECT 205.635 99.330 206.310 99.490 ;
        RECT 203.615 98.900 204.415 99.070 ;
        RECT 203.735 98.350 204.065 98.730 ;
        RECT 204.245 98.610 204.415 98.900 ;
        RECT 205.005 98.860 205.175 99.240 ;
        RECT 205.345 99.320 206.310 99.330 ;
        RECT 206.500 100.150 206.760 100.540 ;
        RECT 206.970 100.440 207.300 100.900 ;
        RECT 208.175 100.510 209.030 100.680 ;
        RECT 209.235 100.510 209.730 100.680 ;
        RECT 209.900 100.540 210.230 100.900 ;
        RECT 206.500 99.460 206.670 100.150 ;
        RECT 206.840 99.800 207.010 99.980 ;
        RECT 207.180 99.970 207.970 100.220 ;
        RECT 208.175 99.800 208.345 100.510 ;
        RECT 208.515 100.000 208.870 100.220 ;
        RECT 206.840 99.630 208.530 99.800 ;
        RECT 205.345 99.030 205.805 99.320 ;
        RECT 206.500 99.290 208.000 99.460 ;
        RECT 206.500 99.150 206.670 99.290 ;
        RECT 206.110 98.980 206.670 99.150 ;
        RECT 204.585 98.350 204.835 98.810 ;
        RECT 205.005 98.520 205.875 98.860 ;
        RECT 206.110 98.520 206.280 98.980 ;
        RECT 207.115 98.950 208.190 99.120 ;
        RECT 206.450 98.350 206.820 98.810 ;
        RECT 207.115 98.610 207.285 98.950 ;
        RECT 207.455 98.350 207.785 98.780 ;
        RECT 208.020 98.610 208.190 98.950 ;
        RECT 208.360 98.850 208.530 99.630 ;
        RECT 208.700 99.410 208.870 100.000 ;
        RECT 209.040 99.600 209.390 100.220 ;
        RECT 208.700 99.020 209.165 99.410 ;
        RECT 209.560 99.150 209.730 100.510 ;
        RECT 209.900 99.320 210.360 100.370 ;
        RECT 209.335 98.980 209.730 99.150 ;
        RECT 209.335 98.850 209.505 98.980 ;
        RECT 208.360 98.520 209.040 98.850 ;
        RECT 209.255 98.520 209.505 98.850 ;
        RECT 209.675 98.350 209.925 98.810 ;
        RECT 210.095 98.535 210.420 99.320 ;
        RECT 210.590 98.520 210.760 100.640 ;
        RECT 210.930 100.520 211.260 100.900 ;
        RECT 211.430 100.350 211.685 100.640 ;
        RECT 210.935 100.180 211.685 100.350 ;
        RECT 210.935 99.190 211.165 100.180 ;
        RECT 211.865 100.060 212.125 100.900 ;
        RECT 212.300 100.155 212.555 100.730 ;
        RECT 212.725 100.520 213.055 100.900 ;
        RECT 213.270 100.350 213.440 100.730 ;
        RECT 212.725 100.180 213.440 100.350 ;
        RECT 211.335 99.360 211.685 100.010 ;
        RECT 210.935 99.020 211.685 99.190 ;
        RECT 210.930 98.350 211.260 98.850 ;
        RECT 211.430 98.520 211.685 99.020 ;
        RECT 211.865 98.350 212.125 99.500 ;
        RECT 212.300 99.425 212.470 100.155 ;
        RECT 212.725 99.990 212.895 100.180 ;
        RECT 213.700 100.175 213.990 100.900 ;
        RECT 215.085 100.060 215.345 100.900 ;
        RECT 215.520 100.155 215.775 100.730 ;
        RECT 215.945 100.520 216.275 100.900 ;
        RECT 216.490 100.350 216.660 100.730 ;
        RECT 215.945 100.180 216.660 100.350 ;
        RECT 217.385 100.350 217.640 100.640 ;
        RECT 217.810 100.520 218.140 100.900 ;
        RECT 217.385 100.180 218.135 100.350 ;
        RECT 212.640 99.660 212.895 99.990 ;
        RECT 212.725 99.450 212.895 99.660 ;
        RECT 213.175 99.630 213.530 100.000 ;
        RECT 212.300 98.520 212.555 99.425 ;
        RECT 212.725 99.280 213.440 99.450 ;
        RECT 212.725 98.350 213.055 99.110 ;
        RECT 213.270 98.520 213.440 99.280 ;
        RECT 213.700 98.350 213.990 99.515 ;
        RECT 215.085 98.350 215.345 99.500 ;
        RECT 215.520 99.425 215.690 100.155 ;
        RECT 215.945 99.990 216.115 100.180 ;
        RECT 215.860 99.660 216.115 99.990 ;
        RECT 215.945 99.450 216.115 99.660 ;
        RECT 216.395 99.630 216.750 100.000 ;
        RECT 215.520 98.520 215.775 99.425 ;
        RECT 215.945 99.280 216.660 99.450 ;
        RECT 217.385 99.360 217.735 100.010 ;
        RECT 215.945 98.350 216.275 99.110 ;
        RECT 216.490 98.520 216.660 99.280 ;
        RECT 217.905 99.190 218.135 100.180 ;
        RECT 217.385 99.020 218.135 99.190 ;
        RECT 217.385 98.520 217.640 99.020 ;
        RECT 217.810 98.350 218.140 98.850 ;
        RECT 218.310 98.520 218.480 100.640 ;
        RECT 218.840 100.540 219.170 100.900 ;
        RECT 219.340 100.510 219.835 100.680 ;
        RECT 220.040 100.510 220.895 100.680 ;
        RECT 218.710 99.320 219.170 100.370 ;
        RECT 218.650 98.535 218.975 99.320 ;
        RECT 219.340 99.150 219.510 100.510 ;
        RECT 219.680 99.600 220.030 100.220 ;
        RECT 220.200 100.000 220.555 100.220 ;
        RECT 220.200 99.410 220.370 100.000 ;
        RECT 220.725 99.800 220.895 100.510 ;
        RECT 221.770 100.440 222.100 100.900 ;
        RECT 222.310 100.540 222.660 100.710 ;
        RECT 221.100 99.970 221.890 100.220 ;
        RECT 222.310 100.150 222.570 100.540 ;
        RECT 222.880 100.450 223.830 100.730 ;
        RECT 224.000 100.460 224.190 100.900 ;
        RECT 224.360 100.520 225.430 100.690 ;
        RECT 222.060 99.800 222.230 99.980 ;
        RECT 219.340 98.980 219.735 99.150 ;
        RECT 219.905 99.020 220.370 99.410 ;
        RECT 220.540 99.630 222.230 99.800 ;
        RECT 219.565 98.850 219.735 98.980 ;
        RECT 220.540 98.850 220.710 99.630 ;
        RECT 222.400 99.460 222.570 100.150 ;
        RECT 221.070 99.290 222.570 99.460 ;
        RECT 222.760 99.490 222.970 100.280 ;
        RECT 223.140 99.660 223.490 100.280 ;
        RECT 223.660 99.670 223.830 100.450 ;
        RECT 224.360 100.290 224.530 100.520 ;
        RECT 224.000 100.120 224.530 100.290 ;
        RECT 224.000 99.840 224.220 100.120 ;
        RECT 224.700 99.950 224.940 100.350 ;
        RECT 223.660 99.500 224.065 99.670 ;
        RECT 224.400 99.580 224.940 99.950 ;
        RECT 225.110 100.165 225.430 100.520 ;
        RECT 225.675 100.440 225.980 100.900 ;
        RECT 226.150 100.190 226.405 100.720 ;
        RECT 225.110 99.990 225.435 100.165 ;
        RECT 225.110 99.690 226.025 99.990 ;
        RECT 225.285 99.660 226.025 99.690 ;
        RECT 222.760 99.330 223.435 99.490 ;
        RECT 223.895 99.410 224.065 99.500 ;
        RECT 222.760 99.320 223.725 99.330 ;
        RECT 222.400 99.150 222.570 99.290 ;
        RECT 219.145 98.350 219.395 98.810 ;
        RECT 219.565 98.520 219.815 98.850 ;
        RECT 220.030 98.520 220.710 98.850 ;
        RECT 220.880 98.950 221.955 99.120 ;
        RECT 222.400 98.980 222.960 99.150 ;
        RECT 223.265 99.030 223.725 99.320 ;
        RECT 223.895 99.240 225.115 99.410 ;
        RECT 220.880 98.610 221.050 98.950 ;
        RECT 221.285 98.350 221.615 98.780 ;
        RECT 221.785 98.610 221.955 98.950 ;
        RECT 222.250 98.350 222.620 98.810 ;
        RECT 222.790 98.520 222.960 98.980 ;
        RECT 223.895 98.860 224.065 99.240 ;
        RECT 225.285 99.070 225.455 99.660 ;
        RECT 226.195 99.540 226.405 100.190 ;
        RECT 226.580 100.150 227.790 100.900 ;
        RECT 228.050 100.250 228.220 100.730 ;
        RECT 228.390 100.420 228.720 100.900 ;
        RECT 228.945 100.480 230.480 100.730 ;
        RECT 228.945 100.250 229.115 100.480 ;
        RECT 226.580 99.610 227.100 100.150 ;
        RECT 228.050 100.080 229.115 100.250 ;
        RECT 223.195 98.520 224.065 98.860 ;
        RECT 224.655 98.900 225.455 99.070 ;
        RECT 224.235 98.350 224.485 98.810 ;
        RECT 224.655 98.610 224.825 98.900 ;
        RECT 225.005 98.350 225.335 98.730 ;
        RECT 225.675 98.350 225.980 99.490 ;
        RECT 226.150 98.660 226.405 99.540 ;
        RECT 227.270 99.440 227.790 99.980 ;
        RECT 229.295 99.910 229.575 100.310 ;
        RECT 227.965 99.700 228.315 99.910 ;
        RECT 228.485 99.710 228.930 99.910 ;
        RECT 229.100 99.710 229.575 99.910 ;
        RECT 229.845 99.910 230.130 100.310 ;
        RECT 230.310 100.250 230.480 100.480 ;
        RECT 230.650 100.420 230.980 100.900 ;
        RECT 231.195 100.400 231.450 100.730 ;
        RECT 231.265 100.320 231.450 100.400 ;
        RECT 231.640 100.355 236.985 100.900 ;
        RECT 230.310 100.080 231.110 100.250 ;
        RECT 229.845 99.710 230.175 99.910 ;
        RECT 230.345 99.710 230.710 99.910 ;
        RECT 230.940 99.530 231.110 100.080 ;
        RECT 226.580 98.350 227.790 99.440 ;
        RECT 228.050 99.360 231.110 99.530 ;
        RECT 228.050 98.520 228.220 99.360 ;
        RECT 231.280 99.190 231.450 100.320 ;
        RECT 233.225 99.525 233.565 100.355 ;
        RECT 237.160 100.130 238.830 100.900 ;
        RECT 239.460 100.175 239.750 100.900 ;
        RECT 239.925 100.350 240.180 100.640 ;
        RECT 240.350 100.520 240.680 100.900 ;
        RECT 239.925 100.180 240.675 100.350 ;
        RECT 228.390 98.690 228.720 99.190 ;
        RECT 228.890 98.950 230.525 99.190 ;
        RECT 228.890 98.860 229.120 98.950 ;
        RECT 229.230 98.690 229.560 98.730 ;
        RECT 228.390 98.520 229.560 98.690 ;
        RECT 229.750 98.350 230.105 98.770 ;
        RECT 230.275 98.520 230.525 98.950 ;
        RECT 230.695 98.350 231.025 99.110 ;
        RECT 231.195 98.520 231.450 99.190 ;
        RECT 235.045 98.785 235.395 100.035 ;
        RECT 237.160 99.610 237.910 100.130 ;
        RECT 238.080 99.440 238.830 99.960 ;
        RECT 231.640 98.350 236.985 98.785 ;
        RECT 237.160 98.350 238.830 99.440 ;
        RECT 239.460 98.350 239.750 99.515 ;
        RECT 239.925 99.360 240.275 100.010 ;
        RECT 240.445 99.190 240.675 100.180 ;
        RECT 239.925 99.020 240.675 99.190 ;
        RECT 239.925 98.520 240.180 99.020 ;
        RECT 240.350 98.350 240.680 98.850 ;
        RECT 240.850 98.520 241.020 100.640 ;
        RECT 241.380 100.540 241.710 100.900 ;
        RECT 241.880 100.510 242.375 100.680 ;
        RECT 242.580 100.510 243.435 100.680 ;
        RECT 241.250 99.320 241.710 100.370 ;
        RECT 241.190 98.535 241.515 99.320 ;
        RECT 241.880 99.150 242.050 100.510 ;
        RECT 242.220 99.600 242.570 100.220 ;
        RECT 242.740 100.000 243.095 100.220 ;
        RECT 242.740 99.410 242.910 100.000 ;
        RECT 243.265 99.800 243.435 100.510 ;
        RECT 244.310 100.440 244.640 100.900 ;
        RECT 244.850 100.540 245.200 100.710 ;
        RECT 243.640 99.970 244.430 100.220 ;
        RECT 244.850 100.150 245.110 100.540 ;
        RECT 245.420 100.450 246.370 100.730 ;
        RECT 246.540 100.460 246.730 100.900 ;
        RECT 246.900 100.520 247.970 100.690 ;
        RECT 244.600 99.800 244.770 99.980 ;
        RECT 241.880 98.980 242.275 99.150 ;
        RECT 242.445 99.020 242.910 99.410 ;
        RECT 243.080 99.630 244.770 99.800 ;
        RECT 242.105 98.850 242.275 98.980 ;
        RECT 243.080 98.850 243.250 99.630 ;
        RECT 244.940 99.460 245.110 100.150 ;
        RECT 243.610 99.290 245.110 99.460 ;
        RECT 245.300 99.490 245.510 100.280 ;
        RECT 245.680 99.660 246.030 100.280 ;
        RECT 246.200 99.670 246.370 100.450 ;
        RECT 246.900 100.290 247.070 100.520 ;
        RECT 246.540 100.120 247.070 100.290 ;
        RECT 246.540 99.840 246.760 100.120 ;
        RECT 247.240 99.950 247.480 100.350 ;
        RECT 246.200 99.500 246.605 99.670 ;
        RECT 246.940 99.580 247.480 99.950 ;
        RECT 247.650 100.165 247.970 100.520 ;
        RECT 248.215 100.440 248.520 100.900 ;
        RECT 248.690 100.190 248.945 100.720 ;
        RECT 247.650 99.990 247.975 100.165 ;
        RECT 247.650 99.690 248.565 99.990 ;
        RECT 247.825 99.660 248.565 99.690 ;
        RECT 245.300 99.330 245.975 99.490 ;
        RECT 246.435 99.410 246.605 99.500 ;
        RECT 245.300 99.320 246.265 99.330 ;
        RECT 244.940 99.150 245.110 99.290 ;
        RECT 241.685 98.350 241.935 98.810 ;
        RECT 242.105 98.520 242.355 98.850 ;
        RECT 242.570 98.520 243.250 98.850 ;
        RECT 243.420 98.950 244.495 99.120 ;
        RECT 244.940 98.980 245.500 99.150 ;
        RECT 245.805 99.030 246.265 99.320 ;
        RECT 246.435 99.240 247.655 99.410 ;
        RECT 243.420 98.610 243.590 98.950 ;
        RECT 243.825 98.350 244.155 98.780 ;
        RECT 244.325 98.610 244.495 98.950 ;
        RECT 244.790 98.350 245.160 98.810 ;
        RECT 245.330 98.520 245.500 98.980 ;
        RECT 246.435 98.860 246.605 99.240 ;
        RECT 247.825 99.070 247.995 99.660 ;
        RECT 248.735 99.540 248.945 100.190 ;
        RECT 249.125 100.135 249.580 100.900 ;
        RECT 249.855 100.520 251.155 100.730 ;
        RECT 251.410 100.540 251.740 100.900 ;
        RECT 250.985 100.370 251.155 100.520 ;
        RECT 251.910 100.400 252.170 100.730 ;
        RECT 250.055 99.910 250.275 100.310 ;
        RECT 249.120 99.710 249.610 99.910 ;
        RECT 249.800 99.700 250.275 99.910 ;
        RECT 250.520 99.910 250.730 100.310 ;
        RECT 250.985 100.245 251.740 100.370 ;
        RECT 250.985 100.200 251.830 100.245 ;
        RECT 251.560 100.080 251.830 100.200 ;
        RECT 250.520 99.700 250.850 99.910 ;
        RECT 251.020 99.640 251.430 99.945 ;
        RECT 245.735 98.520 246.605 98.860 ;
        RECT 247.195 98.900 247.995 99.070 ;
        RECT 246.775 98.350 247.025 98.810 ;
        RECT 247.195 98.610 247.365 98.900 ;
        RECT 247.545 98.350 247.875 98.730 ;
        RECT 248.215 98.350 248.520 99.490 ;
        RECT 248.690 98.660 248.945 99.540 ;
        RECT 249.125 99.470 250.300 99.530 ;
        RECT 251.660 99.505 251.830 100.080 ;
        RECT 251.630 99.470 251.830 99.505 ;
        RECT 249.125 99.360 251.830 99.470 ;
        RECT 249.125 98.740 249.380 99.360 ;
        RECT 249.970 99.300 251.770 99.360 ;
        RECT 249.970 99.270 250.300 99.300 ;
        RECT 252.000 99.200 252.170 100.400 ;
        RECT 249.630 99.100 249.815 99.190 ;
        RECT 250.405 99.100 251.240 99.110 ;
        RECT 249.630 98.900 251.240 99.100 ;
        RECT 249.630 98.860 249.860 98.900 ;
        RECT 249.125 98.520 249.460 98.740 ;
        RECT 250.465 98.350 250.820 98.730 ;
        RECT 250.990 98.520 251.240 98.900 ;
        RECT 251.490 98.350 251.740 99.130 ;
        RECT 251.910 98.520 252.170 99.200 ;
        RECT 252.345 100.160 252.600 100.730 ;
        RECT 252.770 100.500 253.100 100.900 ;
        RECT 253.525 100.365 254.055 100.730 ;
        RECT 253.525 100.330 253.700 100.365 ;
        RECT 252.770 100.160 253.700 100.330 ;
        RECT 252.345 99.490 252.515 100.160 ;
        RECT 252.770 99.990 252.940 100.160 ;
        RECT 252.685 99.660 252.940 99.990 ;
        RECT 253.165 99.660 253.360 99.990 ;
        RECT 252.345 98.520 252.680 99.490 ;
        RECT 252.850 98.350 253.020 99.490 ;
        RECT 253.190 98.690 253.360 99.660 ;
        RECT 253.530 99.030 253.700 100.160 ;
        RECT 253.870 99.370 254.040 100.170 ;
        RECT 254.245 99.880 254.520 100.730 ;
        RECT 254.240 99.710 254.520 99.880 ;
        RECT 254.245 99.570 254.520 99.710 ;
        RECT 254.690 99.370 254.880 100.730 ;
        RECT 255.060 100.365 255.570 100.900 ;
        RECT 255.790 100.090 256.035 100.695 ;
        RECT 255.080 99.920 256.310 100.090 ;
        RECT 256.485 100.060 256.745 100.900 ;
        RECT 256.920 100.155 257.175 100.730 ;
        RECT 257.345 100.520 257.675 100.900 ;
        RECT 257.890 100.350 258.060 100.730 ;
        RECT 257.345 100.180 258.060 100.350 ;
        RECT 253.870 99.200 254.880 99.370 ;
        RECT 255.050 99.355 255.800 99.545 ;
        RECT 253.530 98.860 254.655 99.030 ;
        RECT 255.050 98.690 255.220 99.355 ;
        RECT 255.970 99.110 256.310 99.920 ;
        RECT 253.190 98.520 255.220 98.690 ;
        RECT 255.390 98.350 255.560 99.110 ;
        RECT 255.795 98.700 256.310 99.110 ;
        RECT 256.485 98.350 256.745 99.500 ;
        RECT 256.920 99.425 257.090 100.155 ;
        RECT 257.345 99.990 257.515 100.180 ;
        RECT 258.595 100.090 258.840 100.695 ;
        RECT 259.060 100.365 259.570 100.900 ;
        RECT 257.260 99.660 257.515 99.990 ;
        RECT 257.345 99.450 257.515 99.660 ;
        RECT 257.795 99.630 258.150 100.000 ;
        RECT 258.320 99.920 259.550 100.090 ;
        RECT 256.920 98.520 257.175 99.425 ;
        RECT 257.345 99.280 258.060 99.450 ;
        RECT 257.345 98.350 257.675 99.110 ;
        RECT 257.890 98.520 258.060 99.280 ;
        RECT 258.320 99.110 258.660 99.920 ;
        RECT 258.830 99.355 259.580 99.545 ;
        RECT 258.320 98.700 258.835 99.110 ;
        RECT 259.070 98.350 259.240 99.110 ;
        RECT 259.410 98.690 259.580 99.355 ;
        RECT 259.750 99.370 259.940 100.730 ;
        RECT 260.110 99.880 260.385 100.730 ;
        RECT 260.575 100.365 261.105 100.730 ;
        RECT 261.530 100.500 261.860 100.900 ;
        RECT 260.930 100.330 261.105 100.365 ;
        RECT 260.110 99.710 260.390 99.880 ;
        RECT 260.110 99.570 260.385 99.710 ;
        RECT 260.590 99.370 260.760 100.170 ;
        RECT 259.750 99.200 260.760 99.370 ;
        RECT 260.930 100.160 261.860 100.330 ;
        RECT 262.030 100.160 262.285 100.730 ;
        RECT 260.930 99.030 261.100 100.160 ;
        RECT 261.690 99.990 261.860 100.160 ;
        RECT 259.975 98.860 261.100 99.030 ;
        RECT 261.270 99.660 261.465 99.990 ;
        RECT 261.690 99.660 261.945 99.990 ;
        RECT 261.270 98.690 261.440 99.660 ;
        RECT 262.115 99.490 262.285 100.160 ;
        RECT 262.465 100.060 262.725 100.900 ;
        RECT 262.900 100.155 263.155 100.730 ;
        RECT 263.325 100.520 263.655 100.900 ;
        RECT 263.870 100.350 264.040 100.730 ;
        RECT 263.325 100.180 264.040 100.350 ;
        RECT 259.410 98.520 261.440 98.690 ;
        RECT 261.610 98.350 261.780 99.490 ;
        RECT 261.950 98.520 262.285 99.490 ;
        RECT 262.465 98.350 262.725 99.500 ;
        RECT 262.900 99.425 263.070 100.155 ;
        RECT 263.325 99.990 263.495 100.180 ;
        RECT 265.220 100.175 265.510 100.900 ;
        RECT 265.685 100.190 265.940 100.720 ;
        RECT 266.110 100.440 266.415 100.900 ;
        RECT 266.660 100.520 267.730 100.690 ;
        RECT 263.240 99.660 263.495 99.990 ;
        RECT 263.325 99.450 263.495 99.660 ;
        RECT 263.775 99.630 264.130 100.000 ;
        RECT 265.685 99.540 265.895 100.190 ;
        RECT 266.660 100.165 266.980 100.520 ;
        RECT 266.655 99.990 266.980 100.165 ;
        RECT 266.065 99.690 266.980 99.990 ;
        RECT 267.150 99.950 267.390 100.350 ;
        RECT 267.560 100.290 267.730 100.520 ;
        RECT 267.900 100.460 268.090 100.900 ;
        RECT 268.260 100.450 269.210 100.730 ;
        RECT 269.430 100.540 269.780 100.710 ;
        RECT 267.560 100.120 268.090 100.290 ;
        RECT 266.065 99.660 266.805 99.690 ;
        RECT 262.900 98.520 263.155 99.425 ;
        RECT 263.325 99.280 264.040 99.450 ;
        RECT 263.325 98.350 263.655 99.110 ;
        RECT 263.870 98.520 264.040 99.280 ;
        RECT 265.220 98.350 265.510 99.515 ;
        RECT 265.685 98.660 265.940 99.540 ;
        RECT 266.110 98.350 266.415 99.490 ;
        RECT 266.635 99.070 266.805 99.660 ;
        RECT 267.150 99.580 267.690 99.950 ;
        RECT 267.870 99.840 268.090 100.120 ;
        RECT 268.260 99.670 268.430 100.450 ;
        RECT 268.025 99.500 268.430 99.670 ;
        RECT 268.600 99.660 268.950 100.280 ;
        RECT 268.025 99.410 268.195 99.500 ;
        RECT 269.120 99.490 269.330 100.280 ;
        RECT 266.975 99.240 268.195 99.410 ;
        RECT 268.655 99.330 269.330 99.490 ;
        RECT 266.635 98.900 267.435 99.070 ;
        RECT 266.755 98.350 267.085 98.730 ;
        RECT 267.265 98.610 267.435 98.900 ;
        RECT 268.025 98.860 268.195 99.240 ;
        RECT 268.365 99.320 269.330 99.330 ;
        RECT 269.520 100.150 269.780 100.540 ;
        RECT 269.990 100.440 270.320 100.900 ;
        RECT 271.195 100.510 272.050 100.680 ;
        RECT 272.255 100.510 272.750 100.680 ;
        RECT 272.920 100.540 273.250 100.900 ;
        RECT 269.520 99.460 269.690 100.150 ;
        RECT 269.860 99.800 270.030 99.980 ;
        RECT 270.200 99.970 270.990 100.220 ;
        RECT 271.195 99.800 271.365 100.510 ;
        RECT 271.535 100.000 271.890 100.220 ;
        RECT 269.860 99.630 271.550 99.800 ;
        RECT 268.365 99.030 268.825 99.320 ;
        RECT 269.520 99.290 271.020 99.460 ;
        RECT 269.520 99.150 269.690 99.290 ;
        RECT 269.130 98.980 269.690 99.150 ;
        RECT 267.605 98.350 267.855 98.810 ;
        RECT 268.025 98.520 268.895 98.860 ;
        RECT 269.130 98.520 269.300 98.980 ;
        RECT 270.135 98.950 271.210 99.120 ;
        RECT 269.470 98.350 269.840 98.810 ;
        RECT 270.135 98.610 270.305 98.950 ;
        RECT 270.475 98.350 270.805 98.780 ;
        RECT 271.040 98.610 271.210 98.950 ;
        RECT 271.380 98.850 271.550 99.630 ;
        RECT 271.720 99.410 271.890 100.000 ;
        RECT 272.060 99.600 272.410 100.220 ;
        RECT 271.720 99.020 272.185 99.410 ;
        RECT 272.580 99.150 272.750 100.510 ;
        RECT 272.920 99.320 273.380 100.370 ;
        RECT 272.355 98.980 272.750 99.150 ;
        RECT 272.355 98.850 272.525 98.980 ;
        RECT 271.380 98.520 272.060 98.850 ;
        RECT 272.275 98.520 272.525 98.850 ;
        RECT 272.695 98.350 272.945 98.810 ;
        RECT 273.115 98.535 273.440 99.320 ;
        RECT 273.610 98.520 273.780 100.640 ;
        RECT 273.950 100.520 274.280 100.900 ;
        RECT 274.450 100.350 274.705 100.640 ;
        RECT 273.955 100.180 274.705 100.350 ;
        RECT 274.885 100.350 275.140 100.640 ;
        RECT 275.310 100.520 275.640 100.900 ;
        RECT 274.885 100.180 275.635 100.350 ;
        RECT 273.955 99.190 274.185 100.180 ;
        RECT 274.355 99.360 274.705 100.010 ;
        RECT 274.885 99.360 275.235 100.010 ;
        RECT 275.405 99.190 275.635 100.180 ;
        RECT 273.955 99.020 274.705 99.190 ;
        RECT 273.950 98.350 274.280 98.850 ;
        RECT 274.450 98.520 274.705 99.020 ;
        RECT 274.885 99.020 275.635 99.190 ;
        RECT 274.885 98.520 275.140 99.020 ;
        RECT 275.310 98.350 275.640 98.850 ;
        RECT 275.810 98.520 275.980 100.640 ;
        RECT 276.340 100.540 276.670 100.900 ;
        RECT 276.840 100.510 277.335 100.680 ;
        RECT 277.540 100.510 278.395 100.680 ;
        RECT 276.210 99.320 276.670 100.370 ;
        RECT 276.150 98.535 276.475 99.320 ;
        RECT 276.840 99.150 277.010 100.510 ;
        RECT 277.180 99.600 277.530 100.220 ;
        RECT 277.700 100.000 278.055 100.220 ;
        RECT 277.700 99.410 277.870 100.000 ;
        RECT 278.225 99.800 278.395 100.510 ;
        RECT 279.270 100.440 279.600 100.900 ;
        RECT 279.810 100.540 280.160 100.710 ;
        RECT 278.600 99.970 279.390 100.220 ;
        RECT 279.810 100.150 280.070 100.540 ;
        RECT 280.380 100.450 281.330 100.730 ;
        RECT 281.500 100.460 281.690 100.900 ;
        RECT 281.860 100.520 282.930 100.690 ;
        RECT 279.560 99.800 279.730 99.980 ;
        RECT 276.840 98.980 277.235 99.150 ;
        RECT 277.405 99.020 277.870 99.410 ;
        RECT 278.040 99.630 279.730 99.800 ;
        RECT 277.065 98.850 277.235 98.980 ;
        RECT 278.040 98.850 278.210 99.630 ;
        RECT 279.900 99.460 280.070 100.150 ;
        RECT 278.570 99.290 280.070 99.460 ;
        RECT 280.260 99.490 280.470 100.280 ;
        RECT 280.640 99.660 280.990 100.280 ;
        RECT 281.160 99.670 281.330 100.450 ;
        RECT 281.860 100.290 282.030 100.520 ;
        RECT 281.500 100.120 282.030 100.290 ;
        RECT 281.500 99.840 281.720 100.120 ;
        RECT 282.200 99.950 282.440 100.350 ;
        RECT 281.160 99.500 281.565 99.670 ;
        RECT 281.900 99.580 282.440 99.950 ;
        RECT 282.610 100.165 282.930 100.520 ;
        RECT 283.175 100.440 283.480 100.900 ;
        RECT 283.650 100.190 283.905 100.720 ;
        RECT 282.610 99.990 282.935 100.165 ;
        RECT 282.610 99.690 283.525 99.990 ;
        RECT 282.785 99.660 283.525 99.690 ;
        RECT 280.260 99.330 280.935 99.490 ;
        RECT 281.395 99.410 281.565 99.500 ;
        RECT 280.260 99.320 281.225 99.330 ;
        RECT 279.900 99.150 280.070 99.290 ;
        RECT 276.645 98.350 276.895 98.810 ;
        RECT 277.065 98.520 277.315 98.850 ;
        RECT 277.530 98.520 278.210 98.850 ;
        RECT 278.380 98.950 279.455 99.120 ;
        RECT 279.900 98.980 280.460 99.150 ;
        RECT 280.765 99.030 281.225 99.320 ;
        RECT 281.395 99.240 282.615 99.410 ;
        RECT 278.380 98.610 278.550 98.950 ;
        RECT 278.785 98.350 279.115 98.780 ;
        RECT 279.285 98.610 279.455 98.950 ;
        RECT 279.750 98.350 280.120 98.810 ;
        RECT 280.290 98.520 280.460 98.980 ;
        RECT 281.395 98.860 281.565 99.240 ;
        RECT 282.785 99.070 282.955 99.660 ;
        RECT 283.695 99.540 283.905 100.190 ;
        RECT 284.355 100.090 284.600 100.695 ;
        RECT 284.820 100.365 285.330 100.900 ;
        RECT 280.695 98.520 281.565 98.860 ;
        RECT 282.155 98.900 282.955 99.070 ;
        RECT 281.735 98.350 281.985 98.810 ;
        RECT 282.155 98.610 282.325 98.900 ;
        RECT 282.505 98.350 282.835 98.730 ;
        RECT 283.175 98.350 283.480 99.490 ;
        RECT 283.650 98.660 283.905 99.540 ;
        RECT 284.080 99.920 285.310 100.090 ;
        RECT 284.080 99.110 284.420 99.920 ;
        RECT 284.590 99.355 285.340 99.545 ;
        RECT 284.080 98.700 284.595 99.110 ;
        RECT 284.830 98.350 285.000 99.110 ;
        RECT 285.170 98.690 285.340 99.355 ;
        RECT 285.510 99.370 285.700 100.730 ;
        RECT 285.870 99.880 286.145 100.730 ;
        RECT 286.335 100.365 286.865 100.730 ;
        RECT 287.290 100.500 287.620 100.900 ;
        RECT 286.690 100.330 286.865 100.365 ;
        RECT 285.870 99.710 286.150 99.880 ;
        RECT 285.870 99.570 286.145 99.710 ;
        RECT 286.350 99.370 286.520 100.170 ;
        RECT 285.510 99.200 286.520 99.370 ;
        RECT 286.690 100.160 287.620 100.330 ;
        RECT 287.790 100.160 288.045 100.730 ;
        RECT 288.310 100.350 288.480 100.730 ;
        RECT 288.695 100.520 289.025 100.900 ;
        RECT 288.310 100.180 289.025 100.350 ;
        RECT 286.690 99.030 286.860 100.160 ;
        RECT 287.450 99.990 287.620 100.160 ;
        RECT 285.735 98.860 286.860 99.030 ;
        RECT 287.030 99.660 287.225 99.990 ;
        RECT 287.450 99.660 287.705 99.990 ;
        RECT 287.030 98.690 287.200 99.660 ;
        RECT 287.875 99.490 288.045 100.160 ;
        RECT 288.220 99.630 288.575 100.000 ;
        RECT 288.855 99.990 289.025 100.180 ;
        RECT 289.195 100.155 289.450 100.730 ;
        RECT 288.855 99.660 289.110 99.990 ;
        RECT 285.170 98.520 287.200 98.690 ;
        RECT 287.370 98.350 287.540 99.490 ;
        RECT 287.710 98.520 288.045 99.490 ;
        RECT 288.855 99.450 289.025 99.660 ;
        RECT 288.310 99.280 289.025 99.450 ;
        RECT 289.280 99.425 289.450 100.155 ;
        RECT 289.625 100.060 289.885 100.900 ;
        RECT 290.980 100.175 291.270 100.900 ;
        RECT 291.530 100.350 291.700 100.730 ;
        RECT 291.915 100.520 292.245 100.900 ;
        RECT 291.530 100.180 292.245 100.350 ;
        RECT 291.440 99.630 291.795 100.000 ;
        RECT 292.075 99.990 292.245 100.180 ;
        RECT 292.415 100.155 292.670 100.730 ;
        RECT 292.075 99.660 292.330 99.990 ;
        RECT 288.310 98.520 288.480 99.280 ;
        RECT 288.695 98.350 289.025 99.110 ;
        RECT 289.195 98.520 289.450 99.425 ;
        RECT 289.625 98.350 289.885 99.500 ;
        RECT 290.980 98.350 291.270 99.515 ;
        RECT 292.075 99.450 292.245 99.660 ;
        RECT 291.530 99.280 292.245 99.450 ;
        RECT 292.500 99.425 292.670 100.155 ;
        RECT 292.845 100.060 293.105 100.900 ;
        RECT 293.745 100.350 294.000 100.640 ;
        RECT 294.170 100.520 294.500 100.900 ;
        RECT 293.745 100.180 294.495 100.350 ;
        RECT 291.530 98.520 291.700 99.280 ;
        RECT 291.915 98.350 292.245 99.110 ;
        RECT 292.415 98.520 292.670 99.425 ;
        RECT 292.845 98.350 293.105 99.500 ;
        RECT 293.745 99.360 294.095 100.010 ;
        RECT 294.265 99.190 294.495 100.180 ;
        RECT 293.745 99.020 294.495 99.190 ;
        RECT 293.745 98.520 294.000 99.020 ;
        RECT 294.170 98.350 294.500 98.850 ;
        RECT 294.670 98.520 294.840 100.640 ;
        RECT 295.200 100.540 295.530 100.900 ;
        RECT 295.700 100.510 296.195 100.680 ;
        RECT 296.400 100.510 297.255 100.680 ;
        RECT 295.070 99.320 295.530 100.370 ;
        RECT 295.010 98.535 295.335 99.320 ;
        RECT 295.700 99.150 295.870 100.510 ;
        RECT 296.040 99.600 296.390 100.220 ;
        RECT 296.560 100.000 296.915 100.220 ;
        RECT 296.560 99.410 296.730 100.000 ;
        RECT 297.085 99.800 297.255 100.510 ;
        RECT 298.130 100.440 298.460 100.900 ;
        RECT 298.670 100.540 299.020 100.710 ;
        RECT 297.460 99.970 298.250 100.220 ;
        RECT 298.670 100.150 298.930 100.540 ;
        RECT 299.240 100.450 300.190 100.730 ;
        RECT 300.360 100.460 300.550 100.900 ;
        RECT 300.720 100.520 301.790 100.690 ;
        RECT 298.420 99.800 298.590 99.980 ;
        RECT 295.700 98.980 296.095 99.150 ;
        RECT 296.265 99.020 296.730 99.410 ;
        RECT 296.900 99.630 298.590 99.800 ;
        RECT 295.925 98.850 296.095 98.980 ;
        RECT 296.900 98.850 297.070 99.630 ;
        RECT 298.760 99.460 298.930 100.150 ;
        RECT 297.430 99.290 298.930 99.460 ;
        RECT 299.120 99.490 299.330 100.280 ;
        RECT 299.500 99.660 299.850 100.280 ;
        RECT 300.020 99.670 300.190 100.450 ;
        RECT 300.720 100.290 300.890 100.520 ;
        RECT 300.360 100.120 300.890 100.290 ;
        RECT 300.360 99.840 300.580 100.120 ;
        RECT 301.060 99.950 301.300 100.350 ;
        RECT 300.020 99.500 300.425 99.670 ;
        RECT 300.760 99.580 301.300 99.950 ;
        RECT 301.470 100.165 301.790 100.520 ;
        RECT 302.035 100.440 302.340 100.900 ;
        RECT 302.510 100.190 302.765 100.720 ;
        RECT 301.470 99.990 301.795 100.165 ;
        RECT 301.470 99.690 302.385 99.990 ;
        RECT 301.645 99.660 302.385 99.690 ;
        RECT 299.120 99.330 299.795 99.490 ;
        RECT 300.255 99.410 300.425 99.500 ;
        RECT 299.120 99.320 300.085 99.330 ;
        RECT 298.760 99.150 298.930 99.290 ;
        RECT 295.505 98.350 295.755 98.810 ;
        RECT 295.925 98.520 296.175 98.850 ;
        RECT 296.390 98.520 297.070 98.850 ;
        RECT 297.240 98.950 298.315 99.120 ;
        RECT 298.760 98.980 299.320 99.150 ;
        RECT 299.625 99.030 300.085 99.320 ;
        RECT 300.255 99.240 301.475 99.410 ;
        RECT 297.240 98.610 297.410 98.950 ;
        RECT 297.645 98.350 297.975 98.780 ;
        RECT 298.145 98.610 298.315 98.950 ;
        RECT 298.610 98.350 298.980 98.810 ;
        RECT 299.150 98.520 299.320 98.980 ;
        RECT 300.255 98.860 300.425 99.240 ;
        RECT 301.645 99.070 301.815 99.660 ;
        RECT 302.555 99.540 302.765 100.190 ;
        RECT 302.945 100.060 303.205 100.900 ;
        RECT 303.380 100.155 303.635 100.730 ;
        RECT 303.805 100.520 304.135 100.900 ;
        RECT 304.350 100.350 304.520 100.730 ;
        RECT 303.805 100.180 304.520 100.350 ;
        RECT 304.870 100.350 305.040 100.730 ;
        RECT 305.255 100.520 305.585 100.900 ;
        RECT 304.870 100.180 305.585 100.350 ;
        RECT 299.555 98.520 300.425 98.860 ;
        RECT 301.015 98.900 301.815 99.070 ;
        RECT 300.595 98.350 300.845 98.810 ;
        RECT 301.015 98.610 301.185 98.900 ;
        RECT 301.365 98.350 301.695 98.730 ;
        RECT 302.035 98.350 302.340 99.490 ;
        RECT 302.510 98.660 302.765 99.540 ;
        RECT 302.945 98.350 303.205 99.500 ;
        RECT 303.380 99.425 303.550 100.155 ;
        RECT 303.805 99.990 303.975 100.180 ;
        RECT 303.720 99.660 303.975 99.990 ;
        RECT 303.805 99.450 303.975 99.660 ;
        RECT 304.255 99.630 304.610 100.000 ;
        RECT 304.780 99.630 305.135 100.000 ;
        RECT 305.415 99.990 305.585 100.180 ;
        RECT 305.755 100.155 306.010 100.730 ;
        RECT 305.415 99.660 305.670 99.990 ;
        RECT 305.415 99.450 305.585 99.660 ;
        RECT 303.380 98.520 303.635 99.425 ;
        RECT 303.805 99.280 304.520 99.450 ;
        RECT 303.805 98.350 304.135 99.110 ;
        RECT 304.350 98.520 304.520 99.280 ;
        RECT 304.870 99.280 305.585 99.450 ;
        RECT 305.840 99.425 306.010 100.155 ;
        RECT 306.185 100.060 306.445 100.900 ;
        RECT 307.170 100.350 307.340 100.730 ;
        RECT 307.555 100.520 307.885 100.900 ;
        RECT 307.170 100.180 307.885 100.350 ;
        RECT 307.080 99.630 307.435 100.000 ;
        RECT 307.715 99.990 307.885 100.180 ;
        RECT 308.055 100.155 308.310 100.730 ;
        RECT 307.715 99.660 307.970 99.990 ;
        RECT 304.870 98.520 305.040 99.280 ;
        RECT 305.255 98.350 305.585 99.110 ;
        RECT 305.755 98.520 306.010 99.425 ;
        RECT 306.185 98.350 306.445 99.500 ;
        RECT 307.715 99.450 307.885 99.660 ;
        RECT 307.170 99.280 307.885 99.450 ;
        RECT 308.140 99.425 308.310 100.155 ;
        RECT 308.485 100.060 308.745 100.900 ;
        RECT 309.840 100.150 311.050 100.900 ;
        RECT 307.170 98.520 307.340 99.280 ;
        RECT 307.555 98.350 307.885 99.110 ;
        RECT 308.055 98.520 308.310 99.425 ;
        RECT 308.485 98.350 308.745 99.500 ;
        RECT 309.840 99.440 310.360 99.980 ;
        RECT 310.530 99.610 311.050 100.150 ;
        RECT 309.840 98.350 311.050 99.440 ;
        RECT 162.095 98.180 311.135 98.350 ;
        RECT 162.180 97.090 163.390 98.180 ;
        RECT 162.180 96.380 162.700 96.920 ;
        RECT 162.870 96.550 163.390 97.090 ;
        RECT 163.565 97.030 163.825 98.180 ;
        RECT 164.000 97.105 164.255 98.010 ;
        RECT 164.425 97.420 164.755 98.180 ;
        RECT 164.970 97.250 165.140 98.010 ;
        RECT 165.865 97.510 166.120 98.010 ;
        RECT 166.290 97.680 166.620 98.180 ;
        RECT 165.865 97.340 166.615 97.510 ;
        RECT 162.180 95.630 163.390 96.380 ;
        RECT 163.565 95.630 163.825 96.470 ;
        RECT 164.000 96.375 164.170 97.105 ;
        RECT 164.425 97.080 165.140 97.250 ;
        RECT 164.425 96.870 164.595 97.080 ;
        RECT 164.340 96.540 164.595 96.870 ;
        RECT 164.000 95.800 164.255 96.375 ;
        RECT 164.425 96.350 164.595 96.540 ;
        RECT 164.875 96.530 165.230 96.900 ;
        RECT 165.865 96.520 166.215 97.170 ;
        RECT 166.385 96.350 166.615 97.340 ;
        RECT 164.425 96.180 165.140 96.350 ;
        RECT 164.425 95.630 164.755 96.010 ;
        RECT 164.970 95.800 165.140 96.180 ;
        RECT 165.865 96.180 166.615 96.350 ;
        RECT 165.865 95.890 166.120 96.180 ;
        RECT 166.290 95.630 166.620 96.010 ;
        RECT 166.790 95.890 166.960 98.010 ;
        RECT 167.130 97.210 167.455 97.995 ;
        RECT 167.625 97.720 167.875 98.180 ;
        RECT 168.045 97.680 168.295 98.010 ;
        RECT 168.510 97.680 169.190 98.010 ;
        RECT 168.045 97.550 168.215 97.680 ;
        RECT 167.820 97.380 168.215 97.550 ;
        RECT 167.190 96.160 167.650 97.210 ;
        RECT 167.820 96.020 167.990 97.380 ;
        RECT 168.385 97.120 168.850 97.510 ;
        RECT 168.160 96.310 168.510 96.930 ;
        RECT 168.680 96.530 168.850 97.120 ;
        RECT 169.020 96.900 169.190 97.680 ;
        RECT 169.360 97.580 169.530 97.920 ;
        RECT 169.765 97.750 170.095 98.180 ;
        RECT 170.265 97.580 170.435 97.920 ;
        RECT 170.730 97.720 171.100 98.180 ;
        RECT 169.360 97.410 170.435 97.580 ;
        RECT 171.270 97.550 171.440 98.010 ;
        RECT 171.675 97.670 172.545 98.010 ;
        RECT 172.715 97.720 172.965 98.180 ;
        RECT 170.880 97.380 171.440 97.550 ;
        RECT 170.880 97.240 171.050 97.380 ;
        RECT 169.550 97.070 171.050 97.240 ;
        RECT 171.745 97.210 172.205 97.500 ;
        RECT 169.020 96.730 170.710 96.900 ;
        RECT 168.680 96.310 169.035 96.530 ;
        RECT 169.205 96.020 169.375 96.730 ;
        RECT 169.580 96.310 170.370 96.560 ;
        RECT 170.540 96.550 170.710 96.730 ;
        RECT 170.880 96.380 171.050 97.070 ;
        RECT 167.320 95.630 167.650 95.990 ;
        RECT 167.820 95.850 168.315 96.020 ;
        RECT 168.520 95.850 169.375 96.020 ;
        RECT 170.250 95.630 170.580 96.090 ;
        RECT 170.790 95.990 171.050 96.380 ;
        RECT 171.240 97.200 172.205 97.210 ;
        RECT 172.375 97.290 172.545 97.670 ;
        RECT 173.135 97.630 173.305 97.920 ;
        RECT 173.485 97.800 173.815 98.180 ;
        RECT 173.135 97.460 173.935 97.630 ;
        RECT 171.240 97.040 171.915 97.200 ;
        RECT 172.375 97.120 173.595 97.290 ;
        RECT 171.240 96.250 171.450 97.040 ;
        RECT 172.375 97.030 172.545 97.120 ;
        RECT 171.620 96.250 171.970 96.870 ;
        RECT 172.140 96.860 172.545 97.030 ;
        RECT 172.140 96.080 172.310 96.860 ;
        RECT 172.480 96.410 172.700 96.690 ;
        RECT 172.880 96.580 173.420 96.950 ;
        RECT 173.765 96.870 173.935 97.460 ;
        RECT 174.155 97.040 174.460 98.180 ;
        RECT 174.630 96.990 174.885 97.870 ;
        RECT 175.060 97.015 175.350 98.180 ;
        RECT 175.525 97.040 175.860 98.010 ;
        RECT 176.030 97.040 176.200 98.180 ;
        RECT 176.370 97.840 178.400 98.010 ;
        RECT 173.765 96.840 174.505 96.870 ;
        RECT 172.480 96.240 173.010 96.410 ;
        RECT 170.790 95.820 171.140 95.990 ;
        RECT 171.360 95.800 172.310 96.080 ;
        RECT 172.480 95.630 172.670 96.070 ;
        RECT 172.840 96.010 173.010 96.240 ;
        RECT 173.180 96.180 173.420 96.580 ;
        RECT 173.590 96.540 174.505 96.840 ;
        RECT 173.590 96.365 173.915 96.540 ;
        RECT 173.590 96.010 173.910 96.365 ;
        RECT 174.675 96.340 174.885 96.990 ;
        RECT 175.525 96.370 175.695 97.040 ;
        RECT 176.370 96.870 176.540 97.840 ;
        RECT 175.865 96.540 176.120 96.870 ;
        RECT 176.345 96.540 176.540 96.870 ;
        RECT 176.710 97.500 177.835 97.670 ;
        RECT 175.950 96.370 176.120 96.540 ;
        RECT 176.710 96.370 176.880 97.500 ;
        RECT 172.840 95.840 173.910 96.010 ;
        RECT 174.155 95.630 174.460 96.090 ;
        RECT 174.630 95.810 174.885 96.340 ;
        RECT 175.060 95.630 175.350 96.355 ;
        RECT 175.525 95.800 175.780 96.370 ;
        RECT 175.950 96.200 176.880 96.370 ;
        RECT 177.050 97.160 178.060 97.330 ;
        RECT 177.050 96.360 177.220 97.160 ;
        RECT 176.705 96.165 176.880 96.200 ;
        RECT 175.950 95.630 176.280 96.030 ;
        RECT 176.705 95.800 177.235 96.165 ;
        RECT 177.425 96.140 177.700 96.960 ;
        RECT 177.420 95.970 177.700 96.140 ;
        RECT 177.425 95.800 177.700 95.970 ;
        RECT 177.870 95.800 178.060 97.160 ;
        RECT 178.230 97.175 178.400 97.840 ;
        RECT 178.570 97.420 178.740 98.180 ;
        RECT 178.975 97.420 179.490 97.830 ;
        RECT 178.230 96.985 178.980 97.175 ;
        RECT 179.150 96.610 179.490 97.420 ;
        RECT 179.660 97.090 181.330 98.180 ;
        RECT 178.260 96.440 179.490 96.610 ;
        RECT 178.240 95.630 178.750 96.165 ;
        RECT 178.970 95.835 179.215 96.440 ;
        RECT 179.660 96.400 180.410 96.920 ;
        RECT 180.580 96.570 181.330 97.090 ;
        RECT 181.500 96.575 181.780 98.010 ;
        RECT 181.950 97.405 182.660 98.180 ;
        RECT 182.830 97.235 183.160 98.010 ;
        RECT 182.010 97.020 183.160 97.235 ;
        RECT 179.660 95.630 181.330 96.400 ;
        RECT 181.500 95.800 181.840 96.575 ;
        RECT 182.010 96.450 182.295 97.020 ;
        RECT 182.480 96.620 182.950 96.850 ;
        RECT 183.355 96.820 183.570 97.935 ;
        RECT 183.750 97.460 184.080 98.180 ;
        RECT 184.265 97.510 184.520 98.010 ;
        RECT 184.690 97.680 185.020 98.180 ;
        RECT 184.265 97.340 185.015 97.510 ;
        RECT 183.860 96.820 184.090 97.160 ;
        RECT 183.120 96.640 183.570 96.820 ;
        RECT 183.120 96.620 183.450 96.640 ;
        RECT 183.760 96.620 184.090 96.820 ;
        RECT 184.265 96.520 184.615 97.170 ;
        RECT 182.010 96.260 182.720 96.450 ;
        RECT 182.420 96.120 182.720 96.260 ;
        RECT 182.910 96.260 184.090 96.450 ;
        RECT 184.785 96.350 185.015 97.340 ;
        RECT 182.910 96.180 183.240 96.260 ;
        RECT 182.420 96.110 182.735 96.120 ;
        RECT 182.420 96.100 182.745 96.110 ;
        RECT 182.420 96.095 182.755 96.100 ;
        RECT 182.010 95.630 182.180 96.090 ;
        RECT 182.420 96.085 182.760 96.095 ;
        RECT 182.420 96.080 182.765 96.085 ;
        RECT 182.420 96.070 182.770 96.080 ;
        RECT 182.420 96.065 182.775 96.070 ;
        RECT 182.420 95.800 182.780 96.065 ;
        RECT 183.410 95.630 183.580 96.090 ;
        RECT 183.750 95.800 184.090 96.260 ;
        RECT 184.265 96.180 185.015 96.350 ;
        RECT 184.265 95.890 184.520 96.180 ;
        RECT 184.690 95.630 185.020 96.010 ;
        RECT 185.190 95.890 185.360 98.010 ;
        RECT 185.530 97.210 185.855 97.995 ;
        RECT 186.025 97.720 186.275 98.180 ;
        RECT 186.445 97.680 186.695 98.010 ;
        RECT 186.910 97.680 187.590 98.010 ;
        RECT 186.445 97.550 186.615 97.680 ;
        RECT 186.220 97.380 186.615 97.550 ;
        RECT 185.590 96.160 186.050 97.210 ;
        RECT 186.220 96.020 186.390 97.380 ;
        RECT 186.785 97.120 187.250 97.510 ;
        RECT 186.560 96.310 186.910 96.930 ;
        RECT 187.080 96.530 187.250 97.120 ;
        RECT 187.420 96.900 187.590 97.680 ;
        RECT 187.760 97.580 187.930 97.920 ;
        RECT 188.165 97.750 188.495 98.180 ;
        RECT 188.665 97.580 188.835 97.920 ;
        RECT 189.130 97.720 189.500 98.180 ;
        RECT 187.760 97.410 188.835 97.580 ;
        RECT 189.670 97.550 189.840 98.010 ;
        RECT 190.075 97.670 190.945 98.010 ;
        RECT 191.115 97.720 191.365 98.180 ;
        RECT 189.280 97.380 189.840 97.550 ;
        RECT 189.280 97.240 189.450 97.380 ;
        RECT 187.950 97.070 189.450 97.240 ;
        RECT 190.145 97.210 190.605 97.500 ;
        RECT 187.420 96.730 189.110 96.900 ;
        RECT 187.080 96.310 187.435 96.530 ;
        RECT 187.605 96.020 187.775 96.730 ;
        RECT 187.980 96.310 188.770 96.560 ;
        RECT 188.940 96.550 189.110 96.730 ;
        RECT 189.280 96.380 189.450 97.070 ;
        RECT 185.720 95.630 186.050 95.990 ;
        RECT 186.220 95.850 186.715 96.020 ;
        RECT 186.920 95.850 187.775 96.020 ;
        RECT 188.650 95.630 188.980 96.090 ;
        RECT 189.190 95.990 189.450 96.380 ;
        RECT 189.640 97.200 190.605 97.210 ;
        RECT 190.775 97.290 190.945 97.670 ;
        RECT 191.535 97.630 191.705 97.920 ;
        RECT 191.885 97.800 192.215 98.180 ;
        RECT 191.535 97.460 192.335 97.630 ;
        RECT 189.640 97.040 190.315 97.200 ;
        RECT 190.775 97.120 191.995 97.290 ;
        RECT 189.640 96.250 189.850 97.040 ;
        RECT 190.775 97.030 190.945 97.120 ;
        RECT 190.020 96.250 190.370 96.870 ;
        RECT 190.540 96.860 190.945 97.030 ;
        RECT 190.540 96.080 190.710 96.860 ;
        RECT 190.880 96.410 191.100 96.690 ;
        RECT 191.280 96.580 191.820 96.950 ;
        RECT 192.165 96.870 192.335 97.460 ;
        RECT 192.555 97.040 192.860 98.180 ;
        RECT 193.030 96.990 193.285 97.870 ;
        RECT 192.165 96.840 192.905 96.870 ;
        RECT 190.880 96.240 191.410 96.410 ;
        RECT 189.190 95.820 189.540 95.990 ;
        RECT 189.760 95.800 190.710 96.080 ;
        RECT 190.880 95.630 191.070 96.070 ;
        RECT 191.240 96.010 191.410 96.240 ;
        RECT 191.580 96.180 191.820 96.580 ;
        RECT 191.990 96.540 192.905 96.840 ;
        RECT 191.990 96.365 192.315 96.540 ;
        RECT 191.990 96.010 192.310 96.365 ;
        RECT 193.075 96.340 193.285 96.990 ;
        RECT 191.240 95.840 192.310 96.010 ;
        RECT 192.555 95.630 192.860 96.090 ;
        RECT 193.030 95.810 193.285 96.340 ;
        RECT 193.465 97.040 193.800 98.010 ;
        RECT 193.970 97.040 194.140 98.180 ;
        RECT 194.310 97.840 196.340 98.010 ;
        RECT 193.465 96.370 193.635 97.040 ;
        RECT 194.310 96.870 194.480 97.840 ;
        RECT 193.805 96.540 194.060 96.870 ;
        RECT 194.285 96.540 194.480 96.870 ;
        RECT 194.650 97.500 195.775 97.670 ;
        RECT 193.890 96.370 194.060 96.540 ;
        RECT 194.650 96.370 194.820 97.500 ;
        RECT 193.465 95.800 193.720 96.370 ;
        RECT 193.890 96.200 194.820 96.370 ;
        RECT 194.990 97.160 196.000 97.330 ;
        RECT 194.990 96.360 195.160 97.160 ;
        RECT 194.645 96.165 194.820 96.200 ;
        RECT 193.890 95.630 194.220 96.030 ;
        RECT 194.645 95.800 195.175 96.165 ;
        RECT 195.365 96.140 195.640 96.960 ;
        RECT 195.360 95.970 195.640 96.140 ;
        RECT 195.365 95.800 195.640 95.970 ;
        RECT 195.810 95.800 196.000 97.160 ;
        RECT 196.170 97.175 196.340 97.840 ;
        RECT 196.510 97.420 196.680 98.180 ;
        RECT 196.915 97.420 197.430 97.830 ;
        RECT 196.170 96.985 196.920 97.175 ;
        RECT 197.090 96.610 197.430 97.420 ;
        RECT 197.655 97.310 197.940 98.180 ;
        RECT 198.110 97.550 198.370 98.010 ;
        RECT 198.545 97.720 198.800 98.180 ;
        RECT 198.970 97.550 199.230 98.010 ;
        RECT 198.110 97.380 199.230 97.550 ;
        RECT 199.400 97.380 199.710 98.180 ;
        RECT 198.110 97.130 198.370 97.380 ;
        RECT 199.880 97.210 200.190 98.010 ;
        RECT 196.200 96.440 197.430 96.610 ;
        RECT 197.615 96.960 198.370 97.130 ;
        RECT 199.160 97.040 200.190 97.210 ;
        RECT 197.615 96.450 198.020 96.960 ;
        RECT 199.160 96.790 199.330 97.040 ;
        RECT 198.190 96.620 199.330 96.790 ;
        RECT 196.180 95.630 196.690 96.165 ;
        RECT 196.910 95.835 197.155 96.440 ;
        RECT 197.615 96.280 199.265 96.450 ;
        RECT 199.500 96.300 199.850 96.870 ;
        RECT 197.660 95.630 197.940 96.110 ;
        RECT 198.110 95.890 198.370 96.280 ;
        RECT 198.545 95.630 198.800 96.110 ;
        RECT 198.970 95.890 199.265 96.280 ;
        RECT 200.020 96.130 200.190 97.040 ;
        RECT 200.820 97.015 201.110 98.180 ;
        RECT 201.280 97.090 202.490 98.180 ;
        RECT 201.280 96.380 201.800 96.920 ;
        RECT 201.970 96.550 202.490 97.090 ;
        RECT 199.445 95.630 199.720 96.110 ;
        RECT 199.890 95.800 200.190 96.130 ;
        RECT 200.820 95.630 201.110 96.355 ;
        RECT 201.280 95.630 202.490 96.380 ;
        RECT 202.670 95.810 202.930 98.000 ;
        RECT 203.100 97.450 203.440 98.180 ;
        RECT 203.620 97.270 203.890 98.000 ;
        RECT 203.120 97.050 203.890 97.270 ;
        RECT 204.070 97.290 204.300 98.000 ;
        RECT 204.470 97.470 204.800 98.180 ;
        RECT 204.970 97.290 205.230 98.000 ;
        RECT 204.070 97.050 205.230 97.290 ;
        RECT 205.420 97.330 205.680 98.010 ;
        RECT 205.850 97.400 206.100 98.180 ;
        RECT 206.350 97.630 206.600 98.010 ;
        RECT 206.770 97.800 207.125 98.180 ;
        RECT 208.130 97.790 208.465 98.010 ;
        RECT 207.730 97.630 207.960 97.670 ;
        RECT 206.350 97.430 207.960 97.630 ;
        RECT 206.350 97.420 207.185 97.430 ;
        RECT 207.775 97.340 207.960 97.430 ;
        RECT 203.120 96.380 203.410 97.050 ;
        RECT 203.590 96.560 204.055 96.870 ;
        RECT 204.235 96.560 204.760 96.870 ;
        RECT 203.120 96.180 204.350 96.380 ;
        RECT 203.190 95.630 203.860 96.000 ;
        RECT 204.040 95.810 204.350 96.180 ;
        RECT 204.530 95.920 204.760 96.560 ;
        RECT 204.940 96.540 205.240 96.870 ;
        RECT 204.940 95.630 205.230 96.360 ;
        RECT 205.420 96.140 205.590 97.330 ;
        RECT 207.290 97.230 207.620 97.260 ;
        RECT 205.820 97.170 207.620 97.230 ;
        RECT 208.210 97.170 208.465 97.790 ;
        RECT 208.755 97.550 209.040 98.010 ;
        RECT 209.210 97.720 209.480 98.180 ;
        RECT 208.755 97.330 209.710 97.550 ;
        RECT 205.760 97.060 208.465 97.170 ;
        RECT 205.760 97.025 205.960 97.060 ;
        RECT 205.760 96.450 205.930 97.025 ;
        RECT 207.290 97.000 208.465 97.060 ;
        RECT 206.160 96.585 206.570 96.890 ;
        RECT 206.740 96.620 207.070 96.830 ;
        RECT 205.760 96.330 206.030 96.450 ;
        RECT 205.760 96.285 206.605 96.330 ;
        RECT 205.850 96.160 206.605 96.285 ;
        RECT 206.860 96.220 207.070 96.620 ;
        RECT 207.315 96.620 207.790 96.830 ;
        RECT 207.980 96.620 208.470 96.820 ;
        RECT 207.315 96.220 207.535 96.620 ;
        RECT 208.640 96.600 209.330 97.160 ;
        RECT 209.500 96.430 209.710 97.330 ;
        RECT 205.420 96.130 205.650 96.140 ;
        RECT 205.420 95.800 205.680 96.130 ;
        RECT 206.435 96.010 206.605 96.160 ;
        RECT 205.850 95.630 206.180 95.990 ;
        RECT 206.435 95.800 207.735 96.010 ;
        RECT 208.010 95.630 208.465 96.395 ;
        RECT 208.755 96.260 209.710 96.430 ;
        RECT 209.880 97.160 210.280 98.010 ;
        RECT 210.470 97.550 210.750 98.010 ;
        RECT 211.270 97.720 211.595 98.180 ;
        RECT 210.470 97.330 211.595 97.550 ;
        RECT 209.880 96.600 210.975 97.160 ;
        RECT 211.145 96.870 211.595 97.330 ;
        RECT 211.765 97.040 212.150 98.010 ;
        RECT 212.320 97.745 217.665 98.180 ;
        RECT 208.755 95.800 209.040 96.260 ;
        RECT 209.210 95.630 209.480 96.090 ;
        RECT 209.880 95.800 210.280 96.600 ;
        RECT 211.145 96.540 211.700 96.870 ;
        RECT 211.145 96.430 211.595 96.540 ;
        RECT 210.470 96.260 211.595 96.430 ;
        RECT 211.870 96.370 212.150 97.040 ;
        RECT 210.470 95.800 210.750 96.260 ;
        RECT 211.270 95.630 211.595 96.090 ;
        RECT 211.765 95.800 212.150 96.370 ;
        RECT 213.905 96.175 214.245 97.005 ;
        RECT 215.725 96.495 216.075 97.745 ;
        RECT 217.840 97.090 220.430 98.180 ;
        RECT 217.840 96.400 219.050 96.920 ;
        RECT 219.220 96.570 220.430 97.090 ;
        RECT 220.600 96.575 220.880 98.010 ;
        RECT 221.050 97.405 221.760 98.180 ;
        RECT 221.930 97.235 222.260 98.010 ;
        RECT 221.110 97.020 222.260 97.235 ;
        RECT 212.320 95.630 217.665 96.175 ;
        RECT 217.840 95.630 220.430 96.400 ;
        RECT 220.600 95.800 220.940 96.575 ;
        RECT 221.110 96.450 221.395 97.020 ;
        RECT 221.580 96.620 222.050 96.850 ;
        RECT 222.455 96.820 222.670 97.935 ;
        RECT 222.850 97.460 223.180 98.180 ;
        RECT 223.365 97.790 223.700 98.010 ;
        RECT 224.705 97.800 225.060 98.180 ;
        RECT 223.365 97.170 223.620 97.790 ;
        RECT 223.870 97.630 224.100 97.670 ;
        RECT 225.230 97.630 225.480 98.010 ;
        RECT 223.870 97.430 225.480 97.630 ;
        RECT 223.870 97.340 224.055 97.430 ;
        RECT 224.645 97.420 225.480 97.430 ;
        RECT 225.730 97.400 225.980 98.180 ;
        RECT 226.150 97.330 226.410 98.010 ;
        RECT 224.210 97.230 224.540 97.260 ;
        RECT 224.210 97.170 226.010 97.230 ;
        RECT 222.960 96.820 223.190 97.160 ;
        RECT 223.365 97.060 226.070 97.170 ;
        RECT 223.365 97.000 224.540 97.060 ;
        RECT 225.870 97.025 226.070 97.060 ;
        RECT 222.220 96.640 222.670 96.820 ;
        RECT 222.220 96.620 222.550 96.640 ;
        RECT 222.860 96.620 223.190 96.820 ;
        RECT 223.360 96.620 223.850 96.820 ;
        RECT 224.040 96.620 224.515 96.830 ;
        RECT 221.110 96.260 221.820 96.450 ;
        RECT 221.520 96.120 221.820 96.260 ;
        RECT 222.010 96.260 223.190 96.450 ;
        RECT 222.010 96.180 222.340 96.260 ;
        RECT 221.520 96.110 221.835 96.120 ;
        RECT 221.520 96.100 221.845 96.110 ;
        RECT 221.520 96.095 221.855 96.100 ;
        RECT 221.110 95.630 221.280 96.090 ;
        RECT 221.520 96.085 221.860 96.095 ;
        RECT 221.520 96.080 221.865 96.085 ;
        RECT 221.520 96.070 221.870 96.080 ;
        RECT 221.520 96.065 221.875 96.070 ;
        RECT 221.520 95.800 221.880 96.065 ;
        RECT 222.510 95.630 222.680 96.090 ;
        RECT 222.850 95.800 223.190 96.260 ;
        RECT 223.365 95.630 223.820 96.395 ;
        RECT 224.295 96.220 224.515 96.620 ;
        RECT 224.760 96.620 225.090 96.830 ;
        RECT 224.760 96.220 224.970 96.620 ;
        RECT 225.260 96.585 225.670 96.890 ;
        RECT 225.900 96.450 226.070 97.025 ;
        RECT 225.800 96.330 226.070 96.450 ;
        RECT 225.225 96.285 226.070 96.330 ;
        RECT 225.225 96.160 225.980 96.285 ;
        RECT 225.225 96.010 225.395 96.160 ;
        RECT 226.240 96.130 226.410 97.330 ;
        RECT 226.580 97.015 226.870 98.180 ;
        RECT 227.060 97.340 227.315 98.010 ;
        RECT 227.485 97.420 227.815 98.180 ;
        RECT 227.985 97.580 228.235 98.010 ;
        RECT 228.405 97.760 228.760 98.180 ;
        RECT 228.950 97.840 230.120 98.010 ;
        RECT 228.950 97.800 229.280 97.840 ;
        RECT 229.390 97.580 229.620 97.670 ;
        RECT 227.985 97.340 229.620 97.580 ;
        RECT 229.790 97.340 230.120 97.840 ;
        RECT 224.095 95.800 225.395 96.010 ;
        RECT 225.650 95.630 225.980 95.990 ;
        RECT 226.150 95.800 226.410 96.130 ;
        RECT 226.580 95.630 226.870 96.355 ;
        RECT 227.060 96.210 227.230 97.340 ;
        RECT 230.290 97.170 230.460 98.010 ;
        RECT 230.720 97.745 236.065 98.180 ;
        RECT 236.240 97.745 241.585 98.180 ;
        RECT 227.400 97.000 230.460 97.170 ;
        RECT 227.400 96.450 227.570 97.000 ;
        RECT 227.790 96.650 228.165 96.820 ;
        RECT 227.800 96.620 228.165 96.650 ;
        RECT 228.335 96.620 228.665 96.820 ;
        RECT 227.400 96.280 228.200 96.450 ;
        RECT 227.060 96.140 227.245 96.210 ;
        RECT 227.060 96.130 227.270 96.140 ;
        RECT 227.060 95.800 227.315 96.130 ;
        RECT 227.530 95.630 227.860 96.110 ;
        RECT 228.030 96.050 228.200 96.280 ;
        RECT 228.380 96.220 228.665 96.620 ;
        RECT 228.935 96.620 229.410 96.820 ;
        RECT 229.580 96.620 230.025 96.820 ;
        RECT 230.195 96.620 230.545 96.830 ;
        RECT 228.935 96.220 229.215 96.620 ;
        RECT 229.395 96.280 230.460 96.450 ;
        RECT 229.395 96.050 229.565 96.280 ;
        RECT 228.030 95.800 229.565 96.050 ;
        RECT 229.790 95.630 230.120 96.110 ;
        RECT 230.290 95.800 230.460 96.280 ;
        RECT 232.305 96.175 232.645 97.005 ;
        RECT 234.125 96.495 234.475 97.745 ;
        RECT 237.825 96.175 238.165 97.005 ;
        RECT 239.645 96.495 239.995 97.745 ;
        RECT 241.760 97.090 242.970 98.180 ;
        RECT 241.760 96.380 242.280 96.920 ;
        RECT 242.450 96.550 242.970 97.090 ;
        RECT 243.140 97.330 243.400 98.010 ;
        RECT 243.570 97.400 243.820 98.180 ;
        RECT 244.070 97.630 244.320 98.010 ;
        RECT 244.490 97.800 244.845 98.180 ;
        RECT 245.850 97.790 246.185 98.010 ;
        RECT 245.450 97.630 245.680 97.670 ;
        RECT 244.070 97.430 245.680 97.630 ;
        RECT 244.070 97.420 244.905 97.430 ;
        RECT 245.495 97.340 245.680 97.430 ;
        RECT 230.720 95.630 236.065 96.175 ;
        RECT 236.240 95.630 241.585 96.175 ;
        RECT 241.760 95.630 242.970 96.380 ;
        RECT 243.140 96.130 243.310 97.330 ;
        RECT 245.010 97.230 245.340 97.260 ;
        RECT 243.540 97.170 245.340 97.230 ;
        RECT 245.930 97.170 246.185 97.790 ;
        RECT 243.480 97.060 246.185 97.170 ;
        RECT 243.480 97.025 243.680 97.060 ;
        RECT 243.480 96.450 243.650 97.025 ;
        RECT 245.010 97.000 246.185 97.060 ;
        RECT 246.450 97.170 246.620 98.010 ;
        RECT 246.790 97.840 247.960 98.010 ;
        RECT 246.790 97.340 247.120 97.840 ;
        RECT 247.630 97.800 247.960 97.840 ;
        RECT 248.150 97.760 248.505 98.180 ;
        RECT 247.290 97.580 247.520 97.670 ;
        RECT 248.675 97.580 248.925 98.010 ;
        RECT 247.290 97.340 248.925 97.580 ;
        RECT 249.095 97.420 249.425 98.180 ;
        RECT 249.595 97.340 249.850 98.010 ;
        RECT 246.450 97.000 249.510 97.170 ;
        RECT 243.880 96.585 244.290 96.890 ;
        RECT 244.460 96.620 244.790 96.830 ;
        RECT 243.480 96.330 243.750 96.450 ;
        RECT 243.480 96.285 244.325 96.330 ;
        RECT 243.570 96.160 244.325 96.285 ;
        RECT 244.580 96.220 244.790 96.620 ;
        RECT 245.035 96.620 245.510 96.830 ;
        RECT 245.700 96.620 246.190 96.820 ;
        RECT 246.365 96.620 246.715 96.830 ;
        RECT 246.885 96.620 247.330 96.820 ;
        RECT 247.500 96.620 247.975 96.820 ;
        RECT 245.035 96.220 245.255 96.620 ;
        RECT 243.140 95.800 243.400 96.130 ;
        RECT 244.155 96.010 244.325 96.160 ;
        RECT 243.570 95.630 243.900 95.990 ;
        RECT 244.155 95.800 245.455 96.010 ;
        RECT 245.730 95.630 246.185 96.395 ;
        RECT 246.450 96.280 247.515 96.450 ;
        RECT 246.450 95.800 246.620 96.280 ;
        RECT 246.790 95.630 247.120 96.110 ;
        RECT 247.345 96.050 247.515 96.280 ;
        RECT 247.695 96.220 247.975 96.620 ;
        RECT 248.245 96.620 248.575 96.820 ;
        RECT 248.745 96.620 249.110 96.820 ;
        RECT 248.245 96.220 248.530 96.620 ;
        RECT 249.340 96.450 249.510 97.000 ;
        RECT 248.710 96.280 249.510 96.450 ;
        RECT 248.710 96.050 248.880 96.280 ;
        RECT 249.680 96.210 249.850 97.340 ;
        RECT 250.040 97.090 251.710 98.180 ;
        RECT 249.665 96.140 249.850 96.210 ;
        RECT 249.640 96.130 249.850 96.140 ;
        RECT 247.345 95.800 248.880 96.050 ;
        RECT 249.050 95.630 249.380 96.110 ;
        RECT 249.595 95.800 249.850 96.130 ;
        RECT 250.040 96.400 250.790 96.920 ;
        RECT 250.960 96.570 251.710 97.090 ;
        RECT 252.340 97.015 252.630 98.180 ;
        RECT 252.820 97.340 253.075 98.010 ;
        RECT 253.245 97.420 253.575 98.180 ;
        RECT 253.745 97.580 253.995 98.010 ;
        RECT 254.165 97.760 254.520 98.180 ;
        RECT 254.710 97.840 255.880 98.010 ;
        RECT 254.710 97.800 255.040 97.840 ;
        RECT 255.150 97.580 255.380 97.670 ;
        RECT 253.745 97.340 255.380 97.580 ;
        RECT 255.550 97.340 255.880 97.840 ;
        RECT 250.040 95.630 251.710 96.400 ;
        RECT 252.340 95.630 252.630 96.355 ;
        RECT 252.820 96.210 252.990 97.340 ;
        RECT 256.050 97.170 256.220 98.010 ;
        RECT 253.160 97.000 256.220 97.170 ;
        RECT 257.410 97.115 257.720 98.180 ;
        RECT 257.890 97.510 258.125 98.010 ;
        RECT 258.295 97.720 258.625 98.180 ;
        RECT 258.820 97.840 259.930 98.010 ;
        RECT 258.820 97.680 259.010 97.840 ;
        RECT 259.240 97.510 259.540 97.670 ;
        RECT 257.890 97.330 259.540 97.510 ;
        RECT 259.710 97.330 259.930 97.840 ;
        RECT 260.100 97.330 260.430 98.180 ;
        RECT 260.620 97.745 265.965 98.180 ;
        RECT 266.140 97.745 271.485 98.180 ;
        RECT 253.160 96.450 253.330 97.000 ;
        RECT 253.560 96.620 253.925 96.820 ;
        RECT 254.095 96.620 254.425 96.820 ;
        RECT 253.160 96.280 253.960 96.450 ;
        RECT 252.820 96.140 253.005 96.210 ;
        RECT 252.820 96.130 253.030 96.140 ;
        RECT 252.820 95.800 253.075 96.130 ;
        RECT 253.290 95.630 253.620 96.110 ;
        RECT 253.790 96.050 253.960 96.280 ;
        RECT 254.140 96.220 254.425 96.620 ;
        RECT 254.695 96.620 255.170 96.820 ;
        RECT 255.340 96.620 255.785 96.820 ;
        RECT 255.955 96.620 256.305 96.830 ;
        RECT 254.695 96.220 254.975 96.620 ;
        RECT 255.155 96.280 256.220 96.450 ;
        RECT 257.405 96.310 257.720 96.945 ;
        RECT 255.155 96.050 255.325 96.280 ;
        RECT 253.790 95.800 255.325 96.050 ;
        RECT 255.550 95.630 255.880 96.110 ;
        RECT 256.050 95.800 256.220 96.280 ;
        RECT 257.890 96.140 258.100 97.330 ;
        RECT 258.440 96.990 260.415 97.160 ;
        RECT 258.440 96.620 258.935 96.990 ;
        RECT 259.115 96.620 259.915 96.820 ;
        RECT 260.085 96.600 260.415 96.990 ;
        RECT 258.270 96.260 260.430 96.430 ;
        RECT 257.410 95.970 257.720 96.140 ;
        RECT 258.270 95.970 258.600 96.260 ;
        RECT 257.410 95.800 258.600 95.970 ;
        RECT 258.840 95.630 259.010 96.090 ;
        RECT 259.240 95.800 259.570 96.260 ;
        RECT 259.750 95.630 259.920 96.090 ;
        RECT 260.100 95.800 260.430 96.260 ;
        RECT 262.205 96.175 262.545 97.005 ;
        RECT 264.025 96.495 264.375 97.745 ;
        RECT 267.725 96.175 268.065 97.005 ;
        RECT 269.545 96.495 269.895 97.745 ;
        RECT 271.660 97.090 273.330 98.180 ;
        RECT 271.660 96.400 272.410 96.920 ;
        RECT 272.580 96.570 273.330 97.090 ;
        RECT 273.960 97.420 274.475 97.830 ;
        RECT 274.710 97.420 274.880 98.180 ;
        RECT 275.050 97.840 277.080 98.010 ;
        RECT 273.960 96.610 274.300 97.420 ;
        RECT 275.050 97.175 275.220 97.840 ;
        RECT 275.615 97.500 276.740 97.670 ;
        RECT 274.470 96.985 275.220 97.175 ;
        RECT 275.390 97.160 276.400 97.330 ;
        RECT 273.960 96.440 275.190 96.610 ;
        RECT 260.620 95.630 265.965 96.175 ;
        RECT 266.140 95.630 271.485 96.175 ;
        RECT 271.660 95.630 273.330 96.400 ;
        RECT 274.235 95.835 274.480 96.440 ;
        RECT 274.700 95.630 275.210 96.165 ;
        RECT 275.390 95.800 275.580 97.160 ;
        RECT 275.750 96.820 276.025 96.960 ;
        RECT 275.750 96.650 276.030 96.820 ;
        RECT 275.750 95.800 276.025 96.650 ;
        RECT 276.230 96.360 276.400 97.160 ;
        RECT 276.570 96.370 276.740 97.500 ;
        RECT 276.910 96.870 277.080 97.840 ;
        RECT 277.250 97.040 277.420 98.180 ;
        RECT 277.590 97.040 277.925 98.010 ;
        RECT 276.910 96.540 277.105 96.870 ;
        RECT 277.330 96.540 277.585 96.870 ;
        RECT 277.330 96.370 277.500 96.540 ;
        RECT 277.755 96.370 277.925 97.040 ;
        RECT 278.100 97.015 278.390 98.180 ;
        RECT 279.025 97.510 279.280 98.010 ;
        RECT 279.450 97.680 279.780 98.180 ;
        RECT 279.025 97.340 279.775 97.510 ;
        RECT 279.025 96.520 279.375 97.170 ;
        RECT 276.570 96.200 277.500 96.370 ;
        RECT 276.570 96.165 276.745 96.200 ;
        RECT 276.215 95.800 276.745 96.165 ;
        RECT 277.170 95.630 277.500 96.030 ;
        RECT 277.670 95.800 277.925 96.370 ;
        RECT 278.100 95.630 278.390 96.355 ;
        RECT 279.545 96.350 279.775 97.340 ;
        RECT 279.025 96.180 279.775 96.350 ;
        RECT 279.025 95.890 279.280 96.180 ;
        RECT 279.450 95.630 279.780 96.010 ;
        RECT 279.950 95.890 280.120 98.010 ;
        RECT 280.290 97.210 280.615 97.995 ;
        RECT 280.785 97.720 281.035 98.180 ;
        RECT 281.205 97.680 281.455 98.010 ;
        RECT 281.670 97.680 282.350 98.010 ;
        RECT 281.205 97.550 281.375 97.680 ;
        RECT 280.980 97.380 281.375 97.550 ;
        RECT 280.350 96.160 280.810 97.210 ;
        RECT 280.980 96.020 281.150 97.380 ;
        RECT 281.545 97.120 282.010 97.510 ;
        RECT 281.320 96.310 281.670 96.930 ;
        RECT 281.840 96.530 282.010 97.120 ;
        RECT 282.180 96.900 282.350 97.680 ;
        RECT 282.520 97.580 282.690 97.920 ;
        RECT 282.925 97.750 283.255 98.180 ;
        RECT 283.425 97.580 283.595 97.920 ;
        RECT 283.890 97.720 284.260 98.180 ;
        RECT 282.520 97.410 283.595 97.580 ;
        RECT 284.430 97.550 284.600 98.010 ;
        RECT 284.835 97.670 285.705 98.010 ;
        RECT 285.875 97.720 286.125 98.180 ;
        RECT 284.040 97.380 284.600 97.550 ;
        RECT 284.040 97.240 284.210 97.380 ;
        RECT 282.710 97.070 284.210 97.240 ;
        RECT 284.905 97.210 285.365 97.500 ;
        RECT 282.180 96.730 283.870 96.900 ;
        RECT 281.840 96.310 282.195 96.530 ;
        RECT 282.365 96.020 282.535 96.730 ;
        RECT 282.740 96.310 283.530 96.560 ;
        RECT 283.700 96.550 283.870 96.730 ;
        RECT 284.040 96.380 284.210 97.070 ;
        RECT 280.480 95.630 280.810 95.990 ;
        RECT 280.980 95.850 281.475 96.020 ;
        RECT 281.680 95.850 282.535 96.020 ;
        RECT 283.410 95.630 283.740 96.090 ;
        RECT 283.950 95.990 284.210 96.380 ;
        RECT 284.400 97.200 285.365 97.210 ;
        RECT 285.535 97.290 285.705 97.670 ;
        RECT 286.295 97.630 286.465 97.920 ;
        RECT 286.645 97.800 286.975 98.180 ;
        RECT 286.295 97.460 287.095 97.630 ;
        RECT 284.400 97.040 285.075 97.200 ;
        RECT 285.535 97.120 286.755 97.290 ;
        RECT 284.400 96.250 284.610 97.040 ;
        RECT 285.535 97.030 285.705 97.120 ;
        RECT 284.780 96.250 285.130 96.870 ;
        RECT 285.300 96.860 285.705 97.030 ;
        RECT 285.300 96.080 285.470 96.860 ;
        RECT 285.640 96.410 285.860 96.690 ;
        RECT 286.040 96.580 286.580 96.950 ;
        RECT 286.925 96.870 287.095 97.460 ;
        RECT 287.315 97.040 287.620 98.180 ;
        RECT 287.790 96.990 288.045 97.870 ;
        RECT 288.310 97.250 288.480 98.010 ;
        RECT 288.695 97.420 289.025 98.180 ;
        RECT 288.310 97.080 289.025 97.250 ;
        RECT 289.195 97.105 289.450 98.010 ;
        RECT 286.925 96.840 287.665 96.870 ;
        RECT 285.640 96.240 286.170 96.410 ;
        RECT 283.950 95.820 284.300 95.990 ;
        RECT 284.520 95.800 285.470 96.080 ;
        RECT 285.640 95.630 285.830 96.070 ;
        RECT 286.000 96.010 286.170 96.240 ;
        RECT 286.340 96.180 286.580 96.580 ;
        RECT 286.750 96.540 287.665 96.840 ;
        RECT 286.750 96.365 287.075 96.540 ;
        RECT 286.750 96.010 287.070 96.365 ;
        RECT 287.835 96.340 288.045 96.990 ;
        RECT 288.220 96.530 288.575 96.900 ;
        RECT 288.855 96.870 289.025 97.080 ;
        RECT 288.855 96.540 289.110 96.870 ;
        RECT 288.855 96.350 289.025 96.540 ;
        RECT 289.280 96.375 289.450 97.105 ;
        RECT 289.625 97.030 289.885 98.180 ;
        RECT 290.065 97.040 290.400 98.010 ;
        RECT 290.570 97.040 290.740 98.180 ;
        RECT 290.910 97.840 292.940 98.010 ;
        RECT 286.000 95.840 287.070 96.010 ;
        RECT 287.315 95.630 287.620 96.090 ;
        RECT 287.790 95.810 288.045 96.340 ;
        RECT 288.310 96.180 289.025 96.350 ;
        RECT 288.310 95.800 288.480 96.180 ;
        RECT 288.695 95.630 289.025 96.010 ;
        RECT 289.195 95.800 289.450 96.375 ;
        RECT 289.625 95.630 289.885 96.470 ;
        RECT 290.065 96.370 290.235 97.040 ;
        RECT 290.910 96.870 291.080 97.840 ;
        RECT 290.405 96.540 290.660 96.870 ;
        RECT 290.885 96.540 291.080 96.870 ;
        RECT 291.250 97.500 292.375 97.670 ;
        RECT 290.490 96.370 290.660 96.540 ;
        RECT 291.250 96.370 291.420 97.500 ;
        RECT 290.065 95.800 290.320 96.370 ;
        RECT 290.490 96.200 291.420 96.370 ;
        RECT 291.590 97.160 292.600 97.330 ;
        RECT 291.590 96.360 291.760 97.160 ;
        RECT 291.245 96.165 291.420 96.200 ;
        RECT 290.490 95.630 290.820 96.030 ;
        RECT 291.245 95.800 291.775 96.165 ;
        RECT 291.965 96.140 292.240 96.960 ;
        RECT 291.960 95.970 292.240 96.140 ;
        RECT 291.965 95.800 292.240 95.970 ;
        RECT 292.410 95.800 292.600 97.160 ;
        RECT 292.770 97.175 292.940 97.840 ;
        RECT 293.110 97.420 293.280 98.180 ;
        RECT 293.515 97.420 294.030 97.830 ;
        RECT 292.770 96.985 293.520 97.175 ;
        RECT 293.690 96.610 294.030 97.420 ;
        RECT 294.665 97.510 294.920 98.010 ;
        RECT 295.090 97.680 295.420 98.180 ;
        RECT 294.665 97.340 295.415 97.510 ;
        RECT 292.800 96.440 294.030 96.610 ;
        RECT 294.665 96.520 295.015 97.170 ;
        RECT 292.780 95.630 293.290 96.165 ;
        RECT 293.510 95.835 293.755 96.440 ;
        RECT 295.185 96.350 295.415 97.340 ;
        RECT 294.665 96.180 295.415 96.350 ;
        RECT 294.665 95.890 294.920 96.180 ;
        RECT 295.090 95.630 295.420 96.010 ;
        RECT 295.590 95.890 295.760 98.010 ;
        RECT 295.930 97.210 296.255 97.995 ;
        RECT 296.425 97.720 296.675 98.180 ;
        RECT 296.845 97.680 297.095 98.010 ;
        RECT 297.310 97.680 297.990 98.010 ;
        RECT 296.845 97.550 297.015 97.680 ;
        RECT 296.620 97.380 297.015 97.550 ;
        RECT 295.990 96.160 296.450 97.210 ;
        RECT 296.620 96.020 296.790 97.380 ;
        RECT 297.185 97.120 297.650 97.510 ;
        RECT 296.960 96.310 297.310 96.930 ;
        RECT 297.480 96.530 297.650 97.120 ;
        RECT 297.820 96.900 297.990 97.680 ;
        RECT 298.160 97.580 298.330 97.920 ;
        RECT 298.565 97.750 298.895 98.180 ;
        RECT 299.065 97.580 299.235 97.920 ;
        RECT 299.530 97.720 299.900 98.180 ;
        RECT 298.160 97.410 299.235 97.580 ;
        RECT 300.070 97.550 300.240 98.010 ;
        RECT 300.475 97.670 301.345 98.010 ;
        RECT 301.515 97.720 301.765 98.180 ;
        RECT 299.680 97.380 300.240 97.550 ;
        RECT 299.680 97.240 299.850 97.380 ;
        RECT 298.350 97.070 299.850 97.240 ;
        RECT 300.545 97.210 301.005 97.500 ;
        RECT 297.820 96.730 299.510 96.900 ;
        RECT 297.480 96.310 297.835 96.530 ;
        RECT 298.005 96.020 298.175 96.730 ;
        RECT 298.380 96.310 299.170 96.560 ;
        RECT 299.340 96.550 299.510 96.730 ;
        RECT 299.680 96.380 299.850 97.070 ;
        RECT 296.120 95.630 296.450 95.990 ;
        RECT 296.620 95.850 297.115 96.020 ;
        RECT 297.320 95.850 298.175 96.020 ;
        RECT 299.050 95.630 299.380 96.090 ;
        RECT 299.590 95.990 299.850 96.380 ;
        RECT 300.040 97.200 301.005 97.210 ;
        RECT 301.175 97.290 301.345 97.670 ;
        RECT 301.935 97.630 302.105 97.920 ;
        RECT 302.285 97.800 302.615 98.180 ;
        RECT 301.935 97.460 302.735 97.630 ;
        RECT 300.040 97.040 300.715 97.200 ;
        RECT 301.175 97.120 302.395 97.290 ;
        RECT 300.040 96.250 300.250 97.040 ;
        RECT 301.175 97.030 301.345 97.120 ;
        RECT 300.420 96.250 300.770 96.870 ;
        RECT 300.940 96.860 301.345 97.030 ;
        RECT 300.940 96.080 301.110 96.860 ;
        RECT 301.280 96.410 301.500 96.690 ;
        RECT 301.680 96.580 302.220 96.950 ;
        RECT 302.565 96.870 302.735 97.460 ;
        RECT 302.955 97.040 303.260 98.180 ;
        RECT 303.430 96.990 303.685 97.870 ;
        RECT 303.860 97.015 304.150 98.180 ;
        RECT 304.325 97.040 304.660 98.010 ;
        RECT 304.830 97.040 305.000 98.180 ;
        RECT 305.170 97.840 307.200 98.010 ;
        RECT 302.565 96.840 303.305 96.870 ;
        RECT 301.280 96.240 301.810 96.410 ;
        RECT 299.590 95.820 299.940 95.990 ;
        RECT 300.160 95.800 301.110 96.080 ;
        RECT 301.280 95.630 301.470 96.070 ;
        RECT 301.640 96.010 301.810 96.240 ;
        RECT 301.980 96.180 302.220 96.580 ;
        RECT 302.390 96.540 303.305 96.840 ;
        RECT 302.390 96.365 302.715 96.540 ;
        RECT 302.390 96.010 302.710 96.365 ;
        RECT 303.475 96.340 303.685 96.990 ;
        RECT 304.325 96.370 304.495 97.040 ;
        RECT 305.170 96.870 305.340 97.840 ;
        RECT 304.665 96.540 304.920 96.870 ;
        RECT 305.145 96.540 305.340 96.870 ;
        RECT 305.510 97.500 306.635 97.670 ;
        RECT 304.750 96.370 304.920 96.540 ;
        RECT 305.510 96.370 305.680 97.500 ;
        RECT 301.640 95.840 302.710 96.010 ;
        RECT 302.955 95.630 303.260 96.090 ;
        RECT 303.430 95.810 303.685 96.340 ;
        RECT 303.860 95.630 304.150 96.355 ;
        RECT 304.325 95.800 304.580 96.370 ;
        RECT 304.750 96.200 305.680 96.370 ;
        RECT 305.850 97.160 306.860 97.330 ;
        RECT 305.850 96.360 306.020 97.160 ;
        RECT 306.225 96.820 306.500 96.960 ;
        RECT 306.220 96.650 306.500 96.820 ;
        RECT 305.505 96.165 305.680 96.200 ;
        RECT 304.750 95.630 305.080 96.030 ;
        RECT 305.505 95.800 306.035 96.165 ;
        RECT 306.225 95.800 306.500 96.650 ;
        RECT 306.670 95.800 306.860 97.160 ;
        RECT 307.030 97.175 307.200 97.840 ;
        RECT 307.370 97.420 307.540 98.180 ;
        RECT 307.775 97.420 308.290 97.830 ;
        RECT 307.030 96.985 307.780 97.175 ;
        RECT 307.950 96.610 308.290 97.420 ;
        RECT 308.460 97.090 309.670 98.180 ;
        RECT 307.060 96.440 308.290 96.610 ;
        RECT 307.040 95.630 307.550 96.165 ;
        RECT 307.770 95.835 308.015 96.440 ;
        RECT 308.460 96.380 308.980 96.920 ;
        RECT 309.150 96.550 309.670 97.090 ;
        RECT 309.840 97.090 311.050 98.180 ;
        RECT 309.840 96.550 310.360 97.090 ;
        RECT 310.530 96.380 311.050 96.920 ;
        RECT 308.460 95.630 309.670 96.380 ;
        RECT 309.840 95.630 311.050 96.380 ;
        RECT 162.095 95.460 311.135 95.630 ;
        RECT 162.180 94.710 163.390 95.460 ;
        RECT 162.180 94.170 162.700 94.710 ;
        RECT 163.565 94.620 163.825 95.460 ;
        RECT 164.000 94.715 164.255 95.290 ;
        RECT 164.425 95.080 164.755 95.460 ;
        RECT 164.970 94.910 165.140 95.290 ;
        RECT 164.425 94.740 165.140 94.910 ;
        RECT 162.870 94.000 163.390 94.540 ;
        RECT 162.180 92.910 163.390 94.000 ;
        RECT 163.565 92.910 163.825 94.060 ;
        RECT 164.000 93.985 164.170 94.715 ;
        RECT 164.425 94.550 164.595 94.740 ;
        RECT 165.400 94.690 168.910 95.460 ;
        RECT 169.085 94.910 169.340 95.200 ;
        RECT 169.510 95.080 169.840 95.460 ;
        RECT 169.085 94.740 169.835 94.910 ;
        RECT 164.340 94.220 164.595 94.550 ;
        RECT 164.425 94.010 164.595 94.220 ;
        RECT 164.875 94.190 165.230 94.560 ;
        RECT 165.400 94.170 167.050 94.690 ;
        RECT 164.000 93.080 164.255 93.985 ;
        RECT 164.425 93.840 165.140 94.010 ;
        RECT 167.220 94.000 168.910 94.520 ;
        RECT 164.425 92.910 164.755 93.670 ;
        RECT 164.970 93.080 165.140 93.840 ;
        RECT 165.400 92.910 168.910 94.000 ;
        RECT 169.085 93.920 169.435 94.570 ;
        RECT 169.605 93.750 169.835 94.740 ;
        RECT 169.085 93.580 169.835 93.750 ;
        RECT 169.085 93.080 169.340 93.580 ;
        RECT 169.510 92.910 169.840 93.410 ;
        RECT 170.010 93.080 170.180 95.200 ;
        RECT 170.540 95.100 170.870 95.460 ;
        RECT 171.040 95.070 171.535 95.240 ;
        RECT 171.740 95.070 172.595 95.240 ;
        RECT 170.410 93.880 170.870 94.930 ;
        RECT 170.350 93.095 170.675 93.880 ;
        RECT 171.040 93.710 171.210 95.070 ;
        RECT 171.380 94.160 171.730 94.780 ;
        RECT 171.900 94.560 172.255 94.780 ;
        RECT 171.900 93.970 172.070 94.560 ;
        RECT 172.425 94.360 172.595 95.070 ;
        RECT 173.470 95.000 173.800 95.460 ;
        RECT 174.010 95.100 174.360 95.270 ;
        RECT 172.800 94.530 173.590 94.780 ;
        RECT 174.010 94.710 174.270 95.100 ;
        RECT 174.580 95.010 175.530 95.290 ;
        RECT 175.700 95.020 175.890 95.460 ;
        RECT 176.060 95.080 177.130 95.250 ;
        RECT 173.760 94.360 173.930 94.540 ;
        RECT 171.040 93.540 171.435 93.710 ;
        RECT 171.605 93.580 172.070 93.970 ;
        RECT 172.240 94.190 173.930 94.360 ;
        RECT 171.265 93.410 171.435 93.540 ;
        RECT 172.240 93.410 172.410 94.190 ;
        RECT 174.100 94.020 174.270 94.710 ;
        RECT 172.770 93.850 174.270 94.020 ;
        RECT 174.460 94.050 174.670 94.840 ;
        RECT 174.840 94.220 175.190 94.840 ;
        RECT 175.360 94.230 175.530 95.010 ;
        RECT 176.060 94.850 176.230 95.080 ;
        RECT 175.700 94.680 176.230 94.850 ;
        RECT 175.700 94.400 175.920 94.680 ;
        RECT 176.400 94.510 176.640 94.910 ;
        RECT 175.360 94.060 175.765 94.230 ;
        RECT 176.100 94.140 176.640 94.510 ;
        RECT 176.810 94.725 177.130 95.080 ;
        RECT 177.375 95.000 177.680 95.460 ;
        RECT 177.850 94.750 178.100 95.280 ;
        RECT 176.810 94.550 177.135 94.725 ;
        RECT 176.810 94.250 177.725 94.550 ;
        RECT 176.985 94.220 177.725 94.250 ;
        RECT 174.460 93.890 175.135 94.050 ;
        RECT 175.595 93.970 175.765 94.060 ;
        RECT 174.460 93.880 175.425 93.890 ;
        RECT 174.100 93.710 174.270 93.850 ;
        RECT 170.845 92.910 171.095 93.370 ;
        RECT 171.265 93.080 171.515 93.410 ;
        RECT 171.730 93.080 172.410 93.410 ;
        RECT 172.580 93.510 173.655 93.680 ;
        RECT 174.100 93.540 174.660 93.710 ;
        RECT 174.965 93.590 175.425 93.880 ;
        RECT 175.595 93.800 176.815 93.970 ;
        RECT 172.580 93.170 172.750 93.510 ;
        RECT 172.985 92.910 173.315 93.340 ;
        RECT 173.485 93.170 173.655 93.510 ;
        RECT 173.950 92.910 174.320 93.370 ;
        RECT 174.490 93.080 174.660 93.540 ;
        RECT 175.595 93.420 175.765 93.800 ;
        RECT 176.985 93.630 177.155 94.220 ;
        RECT 177.895 94.100 178.100 94.750 ;
        RECT 178.270 94.705 178.520 95.460 ;
        RECT 178.740 94.915 184.085 95.460 ;
        RECT 174.895 93.080 175.765 93.420 ;
        RECT 176.355 93.460 177.155 93.630 ;
        RECT 175.935 92.910 176.185 93.370 ;
        RECT 176.355 93.170 176.525 93.460 ;
        RECT 176.705 92.910 177.035 93.290 ;
        RECT 177.375 92.910 177.680 94.050 ;
        RECT 177.850 93.220 178.100 94.100 ;
        RECT 180.325 94.085 180.665 94.915 ;
        RECT 184.260 94.690 187.770 95.460 ;
        RECT 187.940 94.735 188.230 95.460 ;
        RECT 188.405 94.720 188.660 95.290 ;
        RECT 188.830 95.060 189.160 95.460 ;
        RECT 189.585 94.925 190.115 95.290 ;
        RECT 190.305 95.120 190.580 95.290 ;
        RECT 190.300 94.950 190.580 95.120 ;
        RECT 189.585 94.890 189.760 94.925 ;
        RECT 188.830 94.720 189.760 94.890 ;
        RECT 178.270 92.910 178.520 94.050 ;
        RECT 182.145 93.345 182.495 94.595 ;
        RECT 184.260 94.170 185.910 94.690 ;
        RECT 186.080 94.000 187.770 94.520 ;
        RECT 178.740 92.910 184.085 93.345 ;
        RECT 184.260 92.910 187.770 94.000 ;
        RECT 187.940 92.910 188.230 94.075 ;
        RECT 188.405 94.050 188.575 94.720 ;
        RECT 188.830 94.550 189.000 94.720 ;
        RECT 188.745 94.220 189.000 94.550 ;
        RECT 189.225 94.220 189.420 94.550 ;
        RECT 188.405 93.080 188.740 94.050 ;
        RECT 188.910 92.910 189.080 94.050 ;
        RECT 189.250 93.250 189.420 94.220 ;
        RECT 189.590 93.590 189.760 94.720 ;
        RECT 189.930 93.930 190.100 94.730 ;
        RECT 190.305 94.130 190.580 94.950 ;
        RECT 190.750 93.930 190.940 95.290 ;
        RECT 191.120 94.925 191.630 95.460 ;
        RECT 191.850 94.650 192.095 95.255 ;
        RECT 191.140 94.480 192.370 94.650 ;
        RECT 189.930 93.760 190.940 93.930 ;
        RECT 191.110 93.915 191.860 94.105 ;
        RECT 189.590 93.420 190.715 93.590 ;
        RECT 191.110 93.250 191.280 93.915 ;
        RECT 192.030 93.670 192.370 94.480 ;
        RECT 189.250 93.080 191.280 93.250 ;
        RECT 191.450 92.910 191.620 93.670 ;
        RECT 191.855 93.260 192.370 93.670 ;
        RECT 192.540 94.515 192.880 95.290 ;
        RECT 193.050 95.000 193.220 95.460 ;
        RECT 193.460 95.025 193.820 95.290 ;
        RECT 193.460 95.020 193.815 95.025 ;
        RECT 193.460 95.010 193.810 95.020 ;
        RECT 193.460 95.005 193.805 95.010 ;
        RECT 193.460 94.995 193.800 95.005 ;
        RECT 194.450 95.000 194.620 95.460 ;
        RECT 193.460 94.990 193.795 94.995 ;
        RECT 193.460 94.980 193.785 94.990 ;
        RECT 193.460 94.970 193.775 94.980 ;
        RECT 193.460 94.830 193.760 94.970 ;
        RECT 193.050 94.640 193.760 94.830 ;
        RECT 193.950 94.830 194.280 94.910 ;
        RECT 194.790 94.830 195.130 95.290 ;
        RECT 195.300 94.915 200.645 95.460 ;
        RECT 200.820 94.915 206.165 95.460 ;
        RECT 193.950 94.640 195.130 94.830 ;
        RECT 192.540 93.080 192.820 94.515 ;
        RECT 193.050 94.070 193.335 94.640 ;
        RECT 193.520 94.240 193.990 94.470 ;
        RECT 194.160 94.450 194.490 94.470 ;
        RECT 194.160 94.270 194.610 94.450 ;
        RECT 194.800 94.270 195.130 94.470 ;
        RECT 193.050 93.855 194.200 94.070 ;
        RECT 192.990 92.910 193.700 93.685 ;
        RECT 193.870 93.080 194.200 93.855 ;
        RECT 194.395 93.155 194.610 94.270 ;
        RECT 194.900 93.930 195.130 94.270 ;
        RECT 196.885 94.085 197.225 94.915 ;
        RECT 194.790 92.910 195.120 93.630 ;
        RECT 198.705 93.345 199.055 94.595 ;
        RECT 202.405 94.085 202.745 94.915 ;
        RECT 204.225 93.345 204.575 94.595 ;
        RECT 195.300 92.910 200.645 93.345 ;
        RECT 200.820 92.910 206.165 93.345 ;
        RECT 206.350 93.090 206.610 95.280 ;
        RECT 206.870 95.090 207.540 95.460 ;
        RECT 207.720 94.910 208.030 95.280 ;
        RECT 206.800 94.710 208.030 94.910 ;
        RECT 206.800 94.040 207.090 94.710 ;
        RECT 208.210 94.530 208.440 95.170 ;
        RECT 208.620 94.730 208.910 95.460 ;
        RECT 209.105 94.695 209.560 95.460 ;
        RECT 209.835 95.080 211.135 95.290 ;
        RECT 211.390 95.100 211.720 95.460 ;
        RECT 210.965 94.930 211.135 95.080 ;
        RECT 211.890 94.960 212.150 95.290 ;
        RECT 207.270 94.220 207.735 94.530 ;
        RECT 207.915 94.220 208.440 94.530 ;
        RECT 208.620 94.220 208.920 94.550 ;
        RECT 210.035 94.470 210.255 94.870 ;
        RECT 209.100 94.270 209.590 94.470 ;
        RECT 209.780 94.260 210.255 94.470 ;
        RECT 210.500 94.470 210.710 94.870 ;
        RECT 210.965 94.805 211.720 94.930 ;
        RECT 210.965 94.760 211.810 94.805 ;
        RECT 211.540 94.640 211.810 94.760 ;
        RECT 210.500 94.260 210.830 94.470 ;
        RECT 211.000 94.200 211.410 94.505 ;
        RECT 206.800 93.820 207.570 94.040 ;
        RECT 206.780 92.910 207.120 93.640 ;
        RECT 207.300 93.090 207.570 93.820 ;
        RECT 207.750 93.800 208.910 94.040 ;
        RECT 207.750 93.090 207.980 93.800 ;
        RECT 208.150 92.910 208.480 93.620 ;
        RECT 208.650 93.090 208.910 93.800 ;
        RECT 209.105 94.030 210.280 94.090 ;
        RECT 211.640 94.065 211.810 94.640 ;
        RECT 211.610 94.030 211.810 94.065 ;
        RECT 209.105 93.920 211.810 94.030 ;
        RECT 209.105 93.300 209.360 93.920 ;
        RECT 209.950 93.860 211.750 93.920 ;
        RECT 209.950 93.830 210.280 93.860 ;
        RECT 211.980 93.760 212.150 94.960 ;
        RECT 212.320 94.710 213.530 95.460 ;
        RECT 213.700 94.735 213.990 95.460 ;
        RECT 214.160 94.915 219.505 95.460 ;
        RECT 212.320 94.170 212.840 94.710 ;
        RECT 213.010 94.000 213.530 94.540 ;
        RECT 215.745 94.085 216.085 94.915 ;
        RECT 219.680 94.690 223.190 95.460 ;
        RECT 224.280 94.960 224.540 95.290 ;
        RECT 224.710 95.100 225.040 95.460 ;
        RECT 225.295 95.080 226.595 95.290 ;
        RECT 209.610 93.660 209.795 93.750 ;
        RECT 210.385 93.660 211.220 93.670 ;
        RECT 209.610 93.460 211.220 93.660 ;
        RECT 209.610 93.420 209.840 93.460 ;
        RECT 209.105 93.080 209.440 93.300 ;
        RECT 210.445 92.910 210.800 93.290 ;
        RECT 210.970 93.080 211.220 93.460 ;
        RECT 211.470 92.910 211.720 93.690 ;
        RECT 211.890 93.080 212.150 93.760 ;
        RECT 212.320 92.910 213.530 94.000 ;
        RECT 213.700 92.910 213.990 94.075 ;
        RECT 217.565 93.345 217.915 94.595 ;
        RECT 219.680 94.170 221.330 94.690 ;
        RECT 221.500 94.000 223.190 94.520 ;
        RECT 214.160 92.910 219.505 93.345 ;
        RECT 219.680 92.910 223.190 94.000 ;
        RECT 224.280 93.760 224.450 94.960 ;
        RECT 225.295 94.930 225.465 95.080 ;
        RECT 224.710 94.805 225.465 94.930 ;
        RECT 224.620 94.760 225.465 94.805 ;
        RECT 224.620 94.640 224.890 94.760 ;
        RECT 224.620 94.065 224.790 94.640 ;
        RECT 225.020 94.200 225.430 94.505 ;
        RECT 225.720 94.470 225.930 94.870 ;
        RECT 225.600 94.260 225.930 94.470 ;
        RECT 226.175 94.470 226.395 94.870 ;
        RECT 226.870 94.695 227.325 95.460 ;
        RECT 227.505 94.695 227.960 95.460 ;
        RECT 228.235 95.080 229.535 95.290 ;
        RECT 229.790 95.100 230.120 95.460 ;
        RECT 229.365 94.930 229.535 95.080 ;
        RECT 230.290 94.960 230.550 95.290 ;
        RECT 228.435 94.470 228.655 94.870 ;
        RECT 226.175 94.260 226.650 94.470 ;
        RECT 226.840 94.270 227.330 94.470 ;
        RECT 227.500 94.270 227.990 94.470 ;
        RECT 228.180 94.260 228.655 94.470 ;
        RECT 228.900 94.470 229.110 94.870 ;
        RECT 229.365 94.805 230.120 94.930 ;
        RECT 229.365 94.760 230.210 94.805 ;
        RECT 229.940 94.640 230.210 94.760 ;
        RECT 228.900 94.260 229.230 94.470 ;
        RECT 229.400 94.200 229.810 94.505 ;
        RECT 224.620 94.030 224.820 94.065 ;
        RECT 226.150 94.030 227.325 94.090 ;
        RECT 224.620 93.920 227.325 94.030 ;
        RECT 224.680 93.860 226.480 93.920 ;
        RECT 226.150 93.830 226.480 93.860 ;
        RECT 224.280 93.080 224.540 93.760 ;
        RECT 224.710 92.910 224.960 93.690 ;
        RECT 225.210 93.660 226.045 93.670 ;
        RECT 226.635 93.660 226.820 93.750 ;
        RECT 225.210 93.460 226.820 93.660 ;
        RECT 225.210 93.080 225.460 93.460 ;
        RECT 226.590 93.420 226.820 93.460 ;
        RECT 227.070 93.300 227.325 93.920 ;
        RECT 225.630 92.910 225.985 93.290 ;
        RECT 226.990 93.080 227.325 93.300 ;
        RECT 227.505 94.030 228.680 94.090 ;
        RECT 230.040 94.065 230.210 94.640 ;
        RECT 230.010 94.030 230.210 94.065 ;
        RECT 227.505 93.920 230.210 94.030 ;
        RECT 227.505 93.300 227.760 93.920 ;
        RECT 228.350 93.860 230.150 93.920 ;
        RECT 228.350 93.830 228.680 93.860 ;
        RECT 230.380 93.760 230.550 94.960 ;
        RECT 230.720 94.915 236.065 95.460 ;
        RECT 232.305 94.085 232.645 94.915 ;
        RECT 236.240 94.690 238.830 95.460 ;
        RECT 239.460 94.735 239.750 95.460 ;
        RECT 239.920 94.710 241.130 95.460 ;
        RECT 241.320 94.960 241.575 95.290 ;
        RECT 241.790 94.980 242.120 95.460 ;
        RECT 242.290 95.040 243.825 95.290 ;
        RECT 241.320 94.950 241.530 94.960 ;
        RECT 241.320 94.880 241.505 94.950 ;
        RECT 228.010 93.660 228.195 93.750 ;
        RECT 228.785 93.660 229.620 93.670 ;
        RECT 228.010 93.460 229.620 93.660 ;
        RECT 228.010 93.420 228.240 93.460 ;
        RECT 227.505 93.080 227.840 93.300 ;
        RECT 228.845 92.910 229.200 93.290 ;
        RECT 229.370 93.080 229.620 93.460 ;
        RECT 229.870 92.910 230.120 93.690 ;
        RECT 230.290 93.080 230.550 93.760 ;
        RECT 234.125 93.345 234.475 94.595 ;
        RECT 236.240 94.170 237.450 94.690 ;
        RECT 237.620 94.000 238.830 94.520 ;
        RECT 239.920 94.170 240.440 94.710 ;
        RECT 230.720 92.910 236.065 93.345 ;
        RECT 236.240 92.910 238.830 94.000 ;
        RECT 239.460 92.910 239.750 94.075 ;
        RECT 240.610 94.000 241.130 94.540 ;
        RECT 239.920 92.910 241.130 94.000 ;
        RECT 241.320 93.750 241.490 94.880 ;
        RECT 242.290 94.810 242.460 95.040 ;
        RECT 241.660 94.640 242.460 94.810 ;
        RECT 241.660 94.090 241.830 94.640 ;
        RECT 242.640 94.470 242.925 94.870 ;
        RECT 242.060 94.440 242.425 94.470 ;
        RECT 242.050 94.270 242.425 94.440 ;
        RECT 242.595 94.270 242.925 94.470 ;
        RECT 243.195 94.470 243.475 94.870 ;
        RECT 243.655 94.810 243.825 95.040 ;
        RECT 244.050 94.980 244.380 95.460 ;
        RECT 244.550 94.810 244.720 95.290 ;
        RECT 243.655 94.640 244.720 94.810 ;
        RECT 244.985 94.695 245.440 95.460 ;
        RECT 245.715 95.080 247.015 95.290 ;
        RECT 247.270 95.100 247.600 95.460 ;
        RECT 246.845 94.930 247.015 95.080 ;
        RECT 247.770 94.960 248.030 95.290 ;
        RECT 245.915 94.470 246.135 94.870 ;
        RECT 243.195 94.270 243.670 94.470 ;
        RECT 243.840 94.270 244.285 94.470 ;
        RECT 244.455 94.260 244.805 94.470 ;
        RECT 244.980 94.270 245.470 94.470 ;
        RECT 245.660 94.260 246.135 94.470 ;
        RECT 246.380 94.470 246.590 94.870 ;
        RECT 246.845 94.805 247.600 94.930 ;
        RECT 246.845 94.760 247.690 94.805 ;
        RECT 247.420 94.640 247.690 94.760 ;
        RECT 246.380 94.260 246.710 94.470 ;
        RECT 246.880 94.200 247.290 94.505 ;
        RECT 241.660 93.920 244.720 94.090 ;
        RECT 241.320 93.080 241.575 93.750 ;
        RECT 241.745 92.910 242.075 93.670 ;
        RECT 242.245 93.510 243.880 93.750 ;
        RECT 242.245 93.080 242.495 93.510 ;
        RECT 243.650 93.420 243.880 93.510 ;
        RECT 242.665 92.910 243.020 93.330 ;
        RECT 243.210 93.250 243.540 93.290 ;
        RECT 244.050 93.250 244.380 93.750 ;
        RECT 243.210 93.080 244.380 93.250 ;
        RECT 244.550 93.080 244.720 93.920 ;
        RECT 244.985 94.030 246.160 94.090 ;
        RECT 247.520 94.065 247.690 94.640 ;
        RECT 247.490 94.030 247.690 94.065 ;
        RECT 244.985 93.920 247.690 94.030 ;
        RECT 244.985 93.300 245.240 93.920 ;
        RECT 245.830 93.860 247.630 93.920 ;
        RECT 245.830 93.830 246.160 93.860 ;
        RECT 247.860 93.760 248.030 94.960 ;
        RECT 245.490 93.660 245.675 93.750 ;
        RECT 246.265 93.660 247.100 93.670 ;
        RECT 245.490 93.460 247.100 93.660 ;
        RECT 245.490 93.420 245.720 93.460 ;
        RECT 244.985 93.080 245.320 93.300 ;
        RECT 246.325 92.910 246.680 93.290 ;
        RECT 246.850 93.080 247.100 93.460 ;
        RECT 247.350 92.910 247.600 93.690 ;
        RECT 247.770 93.080 248.030 93.760 ;
        RECT 248.220 94.960 248.475 95.290 ;
        RECT 248.690 94.980 249.020 95.460 ;
        RECT 249.190 95.040 250.725 95.290 ;
        RECT 248.220 94.950 248.430 94.960 ;
        RECT 248.220 94.880 248.405 94.950 ;
        RECT 248.220 93.750 248.390 94.880 ;
        RECT 249.190 94.810 249.360 95.040 ;
        RECT 248.560 94.640 249.360 94.810 ;
        RECT 248.560 94.090 248.730 94.640 ;
        RECT 249.540 94.470 249.825 94.870 ;
        RECT 248.960 94.270 249.325 94.470 ;
        RECT 249.495 94.270 249.825 94.470 ;
        RECT 250.095 94.470 250.375 94.870 ;
        RECT 250.555 94.810 250.725 95.040 ;
        RECT 250.950 94.980 251.280 95.460 ;
        RECT 251.450 94.810 251.620 95.290 ;
        RECT 251.880 94.915 257.225 95.460 ;
        RECT 250.555 94.640 251.620 94.810 ;
        RECT 250.095 94.270 250.570 94.470 ;
        RECT 250.740 94.270 251.185 94.470 ;
        RECT 251.355 94.260 251.705 94.470 ;
        RECT 248.560 93.920 251.620 94.090 ;
        RECT 253.465 94.085 253.805 94.915 ;
        RECT 258.410 94.810 258.580 95.290 ;
        RECT 258.750 94.980 259.080 95.460 ;
        RECT 259.305 95.040 260.840 95.290 ;
        RECT 259.305 94.810 259.475 95.040 ;
        RECT 258.410 94.640 259.475 94.810 ;
        RECT 248.220 93.080 248.475 93.750 ;
        RECT 248.645 92.910 248.975 93.670 ;
        RECT 249.145 93.510 250.780 93.750 ;
        RECT 249.145 93.080 249.395 93.510 ;
        RECT 250.550 93.420 250.780 93.510 ;
        RECT 249.565 92.910 249.920 93.330 ;
        RECT 250.110 93.250 250.440 93.290 ;
        RECT 250.950 93.250 251.280 93.750 ;
        RECT 250.110 93.080 251.280 93.250 ;
        RECT 251.450 93.080 251.620 93.920 ;
        RECT 255.285 93.345 255.635 94.595 ;
        RECT 259.655 94.470 259.935 94.870 ;
        RECT 258.325 94.260 258.675 94.470 ;
        RECT 258.845 94.270 259.290 94.470 ;
        RECT 259.460 94.270 259.935 94.470 ;
        RECT 260.205 94.470 260.490 94.870 ;
        RECT 260.670 94.810 260.840 95.040 ;
        RECT 261.010 94.980 261.340 95.460 ;
        RECT 261.555 94.960 261.810 95.290 ;
        RECT 261.625 94.880 261.810 94.960 ;
        RECT 260.670 94.640 261.470 94.810 ;
        RECT 260.205 94.270 260.535 94.470 ;
        RECT 260.705 94.270 261.070 94.470 ;
        RECT 261.300 94.090 261.470 94.640 ;
        RECT 258.410 93.920 261.470 94.090 ;
        RECT 251.880 92.910 257.225 93.345 ;
        RECT 258.410 93.080 258.580 93.920 ;
        RECT 261.640 93.750 261.810 94.880 ;
        RECT 262.005 94.695 262.460 95.460 ;
        RECT 262.735 95.080 264.035 95.290 ;
        RECT 264.290 95.100 264.620 95.460 ;
        RECT 263.865 94.930 264.035 95.080 ;
        RECT 264.790 94.960 265.050 95.290 ;
        RECT 262.935 94.470 263.155 94.870 ;
        RECT 262.000 94.270 262.490 94.470 ;
        RECT 262.680 94.260 263.155 94.470 ;
        RECT 263.400 94.470 263.610 94.870 ;
        RECT 263.865 94.805 264.620 94.930 ;
        RECT 263.865 94.760 264.710 94.805 ;
        RECT 264.440 94.640 264.710 94.760 ;
        RECT 263.400 94.260 263.730 94.470 ;
        RECT 263.900 94.200 264.310 94.505 ;
        RECT 258.750 93.250 259.080 93.750 ;
        RECT 259.250 93.510 260.885 93.750 ;
        RECT 259.250 93.420 259.480 93.510 ;
        RECT 259.590 93.250 259.920 93.290 ;
        RECT 258.750 93.080 259.920 93.250 ;
        RECT 260.110 92.910 260.465 93.330 ;
        RECT 260.635 93.080 260.885 93.510 ;
        RECT 261.055 92.910 261.385 93.670 ;
        RECT 261.555 93.080 261.810 93.750 ;
        RECT 262.005 94.030 263.180 94.090 ;
        RECT 264.540 94.065 264.710 94.640 ;
        RECT 264.510 94.030 264.710 94.065 ;
        RECT 262.005 93.920 264.710 94.030 ;
        RECT 262.005 93.300 262.260 93.920 ;
        RECT 262.850 93.860 264.650 93.920 ;
        RECT 262.850 93.830 263.180 93.860 ;
        RECT 264.880 93.760 265.050 94.960 ;
        RECT 265.220 94.735 265.510 95.460 ;
        RECT 265.680 94.915 271.025 95.460 ;
        RECT 271.200 94.915 276.545 95.460 ;
        RECT 267.265 94.085 267.605 94.915 ;
        RECT 262.510 93.660 262.695 93.750 ;
        RECT 263.285 93.660 264.120 93.670 ;
        RECT 262.510 93.460 264.120 93.660 ;
        RECT 262.510 93.420 262.740 93.460 ;
        RECT 262.005 93.080 262.340 93.300 ;
        RECT 263.345 92.910 263.700 93.290 ;
        RECT 263.870 93.080 264.120 93.460 ;
        RECT 264.370 92.910 264.620 93.690 ;
        RECT 264.790 93.080 265.050 93.760 ;
        RECT 265.220 92.910 265.510 94.075 ;
        RECT 269.085 93.345 269.435 94.595 ;
        RECT 272.785 94.085 273.125 94.915 ;
        RECT 274.605 93.345 274.955 94.595 ;
        RECT 277.180 94.515 277.520 95.290 ;
        RECT 277.690 95.000 277.860 95.460 ;
        RECT 278.100 95.025 278.460 95.290 ;
        RECT 278.100 95.020 278.455 95.025 ;
        RECT 278.100 95.010 278.450 95.020 ;
        RECT 278.100 95.005 278.445 95.010 ;
        RECT 278.100 94.995 278.440 95.005 ;
        RECT 279.090 95.000 279.260 95.460 ;
        RECT 278.100 94.990 278.435 94.995 ;
        RECT 278.100 94.980 278.425 94.990 ;
        RECT 278.100 94.970 278.415 94.980 ;
        RECT 278.100 94.830 278.400 94.970 ;
        RECT 277.690 94.640 278.400 94.830 ;
        RECT 278.590 94.830 278.920 94.910 ;
        RECT 279.430 94.830 279.770 95.290 ;
        RECT 278.590 94.640 279.770 94.830 ;
        RECT 279.945 94.720 280.200 95.290 ;
        RECT 280.370 95.060 280.700 95.460 ;
        RECT 281.125 94.925 281.655 95.290 ;
        RECT 281.125 94.890 281.300 94.925 ;
        RECT 280.370 94.720 281.300 94.890 ;
        RECT 281.845 94.780 282.120 95.290 ;
        RECT 265.680 92.910 271.025 93.345 ;
        RECT 271.200 92.910 276.545 93.345 ;
        RECT 277.180 93.080 277.460 94.515 ;
        RECT 277.690 94.070 277.975 94.640 ;
        RECT 278.160 94.240 278.630 94.470 ;
        RECT 278.800 94.450 279.130 94.470 ;
        RECT 278.800 94.270 279.250 94.450 ;
        RECT 279.440 94.270 279.770 94.470 ;
        RECT 277.690 93.855 278.840 94.070 ;
        RECT 277.630 92.910 278.340 93.685 ;
        RECT 278.510 93.080 278.840 93.855 ;
        RECT 279.035 93.155 279.250 94.270 ;
        RECT 279.540 93.930 279.770 94.270 ;
        RECT 279.945 94.050 280.115 94.720 ;
        RECT 280.370 94.550 280.540 94.720 ;
        RECT 280.285 94.220 280.540 94.550 ;
        RECT 280.765 94.220 280.960 94.550 ;
        RECT 279.430 92.910 279.760 93.630 ;
        RECT 279.945 93.080 280.280 94.050 ;
        RECT 280.450 92.910 280.620 94.050 ;
        RECT 280.790 93.250 280.960 94.220 ;
        RECT 281.130 93.590 281.300 94.720 ;
        RECT 281.470 93.930 281.640 94.730 ;
        RECT 281.840 94.610 282.120 94.780 ;
        RECT 281.845 94.130 282.120 94.610 ;
        RECT 282.290 93.930 282.480 95.290 ;
        RECT 282.660 94.925 283.170 95.460 ;
        RECT 283.390 94.650 283.635 95.255 ;
        RECT 284.080 94.830 284.420 95.290 ;
        RECT 284.590 95.000 284.760 95.460 ;
        RECT 285.390 95.025 285.750 95.290 ;
        RECT 285.395 95.020 285.750 95.025 ;
        RECT 285.400 95.010 285.750 95.020 ;
        RECT 285.405 95.005 285.750 95.010 ;
        RECT 285.410 94.995 285.750 95.005 ;
        RECT 285.990 95.000 286.160 95.460 ;
        RECT 285.415 94.990 285.750 94.995 ;
        RECT 285.425 94.980 285.750 94.990 ;
        RECT 285.435 94.970 285.750 94.980 ;
        RECT 284.930 94.830 285.260 94.910 ;
        RECT 282.680 94.480 283.910 94.650 ;
        RECT 284.080 94.640 285.260 94.830 ;
        RECT 285.450 94.830 285.750 94.970 ;
        RECT 285.450 94.640 286.160 94.830 ;
        RECT 281.470 93.760 282.480 93.930 ;
        RECT 282.650 93.915 283.400 94.105 ;
        RECT 281.130 93.420 282.255 93.590 ;
        RECT 282.650 93.250 282.820 93.915 ;
        RECT 283.570 93.670 283.910 94.480 ;
        RECT 284.080 94.270 284.410 94.470 ;
        RECT 284.720 94.450 285.050 94.470 ;
        RECT 284.600 94.270 285.050 94.450 ;
        RECT 284.080 93.930 284.310 94.270 ;
        RECT 280.790 93.080 282.820 93.250 ;
        RECT 282.990 92.910 283.160 93.670 ;
        RECT 283.395 93.260 283.910 93.670 ;
        RECT 284.090 92.910 284.420 93.630 ;
        RECT 284.600 93.155 284.815 94.270 ;
        RECT 285.220 94.240 285.690 94.470 ;
        RECT 285.875 94.070 286.160 94.640 ;
        RECT 286.330 94.515 286.670 95.290 ;
        RECT 285.010 93.855 286.160 94.070 ;
        RECT 285.010 93.080 285.340 93.855 ;
        RECT 285.510 92.910 286.220 93.685 ;
        RECT 286.390 93.080 286.670 94.515 ;
        RECT 286.840 94.690 290.350 95.460 ;
        RECT 290.980 94.735 291.270 95.460 ;
        RECT 286.840 94.170 288.490 94.690 ;
        RECT 292.635 94.650 292.880 95.255 ;
        RECT 293.100 94.925 293.610 95.460 ;
        RECT 288.660 94.000 290.350 94.520 ;
        RECT 292.360 94.480 293.590 94.650 ;
        RECT 286.840 92.910 290.350 94.000 ;
        RECT 290.980 92.910 291.270 94.075 ;
        RECT 292.360 93.670 292.700 94.480 ;
        RECT 292.870 93.915 293.620 94.105 ;
        RECT 292.360 93.260 292.875 93.670 ;
        RECT 293.110 92.910 293.280 93.670 ;
        RECT 293.450 93.250 293.620 93.915 ;
        RECT 293.790 93.930 293.980 95.290 ;
        RECT 294.150 94.780 294.425 95.290 ;
        RECT 294.615 94.925 295.145 95.290 ;
        RECT 295.570 95.060 295.900 95.460 ;
        RECT 294.970 94.890 295.145 94.925 ;
        RECT 294.150 94.610 294.430 94.780 ;
        RECT 294.150 94.130 294.425 94.610 ;
        RECT 294.630 93.930 294.800 94.730 ;
        RECT 293.790 93.760 294.800 93.930 ;
        RECT 294.970 94.720 295.900 94.890 ;
        RECT 296.070 94.720 296.325 95.290 ;
        RECT 296.505 94.910 296.760 95.200 ;
        RECT 296.930 95.080 297.260 95.460 ;
        RECT 296.505 94.740 297.255 94.910 ;
        RECT 294.970 93.590 295.140 94.720 ;
        RECT 295.730 94.550 295.900 94.720 ;
        RECT 294.015 93.420 295.140 93.590 ;
        RECT 295.310 94.220 295.505 94.550 ;
        RECT 295.730 94.220 295.985 94.550 ;
        RECT 295.310 93.250 295.480 94.220 ;
        RECT 296.155 94.050 296.325 94.720 ;
        RECT 293.450 93.080 295.480 93.250 ;
        RECT 295.650 92.910 295.820 94.050 ;
        RECT 295.990 93.080 296.325 94.050 ;
        RECT 296.505 93.920 296.855 94.570 ;
        RECT 297.025 93.750 297.255 94.740 ;
        RECT 296.505 93.580 297.255 93.750 ;
        RECT 296.505 93.080 296.760 93.580 ;
        RECT 296.930 92.910 297.260 93.410 ;
        RECT 297.430 93.080 297.600 95.200 ;
        RECT 297.960 95.100 298.290 95.460 ;
        RECT 298.460 95.070 298.955 95.240 ;
        RECT 299.160 95.070 300.015 95.240 ;
        RECT 297.830 93.880 298.290 94.930 ;
        RECT 297.770 93.095 298.095 93.880 ;
        RECT 298.460 93.710 298.630 95.070 ;
        RECT 298.800 94.160 299.150 94.780 ;
        RECT 299.320 94.560 299.675 94.780 ;
        RECT 299.320 93.970 299.490 94.560 ;
        RECT 299.845 94.360 300.015 95.070 ;
        RECT 300.890 95.000 301.220 95.460 ;
        RECT 301.430 95.100 301.780 95.270 ;
        RECT 300.220 94.530 301.010 94.780 ;
        RECT 301.430 94.710 301.690 95.100 ;
        RECT 302.000 95.010 302.950 95.290 ;
        RECT 303.120 95.020 303.310 95.460 ;
        RECT 303.480 95.080 304.550 95.250 ;
        RECT 301.180 94.360 301.350 94.540 ;
        RECT 298.460 93.540 298.855 93.710 ;
        RECT 299.025 93.580 299.490 93.970 ;
        RECT 299.660 94.190 301.350 94.360 ;
        RECT 298.685 93.410 298.855 93.540 ;
        RECT 299.660 93.410 299.830 94.190 ;
        RECT 301.520 94.020 301.690 94.710 ;
        RECT 300.190 93.850 301.690 94.020 ;
        RECT 301.880 94.050 302.090 94.840 ;
        RECT 302.260 94.220 302.610 94.840 ;
        RECT 302.780 94.230 302.950 95.010 ;
        RECT 303.480 94.850 303.650 95.080 ;
        RECT 303.120 94.680 303.650 94.850 ;
        RECT 303.120 94.400 303.340 94.680 ;
        RECT 303.820 94.510 304.060 94.910 ;
        RECT 302.780 94.060 303.185 94.230 ;
        RECT 303.520 94.140 304.060 94.510 ;
        RECT 304.230 94.725 304.550 95.080 ;
        RECT 304.795 95.000 305.100 95.460 ;
        RECT 305.270 94.750 305.525 95.280 ;
        RECT 304.230 94.550 304.555 94.725 ;
        RECT 304.230 94.250 305.145 94.550 ;
        RECT 304.405 94.220 305.145 94.250 ;
        RECT 301.880 93.890 302.555 94.050 ;
        RECT 303.015 93.970 303.185 94.060 ;
        RECT 301.880 93.880 302.845 93.890 ;
        RECT 301.520 93.710 301.690 93.850 ;
        RECT 298.265 92.910 298.515 93.370 ;
        RECT 298.685 93.080 298.935 93.410 ;
        RECT 299.150 93.080 299.830 93.410 ;
        RECT 300.000 93.510 301.075 93.680 ;
        RECT 301.520 93.540 302.080 93.710 ;
        RECT 302.385 93.590 302.845 93.880 ;
        RECT 303.015 93.800 304.235 93.970 ;
        RECT 300.000 93.170 300.170 93.510 ;
        RECT 300.405 92.910 300.735 93.340 ;
        RECT 300.905 93.170 301.075 93.510 ;
        RECT 301.370 92.910 301.740 93.370 ;
        RECT 301.910 93.080 302.080 93.540 ;
        RECT 303.015 93.420 303.185 93.800 ;
        RECT 304.405 93.630 304.575 94.220 ;
        RECT 305.315 94.100 305.525 94.750 ;
        RECT 306.250 94.910 306.420 95.290 ;
        RECT 306.635 95.080 306.965 95.460 ;
        RECT 306.250 94.740 306.965 94.910 ;
        RECT 306.160 94.190 306.515 94.560 ;
        RECT 306.795 94.550 306.965 94.740 ;
        RECT 307.135 94.715 307.390 95.290 ;
        RECT 306.795 94.220 307.050 94.550 ;
        RECT 302.315 93.080 303.185 93.420 ;
        RECT 303.775 93.460 304.575 93.630 ;
        RECT 303.355 92.910 303.605 93.370 ;
        RECT 303.775 93.170 303.945 93.460 ;
        RECT 304.125 92.910 304.455 93.290 ;
        RECT 304.795 92.910 305.100 94.050 ;
        RECT 305.270 93.220 305.525 94.100 ;
        RECT 306.795 94.010 306.965 94.220 ;
        RECT 306.250 93.840 306.965 94.010 ;
        RECT 307.220 93.985 307.390 94.715 ;
        RECT 307.565 94.620 307.825 95.460 ;
        RECT 308.090 94.910 308.260 95.290 ;
        RECT 308.475 95.080 308.805 95.460 ;
        RECT 308.090 94.740 308.805 94.910 ;
        RECT 308.000 94.190 308.355 94.560 ;
        RECT 308.635 94.550 308.805 94.740 ;
        RECT 308.975 94.715 309.230 95.290 ;
        RECT 308.635 94.220 308.890 94.550 ;
        RECT 306.250 93.080 306.420 93.840 ;
        RECT 306.635 92.910 306.965 93.670 ;
        RECT 307.135 93.080 307.390 93.985 ;
        RECT 307.565 92.910 307.825 94.060 ;
        RECT 308.635 94.010 308.805 94.220 ;
        RECT 308.090 93.840 308.805 94.010 ;
        RECT 309.060 93.985 309.230 94.715 ;
        RECT 309.405 94.620 309.665 95.460 ;
        RECT 309.840 94.710 311.050 95.460 ;
        RECT 308.090 93.080 308.260 93.840 ;
        RECT 308.475 92.910 308.805 93.670 ;
        RECT 308.975 93.080 309.230 93.985 ;
        RECT 309.405 92.910 309.665 94.060 ;
        RECT 309.840 94.000 310.360 94.540 ;
        RECT 310.530 94.170 311.050 94.710 ;
        RECT 309.840 92.910 311.050 94.000 ;
        RECT 162.095 92.740 311.135 92.910 ;
        RECT 162.180 91.650 163.390 92.740 ;
        RECT 163.560 92.305 168.905 92.740 ;
        RECT 162.180 90.940 162.700 91.480 ;
        RECT 162.870 91.110 163.390 91.650 ;
        RECT 162.180 90.190 163.390 90.940 ;
        RECT 165.145 90.735 165.485 91.565 ;
        RECT 166.965 91.055 167.315 92.305 ;
        RECT 169.080 91.650 170.750 92.740 ;
        RECT 171.495 92.110 171.780 92.570 ;
        RECT 171.950 92.280 172.220 92.740 ;
        RECT 171.495 91.890 172.450 92.110 ;
        RECT 169.080 90.960 169.830 91.480 ;
        RECT 170.000 91.130 170.750 91.650 ;
        RECT 171.380 91.160 172.070 91.720 ;
        RECT 172.240 90.990 172.450 91.890 ;
        RECT 163.560 90.190 168.905 90.735 ;
        RECT 169.080 90.190 170.750 90.960 ;
        RECT 171.495 90.820 172.450 90.990 ;
        RECT 172.620 91.720 173.020 92.570 ;
        RECT 173.210 92.110 173.490 92.570 ;
        RECT 174.010 92.280 174.335 92.740 ;
        RECT 173.210 91.890 174.335 92.110 ;
        RECT 172.620 91.160 173.715 91.720 ;
        RECT 173.885 91.430 174.335 91.890 ;
        RECT 174.505 91.600 174.890 92.570 ;
        RECT 171.495 90.360 171.780 90.820 ;
        RECT 171.950 90.190 172.220 90.650 ;
        RECT 172.620 90.360 173.020 91.160 ;
        RECT 173.885 91.100 174.440 91.430 ;
        RECT 173.885 90.990 174.335 91.100 ;
        RECT 173.210 90.820 174.335 90.990 ;
        RECT 174.610 90.930 174.890 91.600 ;
        RECT 175.060 91.575 175.350 92.740 ;
        RECT 175.525 91.600 175.860 92.570 ;
        RECT 176.030 91.600 176.200 92.740 ;
        RECT 176.370 92.400 178.400 92.570 ;
        RECT 173.210 90.360 173.490 90.820 ;
        RECT 174.010 90.190 174.335 90.650 ;
        RECT 174.505 90.360 174.890 90.930 ;
        RECT 175.525 90.930 175.695 91.600 ;
        RECT 176.370 91.430 176.540 92.400 ;
        RECT 175.865 91.100 176.120 91.430 ;
        RECT 176.345 91.100 176.540 91.430 ;
        RECT 176.710 92.060 177.835 92.230 ;
        RECT 175.950 90.930 176.120 91.100 ;
        RECT 176.710 90.930 176.880 92.060 ;
        RECT 175.060 90.190 175.350 90.915 ;
        RECT 175.525 90.360 175.780 90.930 ;
        RECT 175.950 90.760 176.880 90.930 ;
        RECT 177.050 91.720 178.060 91.890 ;
        RECT 177.050 90.920 177.220 91.720 ;
        RECT 177.425 91.040 177.700 91.520 ;
        RECT 177.420 90.870 177.700 91.040 ;
        RECT 176.705 90.725 176.880 90.760 ;
        RECT 175.950 90.190 176.280 90.590 ;
        RECT 176.705 90.360 177.235 90.725 ;
        RECT 177.425 90.360 177.700 90.870 ;
        RECT 177.870 90.360 178.060 91.720 ;
        RECT 178.230 91.735 178.400 92.400 ;
        RECT 178.570 91.980 178.740 92.740 ;
        RECT 178.975 91.980 179.490 92.390 ;
        RECT 178.230 91.545 178.980 91.735 ;
        RECT 179.150 91.170 179.490 91.980 ;
        RECT 178.260 91.000 179.490 91.170 ;
        RECT 179.660 91.600 180.045 92.570 ;
        RECT 180.215 92.280 180.540 92.740 ;
        RECT 181.060 92.110 181.340 92.570 ;
        RECT 180.215 91.890 181.340 92.110 ;
        RECT 178.240 90.190 178.750 90.725 ;
        RECT 178.970 90.395 179.215 91.000 ;
        RECT 179.660 90.930 179.940 91.600 ;
        RECT 180.215 91.430 180.665 91.890 ;
        RECT 181.530 91.720 181.930 92.570 ;
        RECT 182.330 92.280 182.600 92.740 ;
        RECT 182.770 92.110 183.055 92.570 ;
        RECT 183.340 92.305 188.685 92.740 ;
        RECT 180.110 91.100 180.665 91.430 ;
        RECT 180.835 91.160 181.930 91.720 ;
        RECT 180.215 90.990 180.665 91.100 ;
        RECT 179.660 90.360 180.045 90.930 ;
        RECT 180.215 90.820 181.340 90.990 ;
        RECT 180.215 90.190 180.540 90.650 ;
        RECT 181.060 90.360 181.340 90.820 ;
        RECT 181.530 90.360 181.930 91.160 ;
        RECT 182.100 91.890 183.055 92.110 ;
        RECT 182.100 90.990 182.310 91.890 ;
        RECT 182.480 91.160 183.170 91.720 ;
        RECT 182.100 90.820 183.055 90.990 ;
        RECT 182.330 90.190 182.600 90.650 ;
        RECT 182.770 90.360 183.055 90.820 ;
        RECT 184.925 90.735 185.265 91.565 ;
        RECT 186.745 91.055 187.095 92.305 ;
        RECT 188.860 91.650 192.370 92.740 ;
        RECT 188.860 90.960 190.510 91.480 ;
        RECT 190.680 91.130 192.370 91.650 ;
        RECT 193.185 91.770 193.575 91.945 ;
        RECT 194.060 91.940 194.390 92.740 ;
        RECT 194.560 91.950 195.095 92.570 ;
        RECT 193.185 91.600 194.610 91.770 ;
        RECT 183.340 90.190 188.685 90.735 ;
        RECT 188.860 90.190 192.370 90.960 ;
        RECT 193.060 90.870 193.415 91.430 ;
        RECT 193.585 90.700 193.755 91.600 ;
        RECT 193.925 90.870 194.190 91.430 ;
        RECT 194.440 91.100 194.610 91.600 ;
        RECT 194.780 90.930 195.095 91.950 ;
        RECT 195.505 91.770 195.835 92.570 ;
        RECT 196.005 91.940 196.335 92.740 ;
        RECT 196.635 91.770 196.965 92.570 ;
        RECT 197.610 91.940 197.860 92.740 ;
        RECT 195.505 91.600 197.940 91.770 ;
        RECT 198.130 91.600 198.300 92.740 ;
        RECT 198.470 91.600 198.810 92.570 ;
        RECT 198.980 91.650 200.650 92.740 ;
        RECT 195.300 91.180 195.650 91.430 ;
        RECT 195.835 90.970 196.005 91.600 ;
        RECT 196.175 91.180 196.505 91.380 ;
        RECT 196.675 91.180 197.005 91.380 ;
        RECT 197.175 91.180 197.595 91.380 ;
        RECT 197.770 91.350 197.940 91.600 ;
        RECT 197.770 91.180 198.465 91.350 ;
        RECT 193.165 90.190 193.405 90.700 ;
        RECT 193.585 90.370 193.865 90.700 ;
        RECT 194.095 90.190 194.310 90.700 ;
        RECT 194.480 90.360 195.095 90.930 ;
        RECT 195.505 90.360 196.005 90.970 ;
        RECT 196.635 90.840 197.860 91.010 ;
        RECT 198.635 90.990 198.810 91.600 ;
        RECT 196.635 90.360 196.965 90.840 ;
        RECT 197.135 90.190 197.360 90.650 ;
        RECT 197.530 90.360 197.860 90.840 ;
        RECT 198.050 90.190 198.300 90.990 ;
        RECT 198.470 90.360 198.810 90.990 ;
        RECT 198.980 90.960 199.730 91.480 ;
        RECT 199.900 91.130 200.650 91.650 ;
        RECT 200.820 91.575 201.110 92.740 ;
        RECT 201.280 91.650 202.950 92.740 ;
        RECT 201.280 90.960 202.030 91.480 ;
        RECT 202.200 91.130 202.950 91.650 ;
        RECT 203.670 91.810 203.840 92.570 ;
        RECT 204.055 91.980 204.385 92.740 ;
        RECT 203.670 91.640 204.385 91.810 ;
        RECT 204.555 91.665 204.810 92.570 ;
        RECT 203.580 91.090 203.935 91.460 ;
        RECT 204.215 91.430 204.385 91.640 ;
        RECT 204.215 91.100 204.470 91.430 ;
        RECT 198.980 90.190 200.650 90.960 ;
        RECT 200.820 90.190 201.110 90.915 ;
        RECT 201.280 90.190 202.950 90.960 ;
        RECT 204.215 90.910 204.385 91.100 ;
        RECT 204.640 90.935 204.810 91.665 ;
        RECT 204.985 91.590 205.245 92.740 ;
        RECT 205.420 91.650 207.090 92.740 ;
        RECT 203.670 90.740 204.385 90.910 ;
        RECT 203.670 90.360 203.840 90.740 ;
        RECT 204.055 90.190 204.385 90.570 ;
        RECT 204.555 90.360 204.810 90.935 ;
        RECT 204.985 90.190 205.245 91.030 ;
        RECT 205.420 90.960 206.170 91.480 ;
        RECT 206.340 91.130 207.090 91.650 ;
        RECT 207.280 91.850 207.540 92.560 ;
        RECT 207.710 92.030 208.040 92.740 ;
        RECT 208.210 91.850 208.440 92.560 ;
        RECT 207.280 91.610 208.440 91.850 ;
        RECT 208.620 91.830 208.890 92.560 ;
        RECT 209.070 92.010 209.410 92.740 ;
        RECT 208.620 91.610 209.390 91.830 ;
        RECT 207.270 91.100 207.570 91.430 ;
        RECT 207.750 91.120 208.275 91.430 ;
        RECT 208.455 91.120 208.920 91.430 ;
        RECT 205.420 90.190 207.090 90.960 ;
        RECT 207.280 90.190 207.570 90.920 ;
        RECT 207.750 90.480 207.980 91.120 ;
        RECT 209.100 90.940 209.390 91.610 ;
        RECT 208.160 90.740 209.390 90.940 ;
        RECT 208.160 90.370 208.470 90.740 ;
        RECT 208.650 90.190 209.320 90.560 ;
        RECT 209.580 90.370 209.840 92.560 ;
        RECT 210.175 91.730 210.475 92.570 ;
        RECT 210.670 91.900 210.920 92.740 ;
        RECT 211.510 92.150 212.315 92.570 ;
        RECT 211.090 91.980 212.655 92.150 ;
        RECT 211.090 91.730 211.260 91.980 ;
        RECT 210.175 91.560 211.260 91.730 ;
        RECT 210.020 91.100 210.350 91.390 ;
        RECT 210.520 90.930 210.690 91.560 ;
        RECT 211.430 91.430 211.750 91.810 ;
        RECT 211.940 91.720 212.315 91.810 ;
        RECT 211.920 91.550 212.315 91.720 ;
        RECT 212.485 91.730 212.655 91.980 ;
        RECT 212.825 91.900 213.155 92.740 ;
        RECT 213.325 91.980 213.990 92.570 ;
        RECT 214.160 92.305 219.505 92.740 ;
        RECT 219.680 92.305 225.025 92.740 ;
        RECT 212.485 91.560 213.405 91.730 ;
        RECT 210.860 91.180 211.190 91.390 ;
        RECT 211.370 91.180 211.750 91.430 ;
        RECT 211.940 91.390 212.315 91.550 ;
        RECT 213.235 91.390 213.405 91.560 ;
        RECT 211.940 91.180 212.425 91.390 ;
        RECT 212.615 91.180 213.065 91.390 ;
        RECT 213.235 91.180 213.570 91.390 ;
        RECT 213.740 91.010 213.990 91.980 ;
        RECT 210.180 90.750 210.690 90.930 ;
        RECT 211.095 90.840 212.795 91.010 ;
        RECT 211.095 90.750 211.480 90.840 ;
        RECT 210.180 90.360 210.510 90.750 ;
        RECT 210.680 90.410 211.865 90.580 ;
        RECT 212.125 90.190 212.295 90.660 ;
        RECT 212.465 90.375 212.795 90.840 ;
        RECT 212.965 90.190 213.135 91.010 ;
        RECT 213.305 90.370 213.990 91.010 ;
        RECT 215.745 90.735 216.085 91.565 ;
        RECT 217.565 91.055 217.915 92.305 ;
        RECT 221.265 90.735 221.605 91.565 ;
        RECT 223.085 91.055 223.435 92.305 ;
        RECT 225.200 91.650 226.410 92.740 ;
        RECT 225.200 90.940 225.720 91.480 ;
        RECT 225.890 91.110 226.410 91.650 ;
        RECT 226.580 91.575 226.870 92.740 ;
        RECT 227.060 91.900 227.315 92.570 ;
        RECT 227.485 91.980 227.815 92.740 ;
        RECT 227.985 92.140 228.235 92.570 ;
        RECT 228.405 92.320 228.760 92.740 ;
        RECT 228.950 92.400 230.120 92.570 ;
        RECT 228.950 92.360 229.280 92.400 ;
        RECT 229.390 92.140 229.620 92.230 ;
        RECT 227.985 91.900 229.620 92.140 ;
        RECT 229.790 91.900 230.120 92.400 ;
        RECT 214.160 90.190 219.505 90.735 ;
        RECT 219.680 90.190 225.025 90.735 ;
        RECT 225.200 90.190 226.410 90.940 ;
        RECT 226.580 90.190 226.870 90.915 ;
        RECT 227.060 90.770 227.230 91.900 ;
        RECT 230.290 91.730 230.460 92.570 ;
        RECT 227.400 91.560 230.460 91.730 ;
        RECT 230.720 91.890 230.980 92.570 ;
        RECT 231.150 91.960 231.400 92.740 ;
        RECT 231.650 92.190 231.900 92.570 ;
        RECT 232.070 92.360 232.425 92.740 ;
        RECT 233.430 92.350 233.765 92.570 ;
        RECT 233.030 92.190 233.260 92.230 ;
        RECT 231.650 91.990 233.260 92.190 ;
        RECT 231.650 91.980 232.485 91.990 ;
        RECT 233.075 91.900 233.260 91.990 ;
        RECT 227.400 91.010 227.570 91.560 ;
        RECT 227.800 91.180 228.165 91.380 ;
        RECT 228.335 91.180 228.665 91.380 ;
        RECT 227.400 90.840 228.200 91.010 ;
        RECT 227.060 90.700 227.245 90.770 ;
        RECT 227.060 90.690 227.270 90.700 ;
        RECT 227.060 90.360 227.315 90.690 ;
        RECT 227.530 90.190 227.860 90.670 ;
        RECT 228.030 90.610 228.200 90.840 ;
        RECT 228.380 90.780 228.665 91.180 ;
        RECT 228.935 91.180 229.410 91.380 ;
        RECT 229.580 91.180 230.025 91.380 ;
        RECT 230.195 91.180 230.545 91.390 ;
        RECT 228.935 90.780 229.215 91.180 ;
        RECT 229.395 90.840 230.460 91.010 ;
        RECT 229.395 90.610 229.565 90.840 ;
        RECT 228.030 90.360 229.565 90.610 ;
        RECT 229.790 90.190 230.120 90.670 ;
        RECT 230.290 90.360 230.460 90.840 ;
        RECT 230.720 90.700 230.890 91.890 ;
        RECT 232.590 91.790 232.920 91.820 ;
        RECT 231.120 91.730 232.920 91.790 ;
        RECT 233.510 91.730 233.765 92.350 ;
        RECT 233.940 92.305 239.285 92.740 ;
        RECT 231.060 91.620 233.765 91.730 ;
        RECT 231.060 91.585 231.260 91.620 ;
        RECT 231.060 91.010 231.230 91.585 ;
        RECT 232.590 91.560 233.765 91.620 ;
        RECT 231.460 91.145 231.870 91.450 ;
        RECT 232.040 91.180 232.370 91.390 ;
        RECT 231.060 90.890 231.330 91.010 ;
        RECT 231.060 90.845 231.905 90.890 ;
        RECT 231.150 90.720 231.905 90.845 ;
        RECT 232.160 90.780 232.370 91.180 ;
        RECT 232.615 91.180 233.090 91.390 ;
        RECT 233.280 91.180 233.770 91.380 ;
        RECT 232.615 90.780 232.835 91.180 ;
        RECT 230.720 90.690 230.950 90.700 ;
        RECT 230.720 90.360 230.980 90.690 ;
        RECT 231.735 90.570 231.905 90.720 ;
        RECT 231.150 90.190 231.480 90.550 ;
        RECT 231.735 90.360 233.035 90.570 ;
        RECT 233.310 90.190 233.765 90.955 ;
        RECT 235.525 90.735 235.865 91.565 ;
        RECT 237.345 91.055 237.695 92.305 ;
        RECT 239.460 91.650 241.130 92.740 ;
        RECT 239.460 90.960 240.210 91.480 ;
        RECT 240.380 91.130 241.130 91.650 ;
        RECT 241.305 92.020 241.640 92.530 ;
        RECT 233.940 90.190 239.285 90.735 ;
        RECT 239.460 90.190 241.130 90.960 ;
        RECT 241.305 90.665 241.560 92.020 ;
        RECT 241.890 91.940 242.220 92.740 ;
        RECT 242.465 92.150 242.750 92.570 ;
        RECT 243.005 92.320 243.335 92.740 ;
        RECT 243.560 92.400 244.720 92.570 ;
        RECT 243.560 92.150 243.890 92.400 ;
        RECT 242.465 91.980 243.890 92.150 ;
        RECT 244.120 91.770 244.290 92.230 ;
        RECT 244.550 91.900 244.720 92.400 ;
        RECT 245.000 91.900 245.255 92.570 ;
        RECT 245.425 91.980 245.755 92.740 ;
        RECT 245.925 92.140 246.175 92.570 ;
        RECT 246.345 92.320 246.700 92.740 ;
        RECT 246.890 92.400 248.060 92.570 ;
        RECT 246.890 92.360 247.220 92.400 ;
        RECT 247.330 92.140 247.560 92.230 ;
        RECT 245.925 91.900 247.560 92.140 ;
        RECT 247.730 91.900 248.060 92.400 ;
        RECT 241.920 91.600 244.290 91.770 ;
        RECT 245.000 91.890 245.210 91.900 ;
        RECT 241.920 91.430 242.090 91.600 ;
        RECT 244.540 91.550 244.750 91.720 ;
        RECT 244.540 91.430 244.745 91.550 ;
        RECT 241.785 91.100 242.090 91.430 ;
        RECT 242.285 91.380 242.535 91.430 ;
        RECT 242.745 91.380 243.015 91.430 ;
        RECT 242.280 91.210 242.535 91.380 ;
        RECT 242.740 91.210 243.015 91.380 ;
        RECT 242.285 91.100 242.535 91.210 ;
        RECT 241.920 90.930 242.090 91.100 ;
        RECT 241.920 90.760 242.480 90.930 ;
        RECT 242.745 90.770 243.015 91.210 ;
        RECT 243.205 91.040 243.495 91.430 ;
        RECT 243.200 90.870 243.495 91.040 ;
        RECT 243.205 90.770 243.495 90.870 ;
        RECT 243.665 90.765 244.085 91.430 ;
        RECT 244.395 91.100 244.745 91.430 ;
        RECT 241.305 90.405 241.640 90.665 ;
        RECT 242.310 90.590 242.480 90.760 ;
        RECT 241.810 90.190 242.140 90.590 ;
        RECT 242.310 90.420 243.925 90.590 ;
        RECT 244.470 90.190 244.800 90.910 ;
        RECT 245.000 90.770 245.170 91.890 ;
        RECT 248.230 91.730 248.400 92.570 ;
        RECT 245.340 91.560 248.400 91.730 ;
        RECT 248.660 91.650 252.170 92.740 ;
        RECT 245.340 91.010 245.510 91.560 ;
        RECT 245.740 91.180 246.105 91.380 ;
        RECT 246.275 91.180 246.605 91.380 ;
        RECT 245.340 90.840 246.140 91.010 ;
        RECT 245.000 90.690 245.185 90.770 ;
        RECT 245.000 90.360 245.255 90.690 ;
        RECT 245.470 90.190 245.800 90.670 ;
        RECT 245.970 90.610 246.140 90.840 ;
        RECT 246.320 90.780 246.605 91.180 ;
        RECT 246.875 91.180 247.350 91.380 ;
        RECT 247.520 91.180 247.965 91.380 ;
        RECT 248.135 91.180 248.485 91.390 ;
        RECT 246.875 90.780 247.155 91.180 ;
        RECT 247.335 90.840 248.400 91.010 ;
        RECT 247.335 90.610 247.505 90.840 ;
        RECT 245.970 90.360 247.505 90.610 ;
        RECT 247.730 90.190 248.060 90.670 ;
        RECT 248.230 90.360 248.400 90.840 ;
        RECT 248.660 90.960 250.310 91.480 ;
        RECT 250.480 91.130 252.170 91.650 ;
        RECT 252.340 91.575 252.630 92.740 ;
        RECT 252.800 92.305 258.145 92.740 ;
        RECT 248.660 90.190 252.170 90.960 ;
        RECT 252.340 90.190 252.630 90.915 ;
        RECT 254.385 90.735 254.725 91.565 ;
        RECT 256.205 91.055 256.555 92.305 ;
        RECT 258.320 91.650 259.990 92.740 ;
        RECT 258.320 90.960 259.070 91.480 ;
        RECT 259.240 91.130 259.990 91.650 ;
        RECT 260.625 92.350 260.960 92.570 ;
        RECT 261.965 92.360 262.320 92.740 ;
        RECT 260.625 91.730 260.880 92.350 ;
        RECT 261.130 92.190 261.360 92.230 ;
        RECT 262.490 92.190 262.740 92.570 ;
        RECT 261.130 91.990 262.740 92.190 ;
        RECT 261.130 91.900 261.315 91.990 ;
        RECT 261.905 91.980 262.740 91.990 ;
        RECT 262.990 91.960 263.240 92.740 ;
        RECT 263.410 91.890 263.670 92.570 ;
        RECT 261.470 91.790 261.800 91.820 ;
        RECT 261.470 91.730 263.270 91.790 ;
        RECT 260.625 91.620 263.330 91.730 ;
        RECT 260.625 91.560 261.800 91.620 ;
        RECT 263.130 91.585 263.330 91.620 ;
        RECT 260.620 91.180 261.110 91.380 ;
        RECT 261.300 91.180 261.775 91.390 ;
        RECT 252.800 90.190 258.145 90.735 ;
        RECT 258.320 90.190 259.990 90.960 ;
        RECT 260.625 90.190 261.080 90.955 ;
        RECT 261.555 90.780 261.775 91.180 ;
        RECT 262.020 91.180 262.350 91.390 ;
        RECT 262.020 90.780 262.230 91.180 ;
        RECT 262.520 91.145 262.930 91.450 ;
        RECT 263.160 91.010 263.330 91.585 ;
        RECT 263.060 90.890 263.330 91.010 ;
        RECT 262.485 90.845 263.330 90.890 ;
        RECT 262.485 90.720 263.240 90.845 ;
        RECT 262.485 90.570 262.655 90.720 ;
        RECT 263.500 90.690 263.670 91.890 ;
        RECT 263.845 92.350 264.180 92.570 ;
        RECT 265.185 92.360 265.540 92.740 ;
        RECT 263.845 91.730 264.100 92.350 ;
        RECT 264.350 92.190 264.580 92.230 ;
        RECT 265.710 92.190 265.960 92.570 ;
        RECT 264.350 91.990 265.960 92.190 ;
        RECT 264.350 91.900 264.535 91.990 ;
        RECT 265.125 91.980 265.960 91.990 ;
        RECT 266.210 91.960 266.460 92.740 ;
        RECT 266.630 91.890 266.890 92.570 ;
        RECT 267.060 92.230 268.250 92.520 ;
        RECT 264.690 91.790 265.020 91.820 ;
        RECT 264.690 91.730 266.490 91.790 ;
        RECT 263.845 91.620 266.550 91.730 ;
        RECT 263.845 91.560 265.020 91.620 ;
        RECT 266.350 91.585 266.550 91.620 ;
        RECT 263.840 91.180 264.330 91.380 ;
        RECT 264.520 91.180 264.995 91.390 ;
        RECT 261.355 90.360 262.655 90.570 ;
        RECT 262.910 90.190 263.240 90.550 ;
        RECT 263.410 90.360 263.670 90.690 ;
        RECT 263.845 90.190 264.300 90.955 ;
        RECT 264.775 90.780 264.995 91.180 ;
        RECT 265.240 91.180 265.570 91.390 ;
        RECT 265.240 90.780 265.450 91.180 ;
        RECT 265.740 91.145 266.150 91.450 ;
        RECT 266.380 91.010 266.550 91.585 ;
        RECT 266.280 90.890 266.550 91.010 ;
        RECT 265.705 90.845 266.550 90.890 ;
        RECT 265.705 90.720 266.460 90.845 ;
        RECT 265.705 90.570 265.875 90.720 ;
        RECT 266.720 90.700 266.890 91.890 ;
        RECT 267.080 91.890 268.250 92.060 ;
        RECT 268.420 91.940 268.700 92.740 ;
        RECT 267.080 91.600 267.405 91.890 ;
        RECT 268.080 91.770 268.250 91.890 ;
        RECT 267.575 91.430 267.770 91.720 ;
        RECT 268.080 91.600 268.740 91.770 ;
        RECT 268.910 91.600 269.185 92.570 ;
        RECT 269.360 92.305 274.705 92.740 ;
        RECT 268.570 91.430 268.740 91.600 ;
        RECT 267.060 91.100 267.405 91.430 ;
        RECT 267.575 91.100 268.400 91.430 ;
        RECT 268.570 91.100 268.845 91.430 ;
        RECT 268.570 90.930 268.740 91.100 ;
        RECT 266.660 90.690 266.890 90.700 ;
        RECT 264.575 90.360 265.875 90.570 ;
        RECT 266.130 90.190 266.460 90.550 ;
        RECT 266.630 90.360 266.890 90.690 ;
        RECT 267.075 90.760 268.740 90.930 ;
        RECT 269.015 90.865 269.185 91.600 ;
        RECT 267.075 90.410 267.330 90.760 ;
        RECT 267.500 90.190 267.830 90.590 ;
        RECT 268.000 90.410 268.170 90.760 ;
        RECT 268.340 90.190 268.720 90.590 ;
        RECT 268.910 90.520 269.185 90.865 ;
        RECT 270.945 90.735 271.285 91.565 ;
        RECT 272.765 91.055 273.115 92.305 ;
        RECT 274.880 91.650 277.470 92.740 ;
        RECT 274.880 90.960 276.090 91.480 ;
        RECT 276.260 91.130 277.470 91.650 ;
        RECT 278.100 91.575 278.390 92.740 ;
        RECT 278.565 92.020 278.900 92.530 ;
        RECT 269.360 90.190 274.705 90.735 ;
        RECT 274.880 90.190 277.470 90.960 ;
        RECT 278.100 90.190 278.390 90.915 ;
        RECT 278.565 90.665 278.820 92.020 ;
        RECT 279.150 91.940 279.480 92.740 ;
        RECT 279.725 92.150 280.010 92.570 ;
        RECT 280.265 92.320 280.595 92.740 ;
        RECT 280.820 92.400 281.980 92.570 ;
        RECT 280.820 92.150 281.150 92.400 ;
        RECT 279.725 91.980 281.150 92.150 ;
        RECT 281.380 91.770 281.550 92.230 ;
        RECT 281.810 91.900 281.980 92.400 ;
        RECT 282.250 92.020 282.580 92.740 ;
        RECT 279.180 91.600 281.550 91.770 ;
        RECT 279.180 91.430 279.350 91.600 ;
        RECT 281.800 91.550 282.010 91.720 ;
        RECT 281.800 91.430 282.005 91.550 ;
        RECT 279.045 91.100 279.350 91.430 ;
        RECT 279.545 91.380 279.795 91.430 ;
        RECT 279.540 91.210 279.795 91.380 ;
        RECT 279.545 91.100 279.795 91.210 ;
        RECT 279.180 90.930 279.350 91.100 ;
        RECT 280.005 91.040 280.275 91.430 ;
        RECT 280.465 91.040 280.755 91.430 ;
        RECT 279.180 90.760 279.740 90.930 ;
        RECT 280.000 90.870 280.275 91.040 ;
        RECT 280.460 90.870 280.755 91.040 ;
        RECT 280.005 90.770 280.275 90.870 ;
        RECT 280.465 90.770 280.755 90.870 ;
        RECT 280.925 90.765 281.345 91.430 ;
        RECT 281.655 91.100 282.005 91.430 ;
        RECT 282.240 91.380 282.470 91.720 ;
        RECT 282.760 91.380 282.975 92.495 ;
        RECT 283.170 91.795 283.500 92.570 ;
        RECT 283.670 91.965 284.380 92.740 ;
        RECT 283.170 91.580 284.320 91.795 ;
        RECT 282.240 91.180 282.570 91.380 ;
        RECT 282.760 91.200 283.210 91.380 ;
        RECT 282.880 91.180 283.210 91.200 ;
        RECT 283.380 91.180 283.850 91.410 ;
        RECT 284.035 91.010 284.320 91.580 ;
        RECT 284.550 91.135 284.830 92.570 ;
        RECT 285.000 91.650 288.510 92.740 ;
        RECT 288.680 91.650 289.890 92.740 ;
        RECT 278.565 90.405 278.900 90.665 ;
        RECT 279.570 90.590 279.740 90.760 ;
        RECT 279.070 90.190 279.400 90.590 ;
        RECT 279.570 90.420 281.185 90.590 ;
        RECT 281.730 90.190 282.060 90.910 ;
        RECT 282.240 90.820 283.420 91.010 ;
        RECT 282.240 90.360 282.580 90.820 ;
        RECT 283.090 90.740 283.420 90.820 ;
        RECT 283.610 90.820 284.320 91.010 ;
        RECT 283.610 90.680 283.910 90.820 ;
        RECT 283.595 90.670 283.910 90.680 ;
        RECT 283.585 90.660 283.910 90.670 ;
        RECT 283.575 90.655 283.910 90.660 ;
        RECT 282.750 90.190 282.920 90.650 ;
        RECT 283.570 90.645 283.910 90.655 ;
        RECT 283.565 90.640 283.910 90.645 ;
        RECT 283.560 90.630 283.910 90.640 ;
        RECT 283.555 90.625 283.910 90.630 ;
        RECT 283.550 90.360 283.910 90.625 ;
        RECT 284.150 90.190 284.320 90.650 ;
        RECT 284.490 90.360 284.830 91.135 ;
        RECT 285.000 90.960 286.650 91.480 ;
        RECT 286.820 91.130 288.510 91.650 ;
        RECT 285.000 90.190 288.510 90.960 ;
        RECT 288.680 90.940 289.200 91.480 ;
        RECT 289.370 91.110 289.890 91.650 ;
        RECT 290.065 91.600 290.400 92.570 ;
        RECT 290.570 91.600 290.740 92.740 ;
        RECT 290.910 92.400 292.940 92.570 ;
        RECT 288.680 90.190 289.890 90.940 ;
        RECT 290.065 90.930 290.235 91.600 ;
        RECT 290.910 91.430 291.080 92.400 ;
        RECT 290.405 91.100 290.660 91.430 ;
        RECT 290.885 91.100 291.080 91.430 ;
        RECT 291.250 92.060 292.375 92.230 ;
        RECT 290.490 90.930 290.660 91.100 ;
        RECT 291.250 90.930 291.420 92.060 ;
        RECT 290.065 90.360 290.320 90.930 ;
        RECT 290.490 90.760 291.420 90.930 ;
        RECT 291.590 91.720 292.600 91.890 ;
        RECT 291.590 90.920 291.760 91.720 ;
        RECT 291.245 90.725 291.420 90.760 ;
        RECT 290.490 90.190 290.820 90.590 ;
        RECT 291.245 90.360 291.775 90.725 ;
        RECT 291.965 90.700 292.240 91.520 ;
        RECT 291.960 90.530 292.240 90.700 ;
        RECT 291.965 90.360 292.240 90.530 ;
        RECT 292.410 90.360 292.600 91.720 ;
        RECT 292.770 91.735 292.940 92.400 ;
        RECT 293.110 91.980 293.280 92.740 ;
        RECT 293.515 91.980 294.030 92.390 ;
        RECT 292.770 91.545 293.520 91.735 ;
        RECT 293.690 91.170 294.030 91.980 ;
        RECT 294.665 92.070 294.920 92.570 ;
        RECT 295.090 92.240 295.420 92.740 ;
        RECT 294.665 91.900 295.415 92.070 ;
        RECT 292.800 91.000 294.030 91.170 ;
        RECT 294.665 91.080 295.015 91.730 ;
        RECT 292.780 90.190 293.290 90.725 ;
        RECT 293.510 90.395 293.755 91.000 ;
        RECT 295.185 90.910 295.415 91.900 ;
        RECT 294.665 90.740 295.415 90.910 ;
        RECT 294.665 90.450 294.920 90.740 ;
        RECT 295.090 90.190 295.420 90.570 ;
        RECT 295.590 90.450 295.760 92.570 ;
        RECT 295.930 91.770 296.255 92.555 ;
        RECT 296.425 92.280 296.675 92.740 ;
        RECT 296.845 92.240 297.095 92.570 ;
        RECT 297.310 92.240 297.990 92.570 ;
        RECT 296.845 92.110 297.015 92.240 ;
        RECT 296.620 91.940 297.015 92.110 ;
        RECT 295.990 90.720 296.450 91.770 ;
        RECT 296.620 90.580 296.790 91.940 ;
        RECT 297.185 91.680 297.650 92.070 ;
        RECT 296.960 90.870 297.310 91.490 ;
        RECT 297.480 91.090 297.650 91.680 ;
        RECT 297.820 91.460 297.990 92.240 ;
        RECT 298.160 92.140 298.330 92.480 ;
        RECT 298.565 92.310 298.895 92.740 ;
        RECT 299.065 92.140 299.235 92.480 ;
        RECT 299.530 92.280 299.900 92.740 ;
        RECT 298.160 91.970 299.235 92.140 ;
        RECT 300.070 92.110 300.240 92.570 ;
        RECT 300.475 92.230 301.345 92.570 ;
        RECT 301.515 92.280 301.765 92.740 ;
        RECT 299.680 91.940 300.240 92.110 ;
        RECT 299.680 91.800 299.850 91.940 ;
        RECT 298.350 91.630 299.850 91.800 ;
        RECT 300.545 91.770 301.005 92.060 ;
        RECT 297.820 91.290 299.510 91.460 ;
        RECT 297.480 90.870 297.835 91.090 ;
        RECT 298.005 90.580 298.175 91.290 ;
        RECT 298.380 90.870 299.170 91.120 ;
        RECT 299.340 91.110 299.510 91.290 ;
        RECT 299.680 90.940 299.850 91.630 ;
        RECT 296.120 90.190 296.450 90.550 ;
        RECT 296.620 90.410 297.115 90.580 ;
        RECT 297.320 90.410 298.175 90.580 ;
        RECT 299.050 90.190 299.380 90.650 ;
        RECT 299.590 90.550 299.850 90.940 ;
        RECT 300.040 91.760 301.005 91.770 ;
        RECT 301.175 91.850 301.345 92.230 ;
        RECT 301.935 92.190 302.105 92.480 ;
        RECT 302.285 92.360 302.615 92.740 ;
        RECT 301.935 92.020 302.735 92.190 ;
        RECT 300.040 91.600 300.715 91.760 ;
        RECT 301.175 91.680 302.395 91.850 ;
        RECT 300.040 90.810 300.250 91.600 ;
        RECT 301.175 91.590 301.345 91.680 ;
        RECT 300.420 90.810 300.770 91.430 ;
        RECT 300.940 91.420 301.345 91.590 ;
        RECT 300.940 90.640 301.110 91.420 ;
        RECT 301.280 90.970 301.500 91.250 ;
        RECT 301.680 91.140 302.220 91.510 ;
        RECT 302.565 91.430 302.735 92.020 ;
        RECT 302.955 91.600 303.260 92.740 ;
        RECT 303.430 91.550 303.685 92.430 ;
        RECT 303.860 91.575 304.150 92.740 ;
        RECT 304.320 91.650 307.830 92.740 ;
        RECT 302.565 91.400 303.305 91.430 ;
        RECT 301.280 90.800 301.810 90.970 ;
        RECT 299.590 90.380 299.940 90.550 ;
        RECT 300.160 90.360 301.110 90.640 ;
        RECT 301.280 90.190 301.470 90.630 ;
        RECT 301.640 90.570 301.810 90.800 ;
        RECT 301.980 90.740 302.220 91.140 ;
        RECT 302.390 91.100 303.305 91.400 ;
        RECT 302.390 90.925 302.715 91.100 ;
        RECT 302.390 90.570 302.710 90.925 ;
        RECT 303.475 90.900 303.685 91.550 ;
        RECT 304.320 90.960 305.970 91.480 ;
        RECT 306.140 91.130 307.830 91.650 ;
        RECT 308.090 91.810 308.260 92.570 ;
        RECT 308.475 91.980 308.805 92.740 ;
        RECT 308.090 91.640 308.805 91.810 ;
        RECT 308.975 91.665 309.230 92.570 ;
        RECT 308.000 91.090 308.355 91.460 ;
        RECT 308.635 91.430 308.805 91.640 ;
        RECT 308.635 91.100 308.890 91.430 ;
        RECT 301.640 90.400 302.710 90.570 ;
        RECT 302.955 90.190 303.260 90.650 ;
        RECT 303.430 90.370 303.685 90.900 ;
        RECT 303.860 90.190 304.150 90.915 ;
        RECT 304.320 90.190 307.830 90.960 ;
        RECT 308.635 90.910 308.805 91.100 ;
        RECT 309.060 90.935 309.230 91.665 ;
        RECT 309.405 91.590 309.665 92.740 ;
        RECT 309.840 91.650 311.050 92.740 ;
        RECT 309.840 91.110 310.360 91.650 ;
        RECT 308.090 90.740 308.805 90.910 ;
        RECT 308.090 90.360 308.260 90.740 ;
        RECT 308.475 90.190 308.805 90.570 ;
        RECT 308.975 90.360 309.230 90.935 ;
        RECT 309.405 90.190 309.665 91.030 ;
        RECT 310.530 90.940 311.050 91.480 ;
        RECT 309.840 90.190 311.050 90.940 ;
        RECT 162.095 90.020 311.135 90.190 ;
        RECT 162.180 89.270 163.390 90.020 ;
        RECT 163.560 89.475 168.905 90.020 ;
        RECT 162.180 88.730 162.700 89.270 ;
        RECT 162.870 88.560 163.390 89.100 ;
        RECT 165.145 88.645 165.485 89.475 ;
        RECT 169.085 89.310 169.340 89.840 ;
        RECT 169.510 89.560 169.815 90.020 ;
        RECT 170.060 89.640 171.130 89.810 ;
        RECT 162.180 87.470 163.390 88.560 ;
        RECT 166.965 87.905 167.315 89.155 ;
        RECT 169.085 88.660 169.295 89.310 ;
        RECT 170.060 89.285 170.380 89.640 ;
        RECT 170.055 89.110 170.380 89.285 ;
        RECT 169.465 88.810 170.380 89.110 ;
        RECT 170.550 89.070 170.790 89.470 ;
        RECT 170.960 89.410 171.130 89.640 ;
        RECT 171.300 89.580 171.490 90.020 ;
        RECT 171.660 89.570 172.610 89.850 ;
        RECT 172.830 89.660 173.180 89.830 ;
        RECT 170.960 89.240 171.490 89.410 ;
        RECT 169.465 88.780 170.205 88.810 ;
        RECT 163.560 87.470 168.905 87.905 ;
        RECT 169.085 87.780 169.340 88.660 ;
        RECT 169.510 87.470 169.815 88.610 ;
        RECT 170.035 88.190 170.205 88.780 ;
        RECT 170.550 88.700 171.090 89.070 ;
        RECT 171.270 88.960 171.490 89.240 ;
        RECT 171.660 88.790 171.830 89.570 ;
        RECT 171.425 88.620 171.830 88.790 ;
        RECT 172.000 88.780 172.350 89.400 ;
        RECT 171.425 88.530 171.595 88.620 ;
        RECT 172.520 88.610 172.730 89.400 ;
        RECT 170.375 88.360 171.595 88.530 ;
        RECT 172.055 88.450 172.730 88.610 ;
        RECT 170.035 88.020 170.835 88.190 ;
        RECT 170.155 87.470 170.485 87.850 ;
        RECT 170.665 87.730 170.835 88.020 ;
        RECT 171.425 87.980 171.595 88.360 ;
        RECT 171.765 88.440 172.730 88.450 ;
        RECT 172.920 89.270 173.180 89.660 ;
        RECT 173.390 89.560 173.720 90.020 ;
        RECT 174.595 89.630 175.450 89.800 ;
        RECT 175.655 89.630 176.150 89.800 ;
        RECT 176.320 89.660 176.650 90.020 ;
        RECT 172.920 88.580 173.090 89.270 ;
        RECT 173.260 88.920 173.430 89.100 ;
        RECT 173.600 89.090 174.390 89.340 ;
        RECT 174.595 88.920 174.765 89.630 ;
        RECT 174.935 89.120 175.290 89.340 ;
        RECT 173.260 88.750 174.950 88.920 ;
        RECT 171.765 88.150 172.225 88.440 ;
        RECT 172.920 88.410 174.420 88.580 ;
        RECT 172.920 88.270 173.090 88.410 ;
        RECT 172.530 88.100 173.090 88.270 ;
        RECT 171.005 87.470 171.255 87.930 ;
        RECT 171.425 87.640 172.295 87.980 ;
        RECT 172.530 87.640 172.700 88.100 ;
        RECT 173.535 88.070 174.610 88.240 ;
        RECT 172.870 87.470 173.240 87.930 ;
        RECT 173.535 87.730 173.705 88.070 ;
        RECT 173.875 87.470 174.205 87.900 ;
        RECT 174.440 87.730 174.610 88.070 ;
        RECT 174.780 87.970 174.950 88.750 ;
        RECT 175.120 88.530 175.290 89.120 ;
        RECT 175.460 88.720 175.810 89.340 ;
        RECT 175.120 88.140 175.585 88.530 ;
        RECT 175.980 88.270 176.150 89.630 ;
        RECT 176.320 88.440 176.780 89.490 ;
        RECT 175.755 88.100 176.150 88.270 ;
        RECT 175.755 87.970 175.925 88.100 ;
        RECT 174.780 87.640 175.460 87.970 ;
        RECT 175.675 87.640 175.925 87.970 ;
        RECT 176.095 87.470 176.345 87.930 ;
        RECT 176.515 87.655 176.840 88.440 ;
        RECT 177.010 87.640 177.180 89.760 ;
        RECT 177.350 89.640 177.680 90.020 ;
        RECT 177.850 89.470 178.105 89.760 ;
        RECT 177.355 89.300 178.105 89.470 ;
        RECT 177.355 88.310 177.585 89.300 ;
        RECT 178.285 89.280 178.540 89.850 ;
        RECT 178.710 89.620 179.040 90.020 ;
        RECT 179.465 89.485 179.995 89.850 ;
        RECT 180.185 89.680 180.460 89.850 ;
        RECT 180.180 89.510 180.460 89.680 ;
        RECT 179.465 89.450 179.640 89.485 ;
        RECT 178.710 89.280 179.640 89.450 ;
        RECT 177.755 88.480 178.105 89.130 ;
        RECT 178.285 88.610 178.455 89.280 ;
        RECT 178.710 89.110 178.880 89.280 ;
        RECT 178.625 88.780 178.880 89.110 ;
        RECT 179.105 88.780 179.300 89.110 ;
        RECT 177.355 88.140 178.105 88.310 ;
        RECT 177.350 87.470 177.680 87.970 ;
        RECT 177.850 87.640 178.105 88.140 ;
        RECT 178.285 87.640 178.620 88.610 ;
        RECT 178.790 87.470 178.960 88.610 ;
        RECT 179.130 87.810 179.300 88.780 ;
        RECT 179.470 88.150 179.640 89.280 ;
        RECT 179.810 88.490 179.980 89.290 ;
        RECT 180.185 88.690 180.460 89.510 ;
        RECT 180.630 88.490 180.820 89.850 ;
        RECT 181.000 89.485 181.510 90.020 ;
        RECT 181.730 89.210 181.975 89.815 ;
        RECT 182.420 89.475 187.765 90.020 ;
        RECT 181.020 89.040 182.250 89.210 ;
        RECT 179.810 88.320 180.820 88.490 ;
        RECT 180.990 88.475 181.740 88.665 ;
        RECT 179.470 87.980 180.595 88.150 ;
        RECT 180.990 87.810 181.160 88.475 ;
        RECT 181.910 88.230 182.250 89.040 ;
        RECT 184.005 88.645 184.345 89.475 ;
        RECT 187.940 89.295 188.230 90.020 ;
        RECT 188.400 89.220 188.690 90.020 ;
        RECT 188.860 89.560 189.410 89.850 ;
        RECT 189.580 89.560 189.830 90.020 ;
        RECT 179.130 87.640 181.160 87.810 ;
        RECT 181.330 87.470 181.500 88.230 ;
        RECT 181.735 87.820 182.250 88.230 ;
        RECT 185.825 87.905 186.175 89.155 ;
        RECT 182.420 87.470 187.765 87.905 ;
        RECT 187.940 87.470 188.230 88.635 ;
        RECT 188.400 87.470 188.690 88.610 ;
        RECT 188.860 88.190 189.110 89.560 ;
        RECT 190.460 89.390 190.790 89.750 ;
        RECT 191.160 89.475 196.505 90.020 ;
        RECT 196.680 89.475 202.025 90.020 ;
        RECT 202.365 89.510 202.605 90.020 ;
        RECT 202.785 89.510 203.065 89.840 ;
        RECT 203.295 89.510 203.510 90.020 ;
        RECT 189.400 89.200 190.790 89.390 ;
        RECT 189.400 89.110 189.570 89.200 ;
        RECT 189.280 88.780 189.570 89.110 ;
        RECT 189.740 88.780 190.070 89.030 ;
        RECT 190.300 88.780 190.990 89.030 ;
        RECT 189.400 88.530 189.570 88.780 ;
        RECT 189.400 88.360 190.340 88.530 ;
        RECT 188.860 87.640 189.310 88.190 ;
        RECT 189.500 87.470 189.830 88.190 ;
        RECT 190.040 87.810 190.340 88.360 ;
        RECT 190.675 88.340 190.990 88.780 ;
        RECT 192.745 88.645 193.085 89.475 ;
        RECT 190.510 87.470 190.790 88.140 ;
        RECT 194.565 87.905 194.915 89.155 ;
        RECT 198.265 88.645 198.605 89.475 ;
        RECT 200.085 87.905 200.435 89.155 ;
        RECT 202.260 88.780 202.615 89.340 ;
        RECT 202.785 88.610 202.955 89.510 ;
        RECT 203.125 88.780 203.390 89.340 ;
        RECT 203.680 89.280 204.295 89.850 ;
        RECT 204.520 89.290 204.810 90.020 ;
        RECT 203.640 88.610 203.810 89.110 ;
        RECT 202.385 88.440 203.810 88.610 ;
        RECT 202.385 88.265 202.775 88.440 ;
        RECT 191.160 87.470 196.505 87.905 ;
        RECT 196.680 87.470 202.025 87.905 ;
        RECT 203.260 87.470 203.590 88.270 ;
        RECT 203.980 88.260 204.295 89.280 ;
        RECT 204.510 88.780 204.810 89.110 ;
        RECT 204.990 89.090 205.220 89.730 ;
        RECT 205.400 89.470 205.710 89.840 ;
        RECT 205.890 89.650 206.560 90.020 ;
        RECT 205.400 89.270 206.630 89.470 ;
        RECT 204.990 88.780 205.515 89.090 ;
        RECT 205.695 88.780 206.160 89.090 ;
        RECT 206.340 88.600 206.630 89.270 ;
        RECT 203.760 87.640 204.295 88.260 ;
        RECT 204.520 88.360 205.680 88.600 ;
        RECT 204.520 87.650 204.780 88.360 ;
        RECT 204.950 87.470 205.280 88.180 ;
        RECT 205.450 87.650 205.680 88.360 ;
        RECT 205.860 88.380 206.630 88.600 ;
        RECT 205.860 87.650 206.130 88.380 ;
        RECT 206.310 87.470 206.650 88.200 ;
        RECT 206.820 87.650 207.080 89.840 ;
        RECT 207.465 89.240 207.965 89.850 ;
        RECT 207.260 88.780 207.610 89.030 ;
        RECT 207.795 88.610 207.965 89.240 ;
        RECT 208.595 89.370 208.925 89.850 ;
        RECT 209.095 89.560 209.320 90.020 ;
        RECT 209.490 89.370 209.820 89.850 ;
        RECT 208.595 89.200 209.820 89.370 ;
        RECT 210.010 89.220 210.260 90.020 ;
        RECT 210.430 89.220 210.770 89.850 ;
        RECT 208.135 88.830 208.465 89.030 ;
        RECT 208.635 88.830 208.965 89.030 ;
        RECT 209.135 88.830 209.555 89.030 ;
        RECT 209.730 88.860 210.425 89.030 ;
        RECT 209.730 88.610 209.900 88.860 ;
        RECT 210.595 88.610 210.770 89.220 ;
        RECT 210.940 89.250 213.530 90.020 ;
        RECT 213.700 89.295 213.990 90.020 ;
        RECT 214.160 89.270 215.370 90.020 ;
        RECT 215.590 89.480 215.815 89.840 ;
        RECT 215.995 89.650 216.325 90.020 ;
        RECT 216.505 89.480 216.760 89.840 ;
        RECT 217.325 89.650 218.070 90.020 ;
        RECT 215.590 89.290 218.075 89.480 ;
        RECT 210.940 88.730 212.150 89.250 ;
        RECT 207.465 88.440 209.900 88.610 ;
        RECT 207.465 87.640 207.795 88.440 ;
        RECT 207.965 87.470 208.295 88.270 ;
        RECT 208.595 87.640 208.925 88.440 ;
        RECT 209.570 87.470 209.820 88.270 ;
        RECT 210.090 87.470 210.260 88.610 ;
        RECT 210.430 87.640 210.770 88.610 ;
        RECT 212.320 88.560 213.530 89.080 ;
        RECT 214.160 88.730 214.680 89.270 ;
        RECT 210.940 87.470 213.530 88.560 ;
        RECT 213.700 87.470 213.990 88.635 ;
        RECT 214.850 88.560 215.370 89.100 ;
        RECT 215.550 88.780 215.820 89.110 ;
        RECT 216.000 88.780 216.435 89.110 ;
        RECT 216.615 88.780 217.190 89.110 ;
        RECT 217.370 88.780 217.650 89.110 ;
        RECT 217.850 88.600 218.075 89.290 ;
        RECT 214.160 87.470 215.370 88.560 ;
        RECT 215.580 88.420 218.075 88.600 ;
        RECT 218.250 88.420 218.585 89.840 ;
        RECT 218.760 89.475 224.105 90.020 ;
        RECT 220.345 88.645 220.685 89.475 ;
        RECT 224.280 89.250 227.790 90.020 ;
        RECT 227.960 89.270 229.170 90.020 ;
        RECT 229.345 89.345 229.620 89.690 ;
        RECT 229.810 89.620 230.190 90.020 ;
        RECT 230.360 89.450 230.530 89.800 ;
        RECT 230.700 89.620 231.030 90.020 ;
        RECT 231.200 89.450 231.455 89.800 ;
        RECT 231.640 89.475 236.985 90.020 ;
        RECT 215.580 87.650 215.870 88.420 ;
        RECT 216.440 88.010 217.630 88.240 ;
        RECT 216.440 87.650 216.700 88.010 ;
        RECT 216.870 87.470 217.200 87.840 ;
        RECT 217.370 87.650 217.630 88.010 ;
        RECT 217.820 87.470 218.150 88.190 ;
        RECT 218.320 87.650 218.585 88.420 ;
        RECT 222.165 87.905 222.515 89.155 ;
        RECT 224.280 88.730 225.930 89.250 ;
        RECT 226.100 88.560 227.790 89.080 ;
        RECT 227.960 88.730 228.480 89.270 ;
        RECT 228.650 88.560 229.170 89.100 ;
        RECT 218.760 87.470 224.105 87.905 ;
        RECT 224.280 87.470 227.790 88.560 ;
        RECT 227.960 87.470 229.170 88.560 ;
        RECT 229.345 88.610 229.515 89.345 ;
        RECT 229.790 89.280 231.455 89.450 ;
        RECT 229.790 89.110 229.960 89.280 ;
        RECT 229.685 88.780 229.960 89.110 ;
        RECT 230.130 88.780 230.955 89.110 ;
        RECT 231.125 88.780 231.470 89.110 ;
        RECT 229.790 88.610 229.960 88.780 ;
        RECT 229.345 87.640 229.620 88.610 ;
        RECT 229.790 88.440 230.450 88.610 ;
        RECT 230.760 88.490 230.955 88.780 ;
        RECT 233.225 88.645 233.565 89.475 ;
        RECT 237.160 89.250 238.830 90.020 ;
        RECT 239.460 89.295 239.750 90.020 ;
        RECT 239.920 89.250 242.510 90.020 ;
        RECT 230.280 88.320 230.450 88.440 ;
        RECT 231.125 88.320 231.450 88.610 ;
        RECT 229.830 87.470 230.110 88.270 ;
        RECT 230.280 88.150 231.450 88.320 ;
        RECT 230.280 87.690 231.470 87.980 ;
        RECT 235.045 87.905 235.395 89.155 ;
        RECT 237.160 88.730 237.910 89.250 ;
        RECT 238.080 88.560 238.830 89.080 ;
        RECT 239.920 88.730 241.130 89.250 ;
        RECT 231.640 87.470 236.985 87.905 ;
        RECT 237.160 87.470 238.830 88.560 ;
        RECT 239.460 87.470 239.750 88.635 ;
        RECT 241.300 88.560 242.510 89.080 ;
        RECT 239.920 87.470 242.510 88.560 ;
        RECT 242.685 88.420 243.020 89.840 ;
        RECT 243.200 89.650 243.945 90.020 ;
        RECT 244.510 89.480 244.765 89.840 ;
        RECT 244.945 89.650 245.275 90.020 ;
        RECT 245.455 89.480 245.680 89.840 ;
        RECT 243.195 89.290 245.680 89.480 ;
        RECT 245.900 89.475 251.245 90.020 ;
        RECT 251.420 89.475 256.765 90.020 ;
        RECT 243.195 88.600 243.420 89.290 ;
        RECT 243.620 88.780 243.900 89.110 ;
        RECT 244.080 88.780 244.655 89.110 ;
        RECT 244.835 88.780 245.270 89.110 ;
        RECT 245.450 88.780 245.720 89.110 ;
        RECT 247.485 88.645 247.825 89.475 ;
        RECT 243.195 88.420 245.690 88.600 ;
        RECT 242.685 87.650 242.950 88.420 ;
        RECT 243.120 87.470 243.450 88.190 ;
        RECT 243.640 88.010 244.830 88.240 ;
        RECT 243.640 87.650 243.900 88.010 ;
        RECT 244.070 87.470 244.400 87.840 ;
        RECT 244.570 87.650 244.830 88.010 ;
        RECT 245.400 87.650 245.690 88.420 ;
        RECT 249.305 87.905 249.655 89.155 ;
        RECT 253.005 88.645 253.345 89.475 ;
        RECT 256.940 89.250 259.530 90.020 ;
        RECT 260.250 89.370 260.420 89.850 ;
        RECT 260.590 89.540 260.920 90.020 ;
        RECT 261.145 89.600 262.680 89.850 ;
        RECT 261.145 89.370 261.315 89.600 ;
        RECT 254.825 87.905 255.175 89.155 ;
        RECT 256.940 88.730 258.150 89.250 ;
        RECT 260.250 89.200 261.315 89.370 ;
        RECT 258.320 88.560 259.530 89.080 ;
        RECT 261.495 89.030 261.775 89.430 ;
        RECT 260.165 88.820 260.515 89.030 ;
        RECT 260.685 88.830 261.130 89.030 ;
        RECT 261.300 88.830 261.775 89.030 ;
        RECT 262.045 89.030 262.330 89.430 ;
        RECT 262.510 89.370 262.680 89.600 ;
        RECT 262.850 89.540 263.180 90.020 ;
        RECT 263.395 89.520 263.650 89.850 ;
        RECT 263.440 89.510 263.650 89.520 ;
        RECT 263.465 89.440 263.650 89.510 ;
        RECT 262.510 89.200 263.310 89.370 ;
        RECT 262.045 88.830 262.375 89.030 ;
        RECT 262.545 88.830 262.910 89.030 ;
        RECT 263.140 88.650 263.310 89.200 ;
        RECT 245.900 87.470 251.245 87.905 ;
        RECT 251.420 87.470 256.765 87.905 ;
        RECT 256.940 87.470 259.530 88.560 ;
        RECT 260.250 88.480 263.310 88.650 ;
        RECT 260.250 87.640 260.420 88.480 ;
        RECT 263.480 88.310 263.650 89.440 ;
        RECT 263.840 89.270 265.050 90.020 ;
        RECT 265.220 89.295 265.510 90.020 ;
        RECT 265.925 89.540 266.225 90.020 ;
        RECT 266.395 89.370 266.655 89.825 ;
        RECT 266.825 89.540 267.085 90.020 ;
        RECT 267.255 89.370 267.515 89.825 ;
        RECT 267.685 89.540 267.945 90.020 ;
        RECT 268.115 89.370 268.375 89.825 ;
        RECT 268.545 89.540 268.805 90.020 ;
        RECT 268.975 89.370 269.235 89.825 ;
        RECT 269.405 89.495 269.665 90.020 ;
        RECT 263.840 88.730 264.360 89.270 ;
        RECT 265.925 89.200 269.235 89.370 ;
        RECT 264.530 88.560 265.050 89.100 ;
        RECT 260.590 87.810 260.920 88.310 ;
        RECT 261.090 88.070 262.725 88.310 ;
        RECT 261.090 87.980 261.320 88.070 ;
        RECT 261.430 87.810 261.760 87.850 ;
        RECT 260.590 87.640 261.760 87.810 ;
        RECT 261.950 87.470 262.305 87.890 ;
        RECT 262.475 87.640 262.725 88.070 ;
        RECT 262.895 87.470 263.225 88.230 ;
        RECT 263.395 87.640 263.650 88.310 ;
        RECT 263.840 87.470 265.050 88.560 ;
        RECT 265.220 87.470 265.510 88.635 ;
        RECT 265.925 88.610 266.895 89.200 ;
        RECT 269.835 89.030 270.085 89.840 ;
        RECT 270.265 89.560 270.510 90.020 ;
        RECT 267.065 88.780 270.085 89.030 ;
        RECT 270.255 88.780 270.570 89.390 ;
        RECT 270.740 89.250 274.250 90.020 ;
        RECT 275.350 89.520 275.680 90.020 ;
        RECT 275.880 89.450 276.050 89.800 ;
        RECT 276.250 89.620 276.580 90.020 ;
        RECT 276.750 89.450 276.920 89.800 ;
        RECT 277.090 89.620 277.470 90.020 ;
        RECT 265.925 88.370 269.235 88.610 ;
        RECT 265.930 87.470 266.225 88.200 ;
        RECT 266.395 87.645 266.655 88.370 ;
        RECT 266.825 87.470 267.085 88.200 ;
        RECT 267.255 87.645 267.515 88.370 ;
        RECT 267.685 87.470 267.945 88.200 ;
        RECT 268.115 87.645 268.375 88.370 ;
        RECT 268.545 87.470 268.805 88.200 ;
        RECT 268.975 87.645 269.235 88.370 ;
        RECT 269.405 87.470 269.665 88.580 ;
        RECT 269.835 87.645 270.085 88.780 ;
        RECT 270.740 88.730 272.390 89.250 ;
        RECT 270.265 87.470 270.560 88.580 ;
        RECT 272.560 88.560 274.250 89.080 ;
        RECT 275.345 88.780 275.695 89.350 ;
        RECT 275.880 89.280 277.490 89.450 ;
        RECT 277.660 89.345 277.930 89.690 ;
        RECT 278.345 89.540 278.645 90.020 ;
        RECT 278.815 89.370 279.075 89.825 ;
        RECT 279.245 89.540 279.505 90.020 ;
        RECT 279.675 89.370 279.935 89.825 ;
        RECT 280.105 89.540 280.365 90.020 ;
        RECT 280.535 89.370 280.795 89.825 ;
        RECT 280.965 89.540 281.225 90.020 ;
        RECT 281.395 89.370 281.655 89.825 ;
        RECT 281.825 89.495 282.085 90.020 ;
        RECT 277.320 89.110 277.490 89.280 ;
        RECT 275.865 88.660 276.575 89.110 ;
        RECT 276.745 88.780 277.150 89.110 ;
        RECT 277.320 88.780 277.590 89.110 ;
        RECT 270.740 87.470 274.250 88.560 ;
        RECT 275.345 88.320 275.665 88.610 ;
        RECT 275.860 88.490 276.575 88.660 ;
        RECT 277.320 88.610 277.490 88.780 ;
        RECT 277.760 88.610 277.930 89.345 ;
        RECT 276.765 88.440 277.490 88.610 ;
        RECT 276.765 88.320 276.935 88.440 ;
        RECT 275.345 88.150 276.935 88.320 ;
        RECT 275.345 87.690 277.000 87.980 ;
        RECT 277.170 87.470 277.450 88.270 ;
        RECT 277.660 87.640 277.930 88.610 ;
        RECT 278.345 89.200 281.655 89.370 ;
        RECT 278.345 88.610 279.315 89.200 ;
        RECT 282.255 89.030 282.505 89.840 ;
        RECT 282.685 89.560 282.930 90.020 ;
        RECT 279.485 88.780 282.505 89.030 ;
        RECT 282.675 88.780 282.990 89.390 ;
        RECT 283.160 89.250 286.670 90.020 ;
        RECT 278.345 88.370 281.655 88.610 ;
        RECT 278.350 87.470 278.645 88.200 ;
        RECT 278.815 87.645 279.075 88.370 ;
        RECT 279.245 87.470 279.505 88.200 ;
        RECT 279.675 87.645 279.935 88.370 ;
        RECT 280.105 87.470 280.365 88.200 ;
        RECT 280.535 87.645 280.795 88.370 ;
        RECT 280.965 87.470 281.225 88.200 ;
        RECT 281.395 87.645 281.655 88.370 ;
        RECT 281.825 87.470 282.085 88.580 ;
        RECT 282.255 87.645 282.505 88.780 ;
        RECT 283.160 88.730 284.810 89.250 ;
        RECT 287.115 89.210 287.360 89.815 ;
        RECT 287.580 89.485 288.090 90.020 ;
        RECT 282.685 87.470 282.980 88.580 ;
        RECT 284.980 88.560 286.670 89.080 ;
        RECT 283.160 87.470 286.670 88.560 ;
        RECT 286.840 89.040 288.070 89.210 ;
        RECT 286.840 88.230 287.180 89.040 ;
        RECT 287.350 88.475 288.100 88.665 ;
        RECT 286.840 87.820 287.355 88.230 ;
        RECT 287.590 87.470 287.760 88.230 ;
        RECT 287.930 87.810 288.100 88.475 ;
        RECT 288.270 88.490 288.460 89.850 ;
        RECT 288.630 89.000 288.905 89.850 ;
        RECT 289.095 89.485 289.625 89.850 ;
        RECT 290.050 89.620 290.380 90.020 ;
        RECT 289.450 89.450 289.625 89.485 ;
        RECT 288.630 88.830 288.910 89.000 ;
        RECT 288.630 88.690 288.905 88.830 ;
        RECT 289.110 88.490 289.280 89.290 ;
        RECT 288.270 88.320 289.280 88.490 ;
        RECT 289.450 89.280 290.380 89.450 ;
        RECT 290.550 89.280 290.805 89.850 ;
        RECT 290.980 89.295 291.270 90.020 ;
        RECT 289.450 88.150 289.620 89.280 ;
        RECT 290.210 89.110 290.380 89.280 ;
        RECT 288.495 87.980 289.620 88.150 ;
        RECT 289.790 88.780 289.985 89.110 ;
        RECT 290.210 88.780 290.465 89.110 ;
        RECT 289.790 87.810 289.960 88.780 ;
        RECT 290.635 88.610 290.805 89.280 ;
        RECT 291.440 89.250 294.950 90.020 ;
        RECT 295.125 89.470 295.380 89.760 ;
        RECT 295.550 89.640 295.880 90.020 ;
        RECT 295.125 89.300 295.875 89.470 ;
        RECT 291.440 88.730 293.090 89.250 ;
        RECT 287.930 87.640 289.960 87.810 ;
        RECT 290.130 87.470 290.300 88.610 ;
        RECT 290.470 87.640 290.805 88.610 ;
        RECT 290.980 87.470 291.270 88.635 ;
        RECT 293.260 88.560 294.950 89.080 ;
        RECT 291.440 87.470 294.950 88.560 ;
        RECT 295.125 88.480 295.475 89.130 ;
        RECT 295.645 88.310 295.875 89.300 ;
        RECT 295.125 88.140 295.875 88.310 ;
        RECT 295.125 87.640 295.380 88.140 ;
        RECT 295.550 87.470 295.880 87.970 ;
        RECT 296.050 87.640 296.220 89.760 ;
        RECT 296.580 89.660 296.910 90.020 ;
        RECT 297.080 89.630 297.575 89.800 ;
        RECT 297.780 89.630 298.635 89.800 ;
        RECT 296.450 88.440 296.910 89.490 ;
        RECT 296.390 87.655 296.715 88.440 ;
        RECT 297.080 88.270 297.250 89.630 ;
        RECT 297.420 88.720 297.770 89.340 ;
        RECT 297.940 89.120 298.295 89.340 ;
        RECT 297.940 88.530 298.110 89.120 ;
        RECT 298.465 88.920 298.635 89.630 ;
        RECT 299.510 89.560 299.840 90.020 ;
        RECT 300.050 89.660 300.400 89.830 ;
        RECT 298.840 89.090 299.630 89.340 ;
        RECT 300.050 89.270 300.310 89.660 ;
        RECT 300.620 89.570 301.570 89.850 ;
        RECT 301.740 89.580 301.930 90.020 ;
        RECT 302.100 89.640 303.170 89.810 ;
        RECT 299.800 88.920 299.970 89.100 ;
        RECT 297.080 88.100 297.475 88.270 ;
        RECT 297.645 88.140 298.110 88.530 ;
        RECT 298.280 88.750 299.970 88.920 ;
        RECT 297.305 87.970 297.475 88.100 ;
        RECT 298.280 87.970 298.450 88.750 ;
        RECT 300.140 88.580 300.310 89.270 ;
        RECT 298.810 88.410 300.310 88.580 ;
        RECT 300.500 88.610 300.710 89.400 ;
        RECT 300.880 88.780 301.230 89.400 ;
        RECT 301.400 88.790 301.570 89.570 ;
        RECT 302.100 89.410 302.270 89.640 ;
        RECT 301.740 89.240 302.270 89.410 ;
        RECT 301.740 88.960 301.960 89.240 ;
        RECT 302.440 89.070 302.680 89.470 ;
        RECT 301.400 88.620 301.805 88.790 ;
        RECT 302.140 88.700 302.680 89.070 ;
        RECT 302.850 89.285 303.170 89.640 ;
        RECT 303.415 89.560 303.720 90.020 ;
        RECT 303.890 89.310 304.140 89.840 ;
        RECT 302.850 89.110 303.175 89.285 ;
        RECT 302.850 88.810 303.765 89.110 ;
        RECT 303.025 88.780 303.765 88.810 ;
        RECT 300.500 88.450 301.175 88.610 ;
        RECT 301.635 88.530 301.805 88.620 ;
        RECT 300.500 88.440 301.465 88.450 ;
        RECT 300.140 88.270 300.310 88.410 ;
        RECT 296.885 87.470 297.135 87.930 ;
        RECT 297.305 87.640 297.555 87.970 ;
        RECT 297.770 87.640 298.450 87.970 ;
        RECT 298.620 88.070 299.695 88.240 ;
        RECT 300.140 88.100 300.700 88.270 ;
        RECT 301.005 88.150 301.465 88.440 ;
        RECT 301.635 88.360 302.855 88.530 ;
        RECT 298.620 87.730 298.790 88.070 ;
        RECT 299.025 87.470 299.355 87.900 ;
        RECT 299.525 87.730 299.695 88.070 ;
        RECT 299.990 87.470 300.360 87.930 ;
        RECT 300.530 87.640 300.700 88.100 ;
        RECT 301.635 87.980 301.805 88.360 ;
        RECT 303.025 88.190 303.195 88.780 ;
        RECT 303.935 88.660 304.140 89.310 ;
        RECT 304.310 89.265 304.560 90.020 ;
        RECT 304.780 89.520 305.080 89.850 ;
        RECT 305.250 89.540 305.525 90.020 ;
        RECT 300.935 87.640 301.805 87.980 ;
        RECT 302.395 88.020 303.195 88.190 ;
        RECT 301.975 87.470 302.225 87.930 ;
        RECT 302.395 87.730 302.565 88.020 ;
        RECT 302.745 87.470 303.075 87.850 ;
        RECT 303.415 87.470 303.720 88.610 ;
        RECT 303.890 87.780 304.140 88.660 ;
        RECT 304.780 88.610 304.950 89.520 ;
        RECT 305.705 89.370 306.000 89.760 ;
        RECT 306.170 89.540 306.425 90.020 ;
        RECT 306.600 89.370 306.860 89.760 ;
        RECT 307.030 89.540 307.310 90.020 ;
        RECT 305.120 88.780 305.470 89.350 ;
        RECT 305.705 89.200 307.355 89.370 ;
        RECT 305.640 88.860 306.780 89.030 ;
        RECT 305.640 88.610 305.810 88.860 ;
        RECT 306.950 88.690 307.355 89.200 ;
        RECT 307.540 89.250 309.210 90.020 ;
        RECT 309.840 89.270 311.050 90.020 ;
        RECT 307.540 88.730 308.290 89.250 ;
        RECT 304.310 87.470 304.560 88.610 ;
        RECT 304.780 88.440 305.810 88.610 ;
        RECT 306.600 88.520 307.355 88.690 ;
        RECT 308.460 88.560 309.210 89.080 ;
        RECT 304.780 87.640 305.090 88.440 ;
        RECT 306.600 88.270 306.860 88.520 ;
        RECT 305.260 87.470 305.570 88.270 ;
        RECT 305.740 88.100 306.860 88.270 ;
        RECT 305.740 87.640 306.000 88.100 ;
        RECT 306.170 87.470 306.425 87.930 ;
        RECT 306.600 87.640 306.860 88.100 ;
        RECT 307.030 87.470 307.315 88.340 ;
        RECT 307.540 87.470 309.210 88.560 ;
        RECT 309.840 88.560 310.360 89.100 ;
        RECT 310.530 88.730 311.050 89.270 ;
        RECT 309.840 87.470 311.050 88.560 ;
        RECT 162.095 87.300 311.135 87.470 ;
        RECT 162.180 86.210 163.390 87.300 ;
        RECT 163.560 86.210 165.230 87.300 ;
        RECT 162.180 85.500 162.700 86.040 ;
        RECT 162.870 85.670 163.390 86.210 ;
        RECT 163.560 85.520 164.310 86.040 ;
        RECT 164.480 85.690 165.230 86.210 ;
        RECT 165.865 86.110 166.120 86.990 ;
        RECT 166.290 86.160 166.595 87.300 ;
        RECT 166.935 86.920 167.265 87.300 ;
        RECT 167.445 86.750 167.615 87.040 ;
        RECT 167.785 86.840 168.035 87.300 ;
        RECT 166.815 86.580 167.615 86.750 ;
        RECT 168.205 86.790 169.075 87.130 ;
        RECT 162.180 84.750 163.390 85.500 ;
        RECT 163.560 84.750 165.230 85.520 ;
        RECT 165.865 85.460 166.075 86.110 ;
        RECT 166.815 85.990 166.985 86.580 ;
        RECT 168.205 86.410 168.375 86.790 ;
        RECT 169.310 86.670 169.480 87.130 ;
        RECT 169.650 86.840 170.020 87.300 ;
        RECT 170.315 86.700 170.485 87.040 ;
        RECT 170.655 86.870 170.985 87.300 ;
        RECT 171.220 86.700 171.390 87.040 ;
        RECT 167.155 86.240 168.375 86.410 ;
        RECT 168.545 86.330 169.005 86.620 ;
        RECT 169.310 86.500 169.870 86.670 ;
        RECT 170.315 86.530 171.390 86.700 ;
        RECT 171.560 86.800 172.240 87.130 ;
        RECT 172.455 86.800 172.705 87.130 ;
        RECT 172.875 86.840 173.125 87.300 ;
        RECT 169.700 86.360 169.870 86.500 ;
        RECT 168.545 86.320 169.510 86.330 ;
        RECT 168.205 86.150 168.375 86.240 ;
        RECT 168.835 86.160 169.510 86.320 ;
        RECT 166.245 85.960 166.985 85.990 ;
        RECT 166.245 85.660 167.160 85.960 ;
        RECT 166.835 85.485 167.160 85.660 ;
        RECT 165.865 84.930 166.120 85.460 ;
        RECT 166.290 84.750 166.595 85.210 ;
        RECT 166.840 85.130 167.160 85.485 ;
        RECT 167.330 85.700 167.870 86.070 ;
        RECT 168.205 85.980 168.610 86.150 ;
        RECT 167.330 85.300 167.570 85.700 ;
        RECT 168.050 85.530 168.270 85.810 ;
        RECT 167.740 85.360 168.270 85.530 ;
        RECT 167.740 85.130 167.910 85.360 ;
        RECT 168.440 85.200 168.610 85.980 ;
        RECT 168.780 85.370 169.130 85.990 ;
        RECT 169.300 85.370 169.510 86.160 ;
        RECT 169.700 86.190 171.200 86.360 ;
        RECT 169.700 85.500 169.870 86.190 ;
        RECT 171.560 86.020 171.730 86.800 ;
        RECT 172.535 86.670 172.705 86.800 ;
        RECT 170.040 85.850 171.730 86.020 ;
        RECT 171.900 86.240 172.365 86.630 ;
        RECT 172.535 86.500 172.930 86.670 ;
        RECT 170.040 85.670 170.210 85.850 ;
        RECT 166.840 84.960 167.910 85.130 ;
        RECT 168.080 84.750 168.270 85.190 ;
        RECT 168.440 84.920 169.390 85.200 ;
        RECT 169.700 85.110 169.960 85.500 ;
        RECT 170.380 85.430 171.170 85.680 ;
        RECT 169.610 84.940 169.960 85.110 ;
        RECT 170.170 84.750 170.500 85.210 ;
        RECT 171.375 85.140 171.545 85.850 ;
        RECT 171.900 85.650 172.070 86.240 ;
        RECT 171.715 85.430 172.070 85.650 ;
        RECT 172.240 85.430 172.590 86.050 ;
        RECT 172.760 85.140 172.930 86.500 ;
        RECT 173.295 86.330 173.620 87.115 ;
        RECT 173.100 85.280 173.560 86.330 ;
        RECT 171.375 84.970 172.230 85.140 ;
        RECT 172.435 84.970 172.930 85.140 ;
        RECT 173.100 84.750 173.430 85.110 ;
        RECT 173.790 85.010 173.960 87.130 ;
        RECT 174.130 86.800 174.460 87.300 ;
        RECT 174.630 86.630 174.885 87.130 ;
        RECT 174.135 86.460 174.885 86.630 ;
        RECT 174.135 85.470 174.365 86.460 ;
        RECT 174.535 85.640 174.885 86.290 ;
        RECT 175.060 86.135 175.350 87.300 ;
        RECT 175.525 86.160 175.860 87.130 ;
        RECT 176.030 86.160 176.200 87.300 ;
        RECT 176.370 86.960 178.400 87.130 ;
        RECT 175.525 85.490 175.695 86.160 ;
        RECT 176.370 85.990 176.540 86.960 ;
        RECT 175.865 85.660 176.120 85.990 ;
        RECT 176.345 85.660 176.540 85.990 ;
        RECT 176.710 86.620 177.835 86.790 ;
        RECT 175.950 85.490 176.120 85.660 ;
        RECT 176.710 85.490 176.880 86.620 ;
        RECT 174.135 85.300 174.885 85.470 ;
        RECT 174.130 84.750 174.460 85.130 ;
        RECT 174.630 85.010 174.885 85.300 ;
        RECT 175.060 84.750 175.350 85.475 ;
        RECT 175.525 84.920 175.780 85.490 ;
        RECT 175.950 85.320 176.880 85.490 ;
        RECT 177.050 86.280 178.060 86.450 ;
        RECT 177.050 85.480 177.220 86.280 ;
        RECT 177.425 85.940 177.700 86.080 ;
        RECT 177.420 85.770 177.700 85.940 ;
        RECT 176.705 85.285 176.880 85.320 ;
        RECT 175.950 84.750 176.280 85.150 ;
        RECT 176.705 84.920 177.235 85.285 ;
        RECT 177.425 84.920 177.700 85.770 ;
        RECT 177.870 84.920 178.060 86.280 ;
        RECT 178.230 86.295 178.400 86.960 ;
        RECT 178.570 86.540 178.740 87.300 ;
        RECT 178.975 86.540 179.490 86.950 ;
        RECT 178.230 86.105 178.980 86.295 ;
        RECT 179.150 85.730 179.490 86.540 ;
        RECT 178.260 85.560 179.490 85.730 ;
        RECT 179.665 86.160 180.000 87.130 ;
        RECT 180.170 86.160 180.340 87.300 ;
        RECT 180.510 86.960 182.540 87.130 ;
        RECT 178.240 84.750 178.750 85.285 ;
        RECT 178.970 84.955 179.215 85.560 ;
        RECT 179.665 85.490 179.835 86.160 ;
        RECT 180.510 85.990 180.680 86.960 ;
        RECT 180.005 85.660 180.260 85.990 ;
        RECT 180.485 85.660 180.680 85.990 ;
        RECT 180.850 86.620 181.975 86.790 ;
        RECT 180.090 85.490 180.260 85.660 ;
        RECT 180.850 85.490 181.020 86.620 ;
        RECT 179.665 84.920 179.920 85.490 ;
        RECT 180.090 85.320 181.020 85.490 ;
        RECT 181.190 86.280 182.200 86.450 ;
        RECT 181.190 85.480 181.360 86.280 ;
        RECT 181.565 85.600 181.840 86.080 ;
        RECT 181.560 85.430 181.840 85.600 ;
        RECT 180.845 85.285 181.020 85.320 ;
        RECT 180.090 84.750 180.420 85.150 ;
        RECT 180.845 84.920 181.375 85.285 ;
        RECT 181.565 84.920 181.840 85.430 ;
        RECT 182.010 84.920 182.200 86.280 ;
        RECT 182.370 86.295 182.540 86.960 ;
        RECT 182.710 86.540 182.880 87.300 ;
        RECT 183.115 86.540 183.630 86.950 ;
        RECT 182.370 86.105 183.120 86.295 ;
        RECT 183.290 85.730 183.630 86.540 ;
        RECT 183.800 86.210 185.470 87.300 ;
        RECT 182.400 85.560 183.630 85.730 ;
        RECT 182.380 84.750 182.890 85.285 ;
        RECT 183.110 84.955 183.355 85.560 ;
        RECT 183.800 85.520 184.550 86.040 ;
        RECT 184.720 85.690 185.470 86.210 ;
        RECT 185.640 86.160 185.930 87.300 ;
        RECT 186.100 86.580 186.550 87.130 ;
        RECT 186.740 86.580 187.070 87.300 ;
        RECT 183.800 84.750 185.470 85.520 ;
        RECT 185.640 84.750 185.930 85.550 ;
        RECT 186.100 85.210 186.350 86.580 ;
        RECT 187.280 86.410 187.580 86.960 ;
        RECT 187.750 86.630 188.030 87.300 ;
        RECT 186.640 86.240 187.580 86.410 ;
        RECT 186.640 85.990 186.810 86.240 ;
        RECT 187.915 85.990 188.230 86.430 ;
        RECT 188.400 86.160 188.690 87.300 ;
        RECT 188.860 86.580 189.310 87.130 ;
        RECT 189.500 86.580 189.830 87.300 ;
        RECT 186.520 85.660 186.810 85.990 ;
        RECT 186.980 85.740 187.310 85.990 ;
        RECT 187.540 85.740 188.230 85.990 ;
        RECT 186.640 85.570 186.810 85.660 ;
        RECT 186.640 85.380 188.030 85.570 ;
        RECT 186.100 84.920 186.650 85.210 ;
        RECT 186.820 84.750 187.070 85.210 ;
        RECT 187.700 85.020 188.030 85.380 ;
        RECT 188.400 84.750 188.690 85.550 ;
        RECT 188.860 85.210 189.110 86.580 ;
        RECT 190.040 86.410 190.340 86.960 ;
        RECT 190.510 86.630 190.790 87.300 ;
        RECT 189.400 86.240 190.340 86.410 ;
        RECT 189.400 85.990 189.570 86.240 ;
        RECT 190.675 85.990 190.990 86.430 ;
        RECT 191.160 86.210 192.830 87.300 ;
        RECT 189.280 85.660 189.570 85.990 ;
        RECT 189.740 85.740 190.070 85.990 ;
        RECT 190.300 85.740 190.990 85.990 ;
        RECT 189.400 85.570 189.570 85.660 ;
        RECT 189.400 85.380 190.790 85.570 ;
        RECT 188.860 84.920 189.410 85.210 ;
        RECT 189.580 84.750 189.830 85.210 ;
        RECT 190.460 85.020 190.790 85.380 ;
        RECT 191.160 85.520 191.910 86.040 ;
        RECT 192.080 85.690 192.830 86.210 ;
        RECT 193.495 86.510 194.030 87.130 ;
        RECT 191.160 84.750 192.830 85.520 ;
        RECT 193.495 85.490 193.810 86.510 ;
        RECT 194.200 86.500 194.530 87.300 ;
        RECT 195.015 86.330 195.405 86.505 ;
        RECT 193.980 86.160 195.405 86.330 ;
        RECT 195.965 86.330 196.295 87.130 ;
        RECT 196.465 86.500 196.795 87.300 ;
        RECT 197.095 86.330 197.425 87.130 ;
        RECT 198.070 86.500 198.320 87.300 ;
        RECT 195.965 86.160 198.400 86.330 ;
        RECT 198.590 86.160 198.760 87.300 ;
        RECT 198.930 86.160 199.270 87.130 ;
        RECT 199.440 86.210 200.650 87.300 ;
        RECT 193.980 85.660 194.150 86.160 ;
        RECT 193.495 84.920 194.110 85.490 ;
        RECT 194.400 85.430 194.665 85.990 ;
        RECT 194.835 85.260 195.005 86.160 ;
        RECT 195.175 85.430 195.530 85.990 ;
        RECT 195.760 85.740 196.110 85.990 ;
        RECT 196.295 85.530 196.465 86.160 ;
        RECT 196.635 85.740 196.965 85.940 ;
        RECT 197.135 85.740 197.465 85.940 ;
        RECT 197.635 85.740 198.055 85.940 ;
        RECT 198.230 85.910 198.400 86.160 ;
        RECT 198.230 85.740 198.925 85.910 ;
        RECT 194.280 84.750 194.495 85.260 ;
        RECT 194.725 84.930 195.005 85.260 ;
        RECT 195.185 84.750 195.425 85.260 ;
        RECT 195.965 84.920 196.465 85.530 ;
        RECT 197.095 85.400 198.320 85.570 ;
        RECT 199.095 85.550 199.270 86.160 ;
        RECT 197.095 84.920 197.425 85.400 ;
        RECT 197.595 84.750 197.820 85.210 ;
        RECT 197.990 84.920 198.320 85.400 ;
        RECT 198.510 84.750 198.760 85.550 ;
        RECT 198.930 84.920 199.270 85.550 ;
        RECT 199.440 85.500 199.960 86.040 ;
        RECT 200.130 85.670 200.650 86.210 ;
        RECT 200.820 86.135 201.110 87.300 ;
        RECT 202.385 86.330 202.775 86.505 ;
        RECT 203.260 86.500 203.590 87.300 ;
        RECT 203.760 86.510 204.295 87.130 ;
        RECT 202.385 86.160 203.810 86.330 ;
        RECT 199.440 84.750 200.650 85.500 ;
        RECT 200.820 84.750 201.110 85.475 ;
        RECT 202.260 85.430 202.615 85.990 ;
        RECT 202.785 85.260 202.955 86.160 ;
        RECT 203.125 85.430 203.390 85.990 ;
        RECT 203.640 85.660 203.810 86.160 ;
        RECT 203.980 85.490 204.295 86.510 ;
        RECT 205.625 86.330 205.955 87.130 ;
        RECT 206.125 86.500 206.455 87.300 ;
        RECT 206.755 86.330 207.085 87.130 ;
        RECT 207.730 86.500 207.980 87.300 ;
        RECT 205.625 86.160 208.060 86.330 ;
        RECT 208.250 86.160 208.420 87.300 ;
        RECT 208.590 86.160 208.930 87.130 ;
        RECT 209.100 86.210 210.310 87.300 ;
        RECT 205.420 85.740 205.770 85.990 ;
        RECT 205.955 85.530 206.125 86.160 ;
        RECT 206.295 85.740 206.625 85.940 ;
        RECT 206.795 85.740 207.125 85.940 ;
        RECT 207.295 85.740 207.715 85.940 ;
        RECT 207.890 85.910 208.060 86.160 ;
        RECT 207.890 85.740 208.585 85.910 ;
        RECT 202.365 84.750 202.605 85.260 ;
        RECT 202.785 84.930 203.065 85.260 ;
        RECT 203.295 84.750 203.510 85.260 ;
        RECT 203.680 84.920 204.295 85.490 ;
        RECT 205.625 84.920 206.125 85.530 ;
        RECT 206.755 85.400 207.980 85.570 ;
        RECT 208.755 85.550 208.930 86.160 ;
        RECT 206.755 84.920 207.085 85.400 ;
        RECT 207.255 84.750 207.480 85.210 ;
        RECT 207.650 84.920 207.980 85.400 ;
        RECT 208.170 84.750 208.420 85.550 ;
        RECT 208.590 84.920 208.930 85.550 ;
        RECT 209.100 85.500 209.620 86.040 ;
        RECT 209.790 85.670 210.310 86.210 ;
        RECT 210.665 86.330 211.055 86.505 ;
        RECT 211.540 86.500 211.870 87.300 ;
        RECT 212.040 86.510 212.575 87.130 ;
        RECT 212.780 86.865 218.125 87.300 ;
        RECT 218.300 86.865 223.645 87.300 ;
        RECT 210.665 86.160 212.090 86.330 ;
        RECT 209.100 84.750 210.310 85.500 ;
        RECT 210.540 85.430 210.895 85.990 ;
        RECT 211.065 85.260 211.235 86.160 ;
        RECT 211.405 85.430 211.670 85.990 ;
        RECT 211.920 85.660 212.090 86.160 ;
        RECT 212.260 85.490 212.575 86.510 ;
        RECT 210.645 84.750 210.885 85.260 ;
        RECT 211.065 84.930 211.345 85.260 ;
        RECT 211.575 84.750 211.790 85.260 ;
        RECT 211.960 84.920 212.575 85.490 ;
        RECT 214.365 85.295 214.705 86.125 ;
        RECT 216.185 85.615 216.535 86.865 ;
        RECT 219.885 85.295 220.225 86.125 ;
        RECT 221.705 85.615 222.055 86.865 ;
        RECT 223.820 86.210 226.410 87.300 ;
        RECT 223.820 85.520 225.030 86.040 ;
        RECT 225.200 85.690 226.410 86.210 ;
        RECT 226.580 86.135 226.870 87.300 ;
        RECT 227.040 86.865 232.385 87.300 ;
        RECT 232.560 86.865 237.905 87.300 ;
        RECT 212.780 84.750 218.125 85.295 ;
        RECT 218.300 84.750 223.645 85.295 ;
        RECT 223.820 84.750 226.410 85.520 ;
        RECT 226.580 84.750 226.870 85.475 ;
        RECT 228.625 85.295 228.965 86.125 ;
        RECT 230.445 85.615 230.795 86.865 ;
        RECT 234.145 85.295 234.485 86.125 ;
        RECT 235.965 85.615 236.315 86.865 ;
        RECT 238.080 86.210 241.590 87.300 ;
        RECT 238.080 85.520 239.730 86.040 ;
        RECT 239.900 85.690 241.590 86.210 ;
        RECT 242.225 86.150 242.485 87.300 ;
        RECT 242.660 86.225 242.915 87.130 ;
        RECT 243.085 86.540 243.415 87.300 ;
        RECT 243.630 86.370 243.800 87.130 ;
        RECT 244.100 86.960 245.240 87.130 ;
        RECT 244.100 86.500 244.400 86.960 ;
        RECT 227.040 84.750 232.385 85.295 ;
        RECT 232.560 84.750 237.905 85.295 ;
        RECT 238.080 84.750 241.590 85.520 ;
        RECT 242.225 84.750 242.485 85.590 ;
        RECT 242.660 85.495 242.830 86.225 ;
        RECT 243.085 86.200 243.800 86.370 ;
        RECT 244.570 86.330 244.900 86.790 ;
        RECT 243.085 85.990 243.255 86.200 ;
        RECT 244.140 86.110 244.900 86.330 ;
        RECT 245.070 86.330 245.240 86.960 ;
        RECT 245.410 86.500 245.740 87.300 ;
        RECT 245.910 86.330 246.185 87.130 ;
        RECT 247.365 86.680 247.540 87.130 ;
        RECT 247.710 86.860 248.040 87.300 ;
        RECT 248.345 86.710 248.515 87.130 ;
        RECT 248.750 86.890 249.420 87.300 ;
        RECT 249.635 86.710 249.805 87.130 ;
        RECT 250.005 86.890 250.335 87.300 ;
        RECT 247.365 86.510 247.995 86.680 ;
        RECT 245.070 86.120 246.185 86.330 ;
        RECT 243.000 85.660 243.255 85.990 ;
        RECT 242.660 84.920 242.915 85.495 ;
        RECT 243.085 85.470 243.255 85.660 ;
        RECT 243.535 85.650 243.890 86.020 ;
        RECT 244.140 85.570 244.355 86.110 ;
        RECT 244.525 85.740 245.295 85.940 ;
        RECT 245.465 85.740 246.185 85.940 ;
        RECT 247.280 85.660 247.645 86.340 ;
        RECT 247.825 85.990 247.995 86.510 ;
        RECT 248.345 86.540 250.360 86.710 ;
        RECT 247.825 85.660 248.175 85.990 ;
        RECT 243.085 85.300 243.800 85.470 ;
        RECT 244.140 85.400 245.740 85.570 ;
        RECT 243.085 84.750 243.415 85.130 ;
        RECT 243.630 84.920 243.800 85.300 ;
        RECT 244.570 85.390 245.740 85.400 ;
        RECT 244.110 84.750 244.400 85.220 ;
        RECT 244.570 84.920 244.900 85.390 ;
        RECT 245.070 84.750 245.240 85.220 ;
        RECT 245.410 84.920 245.740 85.390 ;
        RECT 245.910 84.750 246.185 85.570 ;
        RECT 247.825 85.490 247.995 85.660 ;
        RECT 247.365 85.320 247.995 85.490 ;
        RECT 247.365 84.920 247.540 85.320 ;
        RECT 248.345 85.250 248.515 86.540 ;
        RECT 247.710 84.750 248.040 85.130 ;
        RECT 248.285 84.920 248.515 85.250 ;
        RECT 248.715 85.085 248.995 86.360 ;
        RECT 249.220 86.280 249.490 86.360 ;
        RECT 249.180 86.110 249.490 86.280 ;
        RECT 249.220 85.085 249.490 86.110 ;
        RECT 249.680 85.330 250.020 86.360 ;
        RECT 250.190 85.990 250.360 86.540 ;
        RECT 250.530 86.160 250.790 87.130 ;
        RECT 250.960 86.210 252.170 87.300 ;
        RECT 250.190 85.660 250.450 85.990 ;
        RECT 250.620 85.470 250.790 86.160 ;
        RECT 249.950 84.750 250.280 85.130 ;
        RECT 250.450 85.005 250.790 85.470 ;
        RECT 250.960 85.500 251.480 86.040 ;
        RECT 251.650 85.670 252.170 86.210 ;
        RECT 252.340 86.135 252.630 87.300 ;
        RECT 252.800 86.865 258.145 87.300 ;
        RECT 258.320 86.865 263.665 87.300 ;
        RECT 250.450 84.960 250.785 85.005 ;
        RECT 250.960 84.750 252.170 85.500 ;
        RECT 252.340 84.750 252.630 85.475 ;
        RECT 254.385 85.295 254.725 86.125 ;
        RECT 256.205 85.615 256.555 86.865 ;
        RECT 259.905 85.295 260.245 86.125 ;
        RECT 261.725 85.615 262.075 86.865 ;
        RECT 264.400 86.840 264.570 87.300 ;
        RECT 264.740 86.350 265.070 87.130 ;
        RECT 265.240 86.500 265.410 87.300 ;
        RECT 264.300 86.330 265.070 86.350 ;
        RECT 265.580 86.330 265.910 87.130 ;
        RECT 266.080 86.500 266.250 87.300 ;
        RECT 266.420 86.330 266.750 87.130 ;
        RECT 264.300 86.160 266.750 86.330 ;
        RECT 267.010 86.160 267.305 87.300 ;
        RECT 267.520 86.865 272.865 87.300 ;
        RECT 264.300 85.570 264.650 86.160 ;
        RECT 264.820 85.740 267.330 85.990 ;
        RECT 264.300 85.390 266.670 85.570 ;
        RECT 252.800 84.750 258.145 85.295 ;
        RECT 258.320 84.750 263.665 85.295 ;
        RECT 264.400 84.750 264.650 85.215 ;
        RECT 264.820 84.920 264.990 85.390 ;
        RECT 265.240 84.750 265.410 85.210 ;
        RECT 265.660 84.920 265.830 85.390 ;
        RECT 266.080 84.750 266.250 85.210 ;
        RECT 266.500 84.920 266.670 85.390 ;
        RECT 269.105 85.295 269.445 86.125 ;
        RECT 270.925 85.615 271.275 86.865 ;
        RECT 273.040 86.210 276.550 87.300 ;
        RECT 276.720 86.210 277.930 87.300 ;
        RECT 273.040 85.520 274.690 86.040 ;
        RECT 274.860 85.690 276.550 86.210 ;
        RECT 267.040 84.750 267.305 85.210 ;
        RECT 267.520 84.750 272.865 85.295 ;
        RECT 273.040 84.750 276.550 85.520 ;
        RECT 276.720 85.500 277.240 86.040 ;
        RECT 277.410 85.670 277.930 86.210 ;
        RECT 278.100 86.135 278.390 87.300 ;
        RECT 278.570 86.160 278.900 87.300 ;
        RECT 276.720 84.750 277.930 85.500 ;
        RECT 278.100 84.750 278.390 85.475 ;
        RECT 278.560 85.410 278.900 85.990 ;
        RECT 279.070 85.960 279.430 87.130 ;
        RECT 279.630 86.130 279.960 87.300 ;
        RECT 280.160 85.960 280.490 87.130 ;
        RECT 280.690 86.130 281.020 87.300 ;
        RECT 279.070 85.680 280.490 85.960 ;
        RECT 279.070 85.345 279.430 85.680 ;
        RECT 278.570 84.750 278.900 85.240 ;
        RECT 279.070 84.920 279.690 85.345 ;
        RECT 280.150 84.750 280.480 85.440 ;
        RECT 281.790 84.930 282.050 87.120 ;
        RECT 282.220 86.570 282.560 87.300 ;
        RECT 282.740 86.390 283.010 87.120 ;
        RECT 282.240 86.170 283.010 86.390 ;
        RECT 283.190 86.410 283.420 87.120 ;
        RECT 283.590 86.590 283.920 87.300 ;
        RECT 284.090 86.410 284.350 87.120 ;
        RECT 283.190 86.170 284.350 86.410 ;
        RECT 284.540 86.210 288.050 87.300 ;
        RECT 288.685 86.630 288.940 87.130 ;
        RECT 289.110 86.800 289.440 87.300 ;
        RECT 288.685 86.460 289.435 86.630 ;
        RECT 282.240 85.500 282.530 86.170 ;
        RECT 282.710 85.680 283.175 85.990 ;
        RECT 283.355 85.680 283.880 85.990 ;
        RECT 282.240 85.300 283.470 85.500 ;
        RECT 282.310 84.750 282.980 85.120 ;
        RECT 283.160 84.930 283.470 85.300 ;
        RECT 283.650 85.040 283.880 85.680 ;
        RECT 284.060 85.660 284.360 85.990 ;
        RECT 284.540 85.520 286.190 86.040 ;
        RECT 286.360 85.690 288.050 86.210 ;
        RECT 288.685 85.640 289.035 86.290 ;
        RECT 284.060 84.750 284.350 85.480 ;
        RECT 284.540 84.750 288.050 85.520 ;
        RECT 289.205 85.470 289.435 86.460 ;
        RECT 288.685 85.300 289.435 85.470 ;
        RECT 288.685 85.010 288.940 85.300 ;
        RECT 289.110 84.750 289.440 85.130 ;
        RECT 289.610 85.010 289.780 87.130 ;
        RECT 289.950 86.330 290.275 87.115 ;
        RECT 290.445 86.840 290.695 87.300 ;
        RECT 290.865 86.800 291.115 87.130 ;
        RECT 291.330 86.800 292.010 87.130 ;
        RECT 290.865 86.670 291.035 86.800 ;
        RECT 290.640 86.500 291.035 86.670 ;
        RECT 290.010 85.280 290.470 86.330 ;
        RECT 290.640 85.140 290.810 86.500 ;
        RECT 291.205 86.240 291.670 86.630 ;
        RECT 290.980 85.430 291.330 86.050 ;
        RECT 291.500 85.650 291.670 86.240 ;
        RECT 291.840 86.020 292.010 86.800 ;
        RECT 292.180 86.700 292.350 87.040 ;
        RECT 292.585 86.870 292.915 87.300 ;
        RECT 293.085 86.700 293.255 87.040 ;
        RECT 293.550 86.840 293.920 87.300 ;
        RECT 292.180 86.530 293.255 86.700 ;
        RECT 294.090 86.670 294.260 87.130 ;
        RECT 294.495 86.790 295.365 87.130 ;
        RECT 295.535 86.840 295.785 87.300 ;
        RECT 293.700 86.500 294.260 86.670 ;
        RECT 293.700 86.360 293.870 86.500 ;
        RECT 292.370 86.190 293.870 86.360 ;
        RECT 294.565 86.330 295.025 86.620 ;
        RECT 291.840 85.850 293.530 86.020 ;
        RECT 291.500 85.430 291.855 85.650 ;
        RECT 292.025 85.140 292.195 85.850 ;
        RECT 292.400 85.430 293.190 85.680 ;
        RECT 293.360 85.670 293.530 85.850 ;
        RECT 293.700 85.500 293.870 86.190 ;
        RECT 290.140 84.750 290.470 85.110 ;
        RECT 290.640 84.970 291.135 85.140 ;
        RECT 291.340 84.970 292.195 85.140 ;
        RECT 293.070 84.750 293.400 85.210 ;
        RECT 293.610 85.110 293.870 85.500 ;
        RECT 294.060 86.320 295.025 86.330 ;
        RECT 295.195 86.410 295.365 86.790 ;
        RECT 295.955 86.750 296.125 87.040 ;
        RECT 296.305 86.920 296.635 87.300 ;
        RECT 295.955 86.580 296.755 86.750 ;
        RECT 294.060 86.160 294.735 86.320 ;
        RECT 295.195 86.240 296.415 86.410 ;
        RECT 294.060 85.370 294.270 86.160 ;
        RECT 295.195 86.150 295.365 86.240 ;
        RECT 294.440 85.370 294.790 85.990 ;
        RECT 294.960 85.980 295.365 86.150 ;
        RECT 294.960 85.200 295.130 85.980 ;
        RECT 295.300 85.530 295.520 85.810 ;
        RECT 295.700 85.700 296.240 86.070 ;
        RECT 296.585 85.990 296.755 86.580 ;
        RECT 296.975 86.160 297.280 87.300 ;
        RECT 297.450 86.110 297.705 86.990 ;
        RECT 296.585 85.960 297.325 85.990 ;
        RECT 295.300 85.360 295.830 85.530 ;
        RECT 293.610 84.940 293.960 85.110 ;
        RECT 294.180 84.920 295.130 85.200 ;
        RECT 295.300 84.750 295.490 85.190 ;
        RECT 295.660 85.130 295.830 85.360 ;
        RECT 296.000 85.300 296.240 85.700 ;
        RECT 296.410 85.660 297.325 85.960 ;
        RECT 296.410 85.485 296.735 85.660 ;
        RECT 296.410 85.130 296.730 85.485 ;
        RECT 297.495 85.460 297.705 86.110 ;
        RECT 295.660 84.960 296.730 85.130 ;
        RECT 296.975 84.750 297.280 85.210 ;
        RECT 297.450 84.930 297.705 85.460 ;
        RECT 297.885 86.160 298.220 87.130 ;
        RECT 298.390 86.160 298.560 87.300 ;
        RECT 298.730 86.960 300.760 87.130 ;
        RECT 297.885 85.490 298.055 86.160 ;
        RECT 298.730 85.990 298.900 86.960 ;
        RECT 298.225 85.660 298.480 85.990 ;
        RECT 298.705 85.660 298.900 85.990 ;
        RECT 299.070 86.620 300.195 86.790 ;
        RECT 298.310 85.490 298.480 85.660 ;
        RECT 299.070 85.490 299.240 86.620 ;
        RECT 297.885 84.920 298.140 85.490 ;
        RECT 298.310 85.320 299.240 85.490 ;
        RECT 299.410 86.280 300.420 86.450 ;
        RECT 299.410 85.480 299.580 86.280 ;
        RECT 299.785 85.600 300.060 86.080 ;
        RECT 299.780 85.430 300.060 85.600 ;
        RECT 299.065 85.285 299.240 85.320 ;
        RECT 298.310 84.750 298.640 85.150 ;
        RECT 299.065 84.920 299.595 85.285 ;
        RECT 299.785 84.920 300.060 85.430 ;
        RECT 300.230 84.920 300.420 86.280 ;
        RECT 300.590 86.295 300.760 86.960 ;
        RECT 300.930 86.540 301.100 87.300 ;
        RECT 301.335 86.540 301.850 86.950 ;
        RECT 300.590 86.105 301.340 86.295 ;
        RECT 301.510 85.730 301.850 86.540 ;
        RECT 302.020 86.210 303.690 87.300 ;
        RECT 300.620 85.560 301.850 85.730 ;
        RECT 300.600 84.750 301.110 85.285 ;
        RECT 301.330 84.955 301.575 85.560 ;
        RECT 302.020 85.520 302.770 86.040 ;
        RECT 302.940 85.690 303.690 86.210 ;
        RECT 303.860 86.135 304.150 87.300 ;
        RECT 304.325 86.160 304.660 87.130 ;
        RECT 304.830 86.160 305.000 87.300 ;
        RECT 305.170 86.960 307.200 87.130 ;
        RECT 302.020 84.750 303.690 85.520 ;
        RECT 304.325 85.490 304.495 86.160 ;
        RECT 305.170 85.990 305.340 86.960 ;
        RECT 304.665 85.660 304.920 85.990 ;
        RECT 305.145 85.660 305.340 85.990 ;
        RECT 305.510 86.620 306.635 86.790 ;
        RECT 304.750 85.490 304.920 85.660 ;
        RECT 305.510 85.490 305.680 86.620 ;
        RECT 303.860 84.750 304.150 85.475 ;
        RECT 304.325 84.920 304.580 85.490 ;
        RECT 304.750 85.320 305.680 85.490 ;
        RECT 305.850 86.280 306.860 86.450 ;
        RECT 305.850 85.480 306.020 86.280 ;
        RECT 306.225 85.940 306.500 86.080 ;
        RECT 306.220 85.770 306.500 85.940 ;
        RECT 305.505 85.285 305.680 85.320 ;
        RECT 304.750 84.750 305.080 85.150 ;
        RECT 305.505 84.920 306.035 85.285 ;
        RECT 306.225 84.920 306.500 85.770 ;
        RECT 306.670 84.920 306.860 86.280 ;
        RECT 307.030 86.295 307.200 86.960 ;
        RECT 307.370 86.540 307.540 87.300 ;
        RECT 307.775 86.540 308.290 86.950 ;
        RECT 307.030 86.105 307.780 86.295 ;
        RECT 307.950 85.730 308.290 86.540 ;
        RECT 307.060 85.560 308.290 85.730 ;
        RECT 308.460 86.225 308.730 87.130 ;
        RECT 308.900 86.540 309.230 87.300 ;
        RECT 309.410 86.370 309.580 87.130 ;
        RECT 307.040 84.750 307.550 85.285 ;
        RECT 307.770 84.955 308.015 85.560 ;
        RECT 308.460 85.425 308.630 86.225 ;
        RECT 308.915 86.200 309.580 86.370 ;
        RECT 309.840 86.210 311.050 87.300 ;
        RECT 308.915 86.055 309.085 86.200 ;
        RECT 308.800 85.725 309.085 86.055 ;
        RECT 308.915 85.470 309.085 85.725 ;
        RECT 309.320 85.650 309.650 86.020 ;
        RECT 309.840 85.670 310.360 86.210 ;
        RECT 310.530 85.500 311.050 86.040 ;
        RECT 308.460 84.920 308.720 85.425 ;
        RECT 308.915 85.300 309.580 85.470 ;
        RECT 308.900 84.750 309.230 85.130 ;
        RECT 309.410 84.920 309.580 85.300 ;
        RECT 309.840 84.750 311.050 85.500 ;
        RECT 162.095 84.580 311.135 84.750 ;
        RECT 162.180 83.830 163.390 84.580 ;
        RECT 163.560 84.035 168.905 84.580 ;
        RECT 162.180 83.290 162.700 83.830 ;
        RECT 162.870 83.120 163.390 83.660 ;
        RECT 165.145 83.205 165.485 84.035 ;
        RECT 169.080 83.810 170.750 84.580 ;
        RECT 170.925 83.870 171.180 84.400 ;
        RECT 171.350 84.120 171.655 84.580 ;
        RECT 171.900 84.200 172.970 84.370 ;
        RECT 162.180 82.030 163.390 83.120 ;
        RECT 166.965 82.465 167.315 83.715 ;
        RECT 169.080 83.290 169.830 83.810 ;
        RECT 170.000 83.120 170.750 83.640 ;
        RECT 163.560 82.030 168.905 82.465 ;
        RECT 169.080 82.030 170.750 83.120 ;
        RECT 170.925 83.220 171.135 83.870 ;
        RECT 171.900 83.845 172.220 84.200 ;
        RECT 171.895 83.670 172.220 83.845 ;
        RECT 171.305 83.370 172.220 83.670 ;
        RECT 172.390 83.630 172.630 84.030 ;
        RECT 172.800 83.970 172.970 84.200 ;
        RECT 173.140 84.140 173.330 84.580 ;
        RECT 173.500 84.130 174.450 84.410 ;
        RECT 174.670 84.220 175.020 84.390 ;
        RECT 172.800 83.800 173.330 83.970 ;
        RECT 171.305 83.340 172.045 83.370 ;
        RECT 170.925 82.340 171.180 83.220 ;
        RECT 171.350 82.030 171.655 83.170 ;
        RECT 171.875 82.750 172.045 83.340 ;
        RECT 172.390 83.260 172.930 83.630 ;
        RECT 173.110 83.520 173.330 83.800 ;
        RECT 173.500 83.350 173.670 84.130 ;
        RECT 173.265 83.180 173.670 83.350 ;
        RECT 173.840 83.340 174.190 83.960 ;
        RECT 173.265 83.090 173.435 83.180 ;
        RECT 174.360 83.170 174.570 83.960 ;
        RECT 172.215 82.920 173.435 83.090 ;
        RECT 173.895 83.010 174.570 83.170 ;
        RECT 171.875 82.580 172.675 82.750 ;
        RECT 171.995 82.030 172.325 82.410 ;
        RECT 172.505 82.290 172.675 82.580 ;
        RECT 173.265 82.540 173.435 82.920 ;
        RECT 173.605 83.000 174.570 83.010 ;
        RECT 174.760 83.830 175.020 84.220 ;
        RECT 175.230 84.120 175.560 84.580 ;
        RECT 176.435 84.190 177.290 84.360 ;
        RECT 177.495 84.190 177.990 84.360 ;
        RECT 178.160 84.220 178.490 84.580 ;
        RECT 174.760 83.140 174.930 83.830 ;
        RECT 175.100 83.480 175.270 83.660 ;
        RECT 175.440 83.650 176.230 83.900 ;
        RECT 176.435 83.480 176.605 84.190 ;
        RECT 176.775 83.680 177.130 83.900 ;
        RECT 175.100 83.310 176.790 83.480 ;
        RECT 173.605 82.710 174.065 83.000 ;
        RECT 174.760 82.970 176.260 83.140 ;
        RECT 174.760 82.830 174.930 82.970 ;
        RECT 174.370 82.660 174.930 82.830 ;
        RECT 172.845 82.030 173.095 82.490 ;
        RECT 173.265 82.200 174.135 82.540 ;
        RECT 174.370 82.200 174.540 82.660 ;
        RECT 175.375 82.630 176.450 82.800 ;
        RECT 174.710 82.030 175.080 82.490 ;
        RECT 175.375 82.290 175.545 82.630 ;
        RECT 175.715 82.030 176.045 82.460 ;
        RECT 176.280 82.290 176.450 82.630 ;
        RECT 176.620 82.530 176.790 83.310 ;
        RECT 176.960 83.090 177.130 83.680 ;
        RECT 177.300 83.280 177.650 83.900 ;
        RECT 176.960 82.700 177.425 83.090 ;
        RECT 177.820 82.830 177.990 84.190 ;
        RECT 178.160 83.000 178.620 84.050 ;
        RECT 177.595 82.660 177.990 82.830 ;
        RECT 177.595 82.530 177.765 82.660 ;
        RECT 176.620 82.200 177.300 82.530 ;
        RECT 177.515 82.200 177.765 82.530 ;
        RECT 177.935 82.030 178.185 82.490 ;
        RECT 178.355 82.215 178.680 83.000 ;
        RECT 178.850 82.200 179.020 84.320 ;
        RECT 179.190 84.200 179.520 84.580 ;
        RECT 179.690 84.030 179.945 84.320 ;
        RECT 179.195 83.860 179.945 84.030 ;
        RECT 179.195 82.870 179.425 83.860 ;
        RECT 180.120 83.810 182.710 84.580 ;
        RECT 179.595 83.040 179.945 83.690 ;
        RECT 180.120 83.290 181.330 83.810 ;
        RECT 181.500 83.120 182.710 83.640 ;
        RECT 179.195 82.700 179.945 82.870 ;
        RECT 179.190 82.030 179.520 82.530 ;
        RECT 179.690 82.200 179.945 82.700 ;
        RECT 180.120 82.030 182.710 83.120 ;
        RECT 183.340 83.635 183.680 84.410 ;
        RECT 183.850 84.120 184.020 84.580 ;
        RECT 184.260 84.145 184.620 84.410 ;
        RECT 184.260 84.140 184.615 84.145 ;
        RECT 184.260 84.130 184.610 84.140 ;
        RECT 184.260 84.125 184.605 84.130 ;
        RECT 184.260 84.115 184.600 84.125 ;
        RECT 185.250 84.120 185.420 84.580 ;
        RECT 184.260 84.110 184.595 84.115 ;
        RECT 184.260 84.100 184.585 84.110 ;
        RECT 184.260 84.090 184.575 84.100 ;
        RECT 184.260 83.950 184.560 84.090 ;
        RECT 183.850 83.760 184.560 83.950 ;
        RECT 184.750 83.950 185.080 84.030 ;
        RECT 185.590 83.950 185.930 84.410 ;
        RECT 184.750 83.760 185.930 83.950 ;
        RECT 186.100 83.810 187.770 84.580 ;
        RECT 187.940 83.855 188.230 84.580 ;
        RECT 183.340 82.200 183.620 83.635 ;
        RECT 183.850 83.190 184.135 83.760 ;
        RECT 184.320 83.360 184.790 83.590 ;
        RECT 184.960 83.570 185.290 83.590 ;
        RECT 184.960 83.390 185.410 83.570 ;
        RECT 185.600 83.390 185.930 83.590 ;
        RECT 183.850 82.975 185.000 83.190 ;
        RECT 183.790 82.030 184.500 82.805 ;
        RECT 184.670 82.200 185.000 82.975 ;
        RECT 185.195 82.275 185.410 83.390 ;
        RECT 185.700 83.050 185.930 83.390 ;
        RECT 186.100 83.290 186.850 83.810 ;
        RECT 188.400 83.780 188.690 84.580 ;
        RECT 188.860 84.120 189.410 84.410 ;
        RECT 189.580 84.120 189.830 84.580 ;
        RECT 187.020 83.120 187.770 83.640 ;
        RECT 185.590 82.030 185.920 82.750 ;
        RECT 186.100 82.030 187.770 83.120 ;
        RECT 187.940 82.030 188.230 83.195 ;
        RECT 188.400 82.030 188.690 83.170 ;
        RECT 188.860 82.750 189.110 84.120 ;
        RECT 190.460 83.950 190.790 84.310 ;
        RECT 191.160 84.035 196.505 84.580 ;
        RECT 196.680 84.035 202.025 84.580 ;
        RECT 189.400 83.760 190.790 83.950 ;
        RECT 189.400 83.670 189.570 83.760 ;
        RECT 189.280 83.340 189.570 83.670 ;
        RECT 189.740 83.340 190.070 83.590 ;
        RECT 190.300 83.340 190.990 83.590 ;
        RECT 189.400 83.090 189.570 83.340 ;
        RECT 189.400 82.920 190.340 83.090 ;
        RECT 188.860 82.200 189.310 82.750 ;
        RECT 189.500 82.030 189.830 82.750 ;
        RECT 190.040 82.370 190.340 82.920 ;
        RECT 190.675 82.900 190.990 83.340 ;
        RECT 192.745 83.205 193.085 84.035 ;
        RECT 190.510 82.030 190.790 82.700 ;
        RECT 194.565 82.465 194.915 83.715 ;
        RECT 198.265 83.205 198.605 84.035 ;
        RECT 202.200 83.810 205.710 84.580 ;
        RECT 206.810 84.090 207.140 84.580 ;
        RECT 207.310 83.985 207.930 84.410 ;
        RECT 200.085 82.465 200.435 83.715 ;
        RECT 202.200 83.290 203.850 83.810 ;
        RECT 204.020 83.120 205.710 83.640 ;
        RECT 206.800 83.340 207.140 83.920 ;
        RECT 207.310 83.650 207.670 83.985 ;
        RECT 208.390 83.890 208.720 84.580 ;
        RECT 210.225 83.800 210.725 84.410 ;
        RECT 207.310 83.370 208.730 83.650 ;
        RECT 191.160 82.030 196.505 82.465 ;
        RECT 196.680 82.030 202.025 82.465 ;
        RECT 202.200 82.030 205.710 83.120 ;
        RECT 206.810 82.030 207.140 83.170 ;
        RECT 207.310 82.200 207.670 83.370 ;
        RECT 207.870 82.030 208.200 83.200 ;
        RECT 208.400 82.200 208.730 83.370 ;
        RECT 210.020 83.340 210.370 83.590 ;
        RECT 208.930 82.030 209.260 83.200 ;
        RECT 210.555 83.170 210.725 83.800 ;
        RECT 211.355 83.930 211.685 84.410 ;
        RECT 211.855 84.120 212.080 84.580 ;
        RECT 212.250 83.930 212.580 84.410 ;
        RECT 211.355 83.760 212.580 83.930 ;
        RECT 212.770 83.780 213.020 84.580 ;
        RECT 213.190 83.780 213.530 84.410 ;
        RECT 213.700 83.855 213.990 84.580 ;
        RECT 210.895 83.390 211.225 83.590 ;
        RECT 211.395 83.390 211.725 83.590 ;
        RECT 211.895 83.390 212.315 83.590 ;
        RECT 212.490 83.420 213.185 83.590 ;
        RECT 212.490 83.170 212.660 83.420 ;
        RECT 213.355 83.170 213.530 83.780 ;
        RECT 214.160 83.780 214.500 84.410 ;
        RECT 214.670 83.780 214.920 84.580 ;
        RECT 215.110 83.930 215.440 84.410 ;
        RECT 215.610 84.120 215.835 84.580 ;
        RECT 216.005 83.930 216.335 84.410 ;
        RECT 210.225 83.000 212.660 83.170 ;
        RECT 210.225 82.200 210.555 83.000 ;
        RECT 210.725 82.030 211.055 82.830 ;
        RECT 211.355 82.200 211.685 83.000 ;
        RECT 212.330 82.030 212.580 82.830 ;
        RECT 212.850 82.030 213.020 83.170 ;
        RECT 213.190 82.200 213.530 83.170 ;
        RECT 213.700 82.030 213.990 83.195 ;
        RECT 214.160 83.170 214.335 83.780 ;
        RECT 215.110 83.760 216.335 83.930 ;
        RECT 216.965 83.800 217.465 84.410 ;
        RECT 217.840 84.035 223.185 84.580 ;
        RECT 214.505 83.420 215.200 83.590 ;
        RECT 215.030 83.170 215.200 83.420 ;
        RECT 215.375 83.390 215.795 83.590 ;
        RECT 215.965 83.390 216.295 83.590 ;
        RECT 216.465 83.390 216.795 83.590 ;
        RECT 216.965 83.170 217.135 83.800 ;
        RECT 217.320 83.340 217.670 83.590 ;
        RECT 219.425 83.205 219.765 84.035 ;
        RECT 223.360 83.810 226.870 84.580 ;
        RECT 227.045 83.815 227.500 84.580 ;
        RECT 227.775 84.200 229.075 84.410 ;
        RECT 229.330 84.220 229.660 84.580 ;
        RECT 228.905 84.050 229.075 84.200 ;
        RECT 229.830 84.080 230.090 84.410 ;
        RECT 214.160 82.200 214.500 83.170 ;
        RECT 214.670 82.030 214.840 83.170 ;
        RECT 215.030 83.000 217.465 83.170 ;
        RECT 215.110 82.030 215.360 82.830 ;
        RECT 216.005 82.200 216.335 83.000 ;
        RECT 216.635 82.030 216.965 82.830 ;
        RECT 217.135 82.200 217.465 83.000 ;
        RECT 221.245 82.465 221.595 83.715 ;
        RECT 223.360 83.290 225.010 83.810 ;
        RECT 225.180 83.120 226.870 83.640 ;
        RECT 227.975 83.590 228.195 83.990 ;
        RECT 227.040 83.390 227.530 83.590 ;
        RECT 227.720 83.380 228.195 83.590 ;
        RECT 228.440 83.590 228.650 83.990 ;
        RECT 228.905 83.925 229.660 84.050 ;
        RECT 228.905 83.880 229.750 83.925 ;
        RECT 229.480 83.760 229.750 83.880 ;
        RECT 228.440 83.380 228.770 83.590 ;
        RECT 228.940 83.320 229.350 83.625 ;
        RECT 217.840 82.030 223.185 82.465 ;
        RECT 223.360 82.030 226.870 83.120 ;
        RECT 227.045 83.150 228.220 83.210 ;
        RECT 229.580 83.185 229.750 83.760 ;
        RECT 229.550 83.150 229.750 83.185 ;
        RECT 227.045 83.040 229.750 83.150 ;
        RECT 227.045 82.420 227.300 83.040 ;
        RECT 227.890 82.980 229.690 83.040 ;
        RECT 227.890 82.950 228.220 82.980 ;
        RECT 229.920 82.880 230.090 84.080 ;
        RECT 230.260 84.035 235.605 84.580 ;
        RECT 231.845 83.205 232.185 84.035 ;
        RECT 235.780 83.810 239.290 84.580 ;
        RECT 239.460 83.855 239.750 84.580 ;
        RECT 240.910 84.180 241.240 84.580 ;
        RECT 241.410 84.010 241.580 84.280 ;
        RECT 241.750 84.180 242.080 84.580 ;
        RECT 242.250 84.010 242.505 84.280 ;
        RECT 227.550 82.780 227.735 82.870 ;
        RECT 228.325 82.780 229.160 82.790 ;
        RECT 227.550 82.580 229.160 82.780 ;
        RECT 227.550 82.540 227.780 82.580 ;
        RECT 227.045 82.200 227.380 82.420 ;
        RECT 228.385 82.030 228.740 82.410 ;
        RECT 228.910 82.200 229.160 82.580 ;
        RECT 229.410 82.030 229.660 82.810 ;
        RECT 229.830 82.200 230.090 82.880 ;
        RECT 233.665 82.465 234.015 83.715 ;
        RECT 235.780 83.290 237.430 83.810 ;
        RECT 237.600 83.120 239.290 83.640 ;
        RECT 230.260 82.030 235.605 82.465 ;
        RECT 235.780 82.030 239.290 83.120 ;
        RECT 239.460 82.030 239.750 83.195 ;
        RECT 240.840 83.000 241.110 84.010 ;
        RECT 241.280 83.840 242.505 84.010 ;
        RECT 242.700 84.080 242.955 84.410 ;
        RECT 243.170 84.100 243.500 84.580 ;
        RECT 243.670 84.160 245.205 84.410 ;
        RECT 242.700 84.000 242.885 84.080 ;
        RECT 241.280 83.170 241.450 83.840 ;
        RECT 241.620 83.340 242.000 83.670 ;
        RECT 242.170 83.340 242.505 83.670 ;
        RECT 241.280 83.000 241.595 83.170 ;
        RECT 240.845 82.030 241.160 82.830 ;
        RECT 241.425 82.385 241.595 83.000 ;
        RECT 241.765 82.660 242.000 83.340 ;
        RECT 242.170 82.385 242.505 83.170 ;
        RECT 241.425 82.215 242.505 82.385 ;
        RECT 242.700 82.870 242.870 84.000 ;
        RECT 243.670 83.930 243.840 84.160 ;
        RECT 243.040 83.760 243.840 83.930 ;
        RECT 243.040 83.210 243.210 83.760 ;
        RECT 244.020 83.590 244.305 83.990 ;
        RECT 243.440 83.390 243.805 83.590 ;
        RECT 243.975 83.390 244.305 83.590 ;
        RECT 244.575 83.590 244.855 83.990 ;
        RECT 245.035 83.930 245.205 84.160 ;
        RECT 245.430 84.100 245.760 84.580 ;
        RECT 245.930 83.930 246.100 84.410 ;
        RECT 245.035 83.760 246.100 83.930 ;
        RECT 246.360 83.920 246.625 84.580 ;
        RECT 246.795 83.950 247.040 84.410 ;
        RECT 247.215 84.085 247.545 84.580 ;
        RECT 246.795 83.740 246.965 83.950 ;
        RECT 247.735 83.900 247.945 84.360 ;
        RECT 244.575 83.390 245.050 83.590 ;
        RECT 245.220 83.390 245.665 83.590 ;
        RECT 245.835 83.380 246.185 83.590 ;
        RECT 246.360 83.220 246.965 83.740 ;
        RECT 243.040 83.040 246.100 83.210 ;
        RECT 242.700 82.200 242.955 82.870 ;
        RECT 243.125 82.030 243.455 82.790 ;
        RECT 243.625 82.630 245.260 82.870 ;
        RECT 243.625 82.200 243.875 82.630 ;
        RECT 245.030 82.540 245.260 82.630 ;
        RECT 244.045 82.030 244.400 82.450 ;
        RECT 244.590 82.370 244.920 82.410 ;
        RECT 245.430 82.370 245.760 82.870 ;
        RECT 244.590 82.200 245.760 82.370 ;
        RECT 245.930 82.200 246.100 83.040 ;
        RECT 246.360 82.030 246.625 83.040 ;
        RECT 246.795 82.880 246.965 83.220 ;
        RECT 247.135 83.240 247.365 83.670 ;
        RECT 247.535 83.420 247.945 83.900 ;
        RECT 248.115 84.095 248.900 84.360 ;
        RECT 248.115 83.240 248.370 84.095 ;
        RECT 249.100 83.650 249.375 84.360 ;
        RECT 249.600 84.090 249.870 84.580 ;
        RECT 250.130 84.030 250.300 84.410 ;
        RECT 250.515 84.200 250.845 84.580 ;
        RECT 248.540 83.420 249.375 83.650 ;
        RECT 247.135 83.070 248.905 83.240 ;
        RECT 246.795 82.870 247.050 82.880 ;
        RECT 246.795 82.200 247.080 82.870 ;
        RECT 247.280 82.030 247.495 82.875 ;
        RECT 247.755 82.775 247.945 83.070 ;
        RECT 248.170 82.710 248.500 82.900 ;
        RECT 247.665 82.200 248.140 82.540 ;
        RECT 248.310 82.535 248.500 82.710 ;
        RECT 248.670 82.705 248.905 83.070 ;
        RECT 249.100 82.760 249.375 83.420 ;
        RECT 249.545 83.340 249.810 83.920 ;
        RECT 250.130 83.860 250.845 84.030 ;
        RECT 250.040 83.310 250.395 83.680 ;
        RECT 250.675 83.670 250.845 83.860 ;
        RECT 251.015 83.835 251.270 84.410 ;
        RECT 250.675 83.340 250.930 83.670 ;
        RECT 250.675 83.130 250.845 83.340 ;
        RECT 248.310 82.030 248.925 82.535 ;
        RECT 249.555 82.030 249.870 83.090 ;
        RECT 250.130 82.960 250.845 83.130 ;
        RECT 251.100 83.105 251.270 83.835 ;
        RECT 251.445 83.740 251.705 84.580 ;
        RECT 251.885 84.180 252.220 84.580 ;
        RECT 252.390 84.010 252.595 84.410 ;
        RECT 252.805 84.100 253.080 84.580 ;
        RECT 253.290 84.080 253.550 84.410 ;
        RECT 251.910 83.840 252.595 84.010 ;
        RECT 250.130 82.200 250.300 82.960 ;
        RECT 250.515 82.030 250.845 82.790 ;
        RECT 251.015 82.200 251.270 83.105 ;
        RECT 251.445 82.030 251.705 83.180 ;
        RECT 251.910 82.810 252.250 83.840 ;
        RECT 252.420 83.170 252.670 83.670 ;
        RECT 252.850 83.340 253.210 83.920 ;
        RECT 253.380 83.170 253.550 84.080 ;
        RECT 253.720 83.810 257.230 84.580 ;
        RECT 257.400 83.830 258.610 84.580 ;
        RECT 253.720 83.290 255.370 83.810 ;
        RECT 252.420 83.000 253.550 83.170 ;
        RECT 255.540 83.120 257.230 83.640 ;
        RECT 257.400 83.290 257.920 83.830 ;
        RECT 258.785 83.815 259.240 84.580 ;
        RECT 259.515 84.200 260.815 84.410 ;
        RECT 261.070 84.220 261.400 84.580 ;
        RECT 260.645 84.050 260.815 84.200 ;
        RECT 261.570 84.080 261.830 84.410 ;
        RECT 262.010 84.080 262.340 84.580 ;
        RECT 258.090 83.120 258.610 83.660 ;
        RECT 259.715 83.590 259.935 83.990 ;
        RECT 258.780 83.390 259.270 83.590 ;
        RECT 259.460 83.380 259.935 83.590 ;
        RECT 260.180 83.590 260.390 83.990 ;
        RECT 260.645 83.925 261.400 84.050 ;
        RECT 260.645 83.880 261.490 83.925 ;
        RECT 261.220 83.760 261.490 83.880 ;
        RECT 260.180 83.380 260.510 83.590 ;
        RECT 260.680 83.320 261.090 83.625 ;
        RECT 251.910 82.635 252.575 82.810 ;
        RECT 251.885 82.030 252.220 82.455 ;
        RECT 252.390 82.230 252.575 82.635 ;
        RECT 252.780 82.030 253.110 82.810 ;
        RECT 253.280 82.230 253.550 83.000 ;
        RECT 253.720 82.030 257.230 83.120 ;
        RECT 257.400 82.030 258.610 83.120 ;
        RECT 258.785 83.150 259.960 83.210 ;
        RECT 261.320 83.185 261.490 83.760 ;
        RECT 261.290 83.150 261.490 83.185 ;
        RECT 258.785 83.040 261.490 83.150 ;
        RECT 258.785 82.420 259.040 83.040 ;
        RECT 259.630 82.980 261.430 83.040 ;
        RECT 259.630 82.950 259.960 82.980 ;
        RECT 261.660 82.880 261.830 84.080 ;
        RECT 262.540 84.010 262.710 84.360 ;
        RECT 262.910 84.180 263.240 84.580 ;
        RECT 263.410 84.010 263.580 84.360 ;
        RECT 263.750 84.180 264.130 84.580 ;
        RECT 262.005 83.340 262.355 83.910 ;
        RECT 262.540 83.840 264.150 84.010 ;
        RECT 264.320 83.905 264.590 84.250 ;
        RECT 263.980 83.670 264.150 83.840 ;
        RECT 259.290 82.780 259.475 82.870 ;
        RECT 260.065 82.780 260.900 82.790 ;
        RECT 259.290 82.580 260.900 82.780 ;
        RECT 259.290 82.540 259.520 82.580 ;
        RECT 258.785 82.200 259.120 82.420 ;
        RECT 260.125 82.030 260.480 82.410 ;
        RECT 260.650 82.200 260.900 82.580 ;
        RECT 261.150 82.030 261.400 82.810 ;
        RECT 261.570 82.200 261.830 82.880 ;
        RECT 262.005 82.880 262.325 83.170 ;
        RECT 262.525 83.050 263.235 83.670 ;
        RECT 263.405 83.340 263.810 83.670 ;
        RECT 263.980 83.340 264.250 83.670 ;
        RECT 263.980 83.170 264.150 83.340 ;
        RECT 264.420 83.170 264.590 83.905 ;
        RECT 265.220 83.855 265.510 84.580 ;
        RECT 265.680 84.120 266.240 84.410 ;
        RECT 266.410 84.120 266.660 84.580 ;
        RECT 263.425 83.000 264.150 83.170 ;
        RECT 263.425 82.880 263.595 83.000 ;
        RECT 262.005 82.710 263.595 82.880 ;
        RECT 262.005 82.250 263.660 82.540 ;
        RECT 263.830 82.030 264.110 82.830 ;
        RECT 264.320 82.200 264.590 83.170 ;
        RECT 265.220 82.030 265.510 83.195 ;
        RECT 265.680 82.750 265.930 84.120 ;
        RECT 267.280 83.950 267.610 84.310 ;
        RECT 267.980 84.035 273.325 84.580 ;
        RECT 273.500 84.035 278.845 84.580 ;
        RECT 279.020 84.035 284.365 84.580 ;
        RECT 266.220 83.760 267.610 83.950 ;
        RECT 266.220 83.670 266.390 83.760 ;
        RECT 266.100 83.340 266.390 83.670 ;
        RECT 266.560 83.340 266.900 83.590 ;
        RECT 267.120 83.340 267.795 83.590 ;
        RECT 266.220 83.090 266.390 83.340 ;
        RECT 266.220 82.920 267.160 83.090 ;
        RECT 267.530 82.980 267.795 83.340 ;
        RECT 269.565 83.205 269.905 84.035 ;
        RECT 265.680 82.200 266.140 82.750 ;
        RECT 266.330 82.030 266.660 82.750 ;
        RECT 266.860 82.370 267.160 82.920 ;
        RECT 267.330 82.030 267.610 82.700 ;
        RECT 271.385 82.465 271.735 83.715 ;
        RECT 275.085 83.205 275.425 84.035 ;
        RECT 276.905 82.465 277.255 83.715 ;
        RECT 280.605 83.205 280.945 84.035 ;
        RECT 284.540 83.810 287.130 84.580 ;
        RECT 287.770 84.090 288.100 84.580 ;
        RECT 288.270 83.985 288.890 84.410 ;
        RECT 282.425 82.465 282.775 83.715 ;
        RECT 284.540 83.290 285.750 83.810 ;
        RECT 285.920 83.120 287.130 83.640 ;
        RECT 287.760 83.340 288.100 83.920 ;
        RECT 288.270 83.650 288.630 83.985 ;
        RECT 289.350 83.890 289.680 84.580 ;
        RECT 290.980 83.855 291.270 84.580 ;
        RECT 291.440 83.810 294.030 84.580 ;
        RECT 294.665 84.030 294.920 84.320 ;
        RECT 295.090 84.200 295.420 84.580 ;
        RECT 294.665 83.860 295.415 84.030 ;
        RECT 288.270 83.370 289.690 83.650 ;
        RECT 267.980 82.030 273.325 82.465 ;
        RECT 273.500 82.030 278.845 82.465 ;
        RECT 279.020 82.030 284.365 82.465 ;
        RECT 284.540 82.030 287.130 83.120 ;
        RECT 287.770 82.030 288.100 83.170 ;
        RECT 288.270 82.200 288.630 83.370 ;
        RECT 288.830 82.030 289.160 83.200 ;
        RECT 289.360 82.200 289.690 83.370 ;
        RECT 291.440 83.290 292.650 83.810 ;
        RECT 289.890 82.030 290.220 83.200 ;
        RECT 290.980 82.030 291.270 83.195 ;
        RECT 292.820 83.120 294.030 83.640 ;
        RECT 291.440 82.030 294.030 83.120 ;
        RECT 294.665 83.040 295.015 83.690 ;
        RECT 295.185 82.870 295.415 83.860 ;
        RECT 294.665 82.700 295.415 82.870 ;
        RECT 294.665 82.200 294.920 82.700 ;
        RECT 295.090 82.030 295.420 82.530 ;
        RECT 295.590 82.200 295.760 84.320 ;
        RECT 296.120 84.220 296.450 84.580 ;
        RECT 296.620 84.190 297.115 84.360 ;
        RECT 297.320 84.190 298.175 84.360 ;
        RECT 295.990 83.000 296.450 84.050 ;
        RECT 295.930 82.215 296.255 83.000 ;
        RECT 296.620 82.830 296.790 84.190 ;
        RECT 296.960 83.280 297.310 83.900 ;
        RECT 297.480 83.680 297.835 83.900 ;
        RECT 297.480 83.090 297.650 83.680 ;
        RECT 298.005 83.480 298.175 84.190 ;
        RECT 299.050 84.120 299.380 84.580 ;
        RECT 299.590 84.220 299.940 84.390 ;
        RECT 298.380 83.650 299.170 83.900 ;
        RECT 299.590 83.830 299.850 84.220 ;
        RECT 300.160 84.130 301.110 84.410 ;
        RECT 301.280 84.140 301.470 84.580 ;
        RECT 301.640 84.200 302.710 84.370 ;
        RECT 299.340 83.480 299.510 83.660 ;
        RECT 296.620 82.660 297.015 82.830 ;
        RECT 297.185 82.700 297.650 83.090 ;
        RECT 297.820 83.310 299.510 83.480 ;
        RECT 296.845 82.530 297.015 82.660 ;
        RECT 297.820 82.530 297.990 83.310 ;
        RECT 299.680 83.140 299.850 83.830 ;
        RECT 298.350 82.970 299.850 83.140 ;
        RECT 300.040 83.170 300.250 83.960 ;
        RECT 300.420 83.340 300.770 83.960 ;
        RECT 300.940 83.350 301.110 84.130 ;
        RECT 301.640 83.970 301.810 84.200 ;
        RECT 301.280 83.800 301.810 83.970 ;
        RECT 301.280 83.520 301.500 83.800 ;
        RECT 301.980 83.630 302.220 84.030 ;
        RECT 300.940 83.180 301.345 83.350 ;
        RECT 301.680 83.260 302.220 83.630 ;
        RECT 302.390 83.845 302.710 84.200 ;
        RECT 302.955 84.120 303.260 84.580 ;
        RECT 303.430 83.870 303.685 84.400 ;
        RECT 302.390 83.670 302.715 83.845 ;
        RECT 302.390 83.370 303.305 83.670 ;
        RECT 302.565 83.340 303.305 83.370 ;
        RECT 300.040 83.010 300.715 83.170 ;
        RECT 301.175 83.090 301.345 83.180 ;
        RECT 300.040 83.000 301.005 83.010 ;
        RECT 299.680 82.830 299.850 82.970 ;
        RECT 296.425 82.030 296.675 82.490 ;
        RECT 296.845 82.200 297.095 82.530 ;
        RECT 297.310 82.200 297.990 82.530 ;
        RECT 298.160 82.630 299.235 82.800 ;
        RECT 299.680 82.660 300.240 82.830 ;
        RECT 300.545 82.710 301.005 83.000 ;
        RECT 301.175 82.920 302.395 83.090 ;
        RECT 298.160 82.290 298.330 82.630 ;
        RECT 298.565 82.030 298.895 82.460 ;
        RECT 299.065 82.290 299.235 82.630 ;
        RECT 299.530 82.030 299.900 82.490 ;
        RECT 300.070 82.200 300.240 82.660 ;
        RECT 301.175 82.540 301.345 82.920 ;
        RECT 302.565 82.750 302.735 83.340 ;
        RECT 303.475 83.220 303.685 83.870 ;
        RECT 300.475 82.200 301.345 82.540 ;
        RECT 301.935 82.580 302.735 82.750 ;
        RECT 301.515 82.030 301.765 82.490 ;
        RECT 301.935 82.290 302.105 82.580 ;
        RECT 302.285 82.030 302.615 82.410 ;
        RECT 302.955 82.030 303.260 83.170 ;
        RECT 303.430 82.340 303.685 83.220 ;
        RECT 303.865 83.840 304.120 84.410 ;
        RECT 304.290 84.180 304.620 84.580 ;
        RECT 305.045 84.045 305.575 84.410 ;
        RECT 305.045 84.010 305.220 84.045 ;
        RECT 304.290 83.840 305.220 84.010 ;
        RECT 305.765 83.900 306.040 84.410 ;
        RECT 303.865 83.170 304.035 83.840 ;
        RECT 304.290 83.670 304.460 83.840 ;
        RECT 304.205 83.340 304.460 83.670 ;
        RECT 304.685 83.340 304.880 83.670 ;
        RECT 303.865 82.200 304.200 83.170 ;
        RECT 304.370 82.030 304.540 83.170 ;
        RECT 304.710 82.370 304.880 83.340 ;
        RECT 305.050 82.710 305.220 83.840 ;
        RECT 305.390 83.050 305.560 83.850 ;
        RECT 305.760 83.730 306.040 83.900 ;
        RECT 305.765 83.250 306.040 83.730 ;
        RECT 306.210 83.050 306.400 84.410 ;
        RECT 306.580 84.045 307.090 84.580 ;
        RECT 307.310 83.770 307.555 84.375 ;
        RECT 308.000 83.810 309.670 84.580 ;
        RECT 309.840 83.830 311.050 84.580 ;
        RECT 306.600 83.600 307.830 83.770 ;
        RECT 305.390 82.880 306.400 83.050 ;
        RECT 306.570 83.035 307.320 83.225 ;
        RECT 305.050 82.540 306.175 82.710 ;
        RECT 306.570 82.370 306.740 83.035 ;
        RECT 307.490 82.790 307.830 83.600 ;
        RECT 308.000 83.290 308.750 83.810 ;
        RECT 308.920 83.120 309.670 83.640 ;
        RECT 304.710 82.200 306.740 82.370 ;
        RECT 306.910 82.030 307.080 82.790 ;
        RECT 307.315 82.380 307.830 82.790 ;
        RECT 308.000 82.030 309.670 83.120 ;
        RECT 309.840 83.120 310.360 83.660 ;
        RECT 310.530 83.290 311.050 83.830 ;
        RECT 309.840 82.030 311.050 83.120 ;
        RECT 162.095 81.860 311.135 82.030 ;
        RECT 162.180 80.770 163.390 81.860 ;
        RECT 163.560 80.770 165.230 81.860 ;
        RECT 162.180 80.060 162.700 80.600 ;
        RECT 162.870 80.230 163.390 80.770 ;
        RECT 163.560 80.080 164.310 80.600 ;
        RECT 164.480 80.250 165.230 80.770 ;
        RECT 165.865 80.670 166.120 81.550 ;
        RECT 166.290 80.720 166.595 81.860 ;
        RECT 166.935 81.480 167.265 81.860 ;
        RECT 167.445 81.310 167.615 81.600 ;
        RECT 167.785 81.400 168.035 81.860 ;
        RECT 166.815 81.140 167.615 81.310 ;
        RECT 168.205 81.350 169.075 81.690 ;
        RECT 162.180 79.310 163.390 80.060 ;
        RECT 163.560 79.310 165.230 80.080 ;
        RECT 165.865 80.020 166.075 80.670 ;
        RECT 166.815 80.550 166.985 81.140 ;
        RECT 168.205 80.970 168.375 81.350 ;
        RECT 169.310 81.230 169.480 81.690 ;
        RECT 169.650 81.400 170.020 81.860 ;
        RECT 170.315 81.260 170.485 81.600 ;
        RECT 170.655 81.430 170.985 81.860 ;
        RECT 171.220 81.260 171.390 81.600 ;
        RECT 167.155 80.800 168.375 80.970 ;
        RECT 168.545 80.890 169.005 81.180 ;
        RECT 169.310 81.060 169.870 81.230 ;
        RECT 170.315 81.090 171.390 81.260 ;
        RECT 171.560 81.360 172.240 81.690 ;
        RECT 172.455 81.360 172.705 81.690 ;
        RECT 172.875 81.400 173.125 81.860 ;
        RECT 169.700 80.920 169.870 81.060 ;
        RECT 168.545 80.880 169.510 80.890 ;
        RECT 168.205 80.710 168.375 80.800 ;
        RECT 168.835 80.720 169.510 80.880 ;
        RECT 166.245 80.520 166.985 80.550 ;
        RECT 166.245 80.220 167.160 80.520 ;
        RECT 166.835 80.045 167.160 80.220 ;
        RECT 165.865 79.490 166.120 80.020 ;
        RECT 166.290 79.310 166.595 79.770 ;
        RECT 166.840 79.690 167.160 80.045 ;
        RECT 167.330 80.260 167.870 80.630 ;
        RECT 168.205 80.540 168.610 80.710 ;
        RECT 167.330 79.860 167.570 80.260 ;
        RECT 168.050 80.090 168.270 80.370 ;
        RECT 167.740 79.920 168.270 80.090 ;
        RECT 167.740 79.690 167.910 79.920 ;
        RECT 168.440 79.760 168.610 80.540 ;
        RECT 168.780 79.930 169.130 80.550 ;
        RECT 169.300 79.930 169.510 80.720 ;
        RECT 169.700 80.750 171.200 80.920 ;
        RECT 169.700 80.060 169.870 80.750 ;
        RECT 171.560 80.580 171.730 81.360 ;
        RECT 172.535 81.230 172.705 81.360 ;
        RECT 170.040 80.410 171.730 80.580 ;
        RECT 171.900 80.800 172.365 81.190 ;
        RECT 172.535 81.060 172.930 81.230 ;
        RECT 170.040 80.230 170.210 80.410 ;
        RECT 166.840 79.520 167.910 79.690 ;
        RECT 168.080 79.310 168.270 79.750 ;
        RECT 168.440 79.480 169.390 79.760 ;
        RECT 169.700 79.670 169.960 80.060 ;
        RECT 170.380 79.990 171.170 80.240 ;
        RECT 169.610 79.500 169.960 79.670 ;
        RECT 170.170 79.310 170.500 79.770 ;
        RECT 171.375 79.700 171.545 80.410 ;
        RECT 171.900 80.210 172.070 80.800 ;
        RECT 171.715 79.990 172.070 80.210 ;
        RECT 172.240 79.990 172.590 80.610 ;
        RECT 172.760 79.700 172.930 81.060 ;
        RECT 173.295 80.890 173.620 81.675 ;
        RECT 173.100 79.840 173.560 80.890 ;
        RECT 171.375 79.530 172.230 79.700 ;
        RECT 172.435 79.530 172.930 79.700 ;
        RECT 173.100 79.310 173.430 79.670 ;
        RECT 173.790 79.570 173.960 81.690 ;
        RECT 174.130 81.360 174.460 81.860 ;
        RECT 174.630 81.190 174.885 81.690 ;
        RECT 174.135 81.020 174.885 81.190 ;
        RECT 174.135 80.030 174.365 81.020 ;
        RECT 174.535 80.200 174.885 80.850 ;
        RECT 175.060 80.695 175.350 81.860 ;
        RECT 175.520 80.770 179.030 81.860 ;
        RECT 179.200 80.770 180.410 81.860 ;
        RECT 175.520 80.080 177.170 80.600 ;
        RECT 177.340 80.250 179.030 80.770 ;
        RECT 174.135 79.860 174.885 80.030 ;
        RECT 174.130 79.310 174.460 79.690 ;
        RECT 174.630 79.570 174.885 79.860 ;
        RECT 175.060 79.310 175.350 80.035 ;
        RECT 175.520 79.310 179.030 80.080 ;
        RECT 179.200 80.060 179.720 80.600 ;
        RECT 179.890 80.230 180.410 80.770 ;
        RECT 180.585 80.720 180.920 81.690 ;
        RECT 181.090 80.720 181.260 81.860 ;
        RECT 181.430 81.520 183.460 81.690 ;
        RECT 179.200 79.310 180.410 80.060 ;
        RECT 180.585 80.050 180.755 80.720 ;
        RECT 181.430 80.550 181.600 81.520 ;
        RECT 180.925 80.220 181.180 80.550 ;
        RECT 181.405 80.220 181.600 80.550 ;
        RECT 181.770 81.180 182.895 81.350 ;
        RECT 181.010 80.050 181.180 80.220 ;
        RECT 181.770 80.050 181.940 81.180 ;
        RECT 180.585 79.480 180.840 80.050 ;
        RECT 181.010 79.880 181.940 80.050 ;
        RECT 182.110 80.840 183.120 81.010 ;
        RECT 182.110 80.040 182.280 80.840 ;
        RECT 182.485 80.160 182.760 80.640 ;
        RECT 182.480 79.990 182.760 80.160 ;
        RECT 181.765 79.845 181.940 79.880 ;
        RECT 181.010 79.310 181.340 79.710 ;
        RECT 181.765 79.480 182.295 79.845 ;
        RECT 182.485 79.480 182.760 79.990 ;
        RECT 182.930 79.480 183.120 80.840 ;
        RECT 183.290 80.855 183.460 81.520 ;
        RECT 183.630 81.100 183.800 81.860 ;
        RECT 184.035 81.100 184.550 81.510 ;
        RECT 184.720 81.425 190.065 81.860 ;
        RECT 183.290 80.665 184.040 80.855 ;
        RECT 184.210 80.290 184.550 81.100 ;
        RECT 183.320 80.120 184.550 80.290 ;
        RECT 183.300 79.310 183.810 79.845 ;
        RECT 184.030 79.515 184.275 80.120 ;
        RECT 186.305 79.855 186.645 80.685 ;
        RECT 188.125 80.175 188.475 81.425 ;
        RECT 190.240 80.770 191.910 81.860 ;
        RECT 192.540 81.350 193.735 81.640 ;
        RECT 190.240 80.080 190.990 80.600 ;
        RECT 191.160 80.250 191.910 80.770 ;
        RECT 192.560 81.010 193.725 81.180 ;
        RECT 193.905 81.060 194.185 81.860 ;
        RECT 192.560 80.720 192.890 81.010 ;
        RECT 193.555 80.890 193.725 81.010 ;
        RECT 193.060 80.550 193.285 80.840 ;
        RECT 193.555 80.720 194.225 80.890 ;
        RECT 194.395 80.720 194.670 81.690 ;
        RECT 194.055 80.550 194.225 80.720 ;
        RECT 192.540 80.220 192.890 80.550 ;
        RECT 193.060 80.220 193.885 80.550 ;
        RECT 194.055 80.220 194.330 80.550 ;
        RECT 184.720 79.310 190.065 79.855 ;
        RECT 190.240 79.310 191.910 80.080 ;
        RECT 194.055 80.050 194.225 80.220 ;
        RECT 192.560 79.880 194.225 80.050 ;
        RECT 194.500 79.985 194.670 80.720 ;
        RECT 194.840 80.655 195.130 81.860 ;
        RECT 195.310 81.140 195.640 81.860 ;
        RECT 195.300 80.500 195.530 80.840 ;
        RECT 195.820 80.500 196.035 81.615 ;
        RECT 196.230 80.915 196.560 81.690 ;
        RECT 196.730 81.085 197.440 81.860 ;
        RECT 196.230 80.700 197.380 80.915 ;
        RECT 195.300 80.300 195.630 80.500 ;
        RECT 195.820 80.320 196.270 80.500 ;
        RECT 195.940 80.300 196.270 80.320 ;
        RECT 196.440 80.300 196.910 80.530 ;
        RECT 192.560 79.530 192.815 79.880 ;
        RECT 192.985 79.310 193.315 79.710 ;
        RECT 193.485 79.530 193.655 79.880 ;
        RECT 193.825 79.310 194.205 79.710 ;
        RECT 194.395 79.640 194.670 79.985 ;
        RECT 194.840 79.310 195.130 80.140 ;
        RECT 197.095 80.130 197.380 80.700 ;
        RECT 197.610 80.255 197.890 81.690 ;
        RECT 198.060 80.770 200.650 81.860 ;
        RECT 195.300 79.940 196.480 80.130 ;
        RECT 195.300 79.480 195.640 79.940 ;
        RECT 196.150 79.860 196.480 79.940 ;
        RECT 196.670 79.940 197.380 80.130 ;
        RECT 196.670 79.800 196.970 79.940 ;
        RECT 196.655 79.790 196.970 79.800 ;
        RECT 196.645 79.780 196.970 79.790 ;
        RECT 196.635 79.775 196.970 79.780 ;
        RECT 195.810 79.310 195.980 79.770 ;
        RECT 196.630 79.765 196.970 79.775 ;
        RECT 196.625 79.760 196.970 79.765 ;
        RECT 196.620 79.750 196.970 79.760 ;
        RECT 196.615 79.745 196.970 79.750 ;
        RECT 196.610 79.480 196.970 79.745 ;
        RECT 197.210 79.310 197.380 79.770 ;
        RECT 197.550 79.480 197.890 80.255 ;
        RECT 198.060 80.080 199.270 80.600 ;
        RECT 199.440 80.250 200.650 80.770 ;
        RECT 200.820 80.695 201.110 81.860 ;
        RECT 201.280 80.890 201.550 81.660 ;
        RECT 201.720 81.080 202.050 81.860 ;
        RECT 202.255 81.255 202.440 81.660 ;
        RECT 202.610 81.435 202.945 81.860 ;
        RECT 202.255 81.080 202.920 81.255 ;
        RECT 201.280 80.720 202.410 80.890 ;
        RECT 198.060 79.310 200.650 80.080 ;
        RECT 200.820 79.310 201.110 80.035 ;
        RECT 201.280 79.810 201.450 80.720 ;
        RECT 201.620 79.970 201.980 80.550 ;
        RECT 202.160 80.220 202.410 80.720 ;
        RECT 202.580 80.050 202.920 81.080 ;
        RECT 204.065 80.850 204.360 81.690 ;
        RECT 204.530 81.020 204.780 81.860 ;
        RECT 204.950 81.190 205.200 81.690 ;
        RECT 205.370 81.360 205.620 81.860 ;
        RECT 205.790 81.190 206.040 81.690 ;
        RECT 206.210 81.360 206.460 81.860 ;
        RECT 206.730 81.520 210.340 81.690 ;
        RECT 206.730 81.360 206.980 81.520 ;
        RECT 207.570 81.360 207.820 81.520 ;
        RECT 207.150 81.190 207.400 81.350 ;
        RECT 207.990 81.190 208.240 81.350 ;
        RECT 204.950 81.020 208.240 81.190 ;
        RECT 208.410 81.020 208.660 81.520 ;
        RECT 208.830 80.850 209.080 81.350 ;
        RECT 209.250 81.020 209.500 81.520 ;
        RECT 209.670 80.850 209.920 81.350 ;
        RECT 210.090 81.020 210.340 81.520 ;
        RECT 210.510 80.850 210.715 81.640 ;
        RECT 204.065 80.680 208.660 80.850 ;
        RECT 208.830 80.680 210.715 80.850 ;
        RECT 204.065 80.300 204.400 80.510 ;
        RECT 204.570 80.130 204.740 80.680 ;
        RECT 208.490 80.510 208.660 80.680 ;
        RECT 204.990 80.300 206.645 80.510 ;
        RECT 206.990 80.300 208.255 80.510 ;
        RECT 208.490 80.300 210.080 80.510 ;
        RECT 210.375 80.130 210.715 80.680 ;
        RECT 202.235 79.880 202.920 80.050 ;
        RECT 204.065 79.960 204.740 80.130 ;
        RECT 201.280 79.480 201.540 79.810 ;
        RECT 201.750 79.310 202.025 79.790 ;
        RECT 202.235 79.480 202.440 79.880 ;
        RECT 202.610 79.310 202.945 79.710 ;
        RECT 204.065 79.480 204.400 79.960 ;
        RECT 204.910 79.950 210.715 80.130 ;
        RECT 204.570 79.310 204.740 79.780 ;
        RECT 204.910 79.480 205.240 79.950 ;
        RECT 205.410 79.310 205.580 79.780 ;
        RECT 205.750 79.480 206.080 79.950 ;
        RECT 206.250 79.310 206.940 79.780 ;
        RECT 207.110 79.480 207.440 79.950 ;
        RECT 207.610 79.310 207.780 79.780 ;
        RECT 207.950 79.480 208.280 79.950 ;
        RECT 208.450 79.310 208.620 79.780 ;
        RECT 208.790 79.480 209.120 79.950 ;
        RECT 209.290 79.310 209.460 79.780 ;
        RECT 209.630 79.480 209.960 79.950 ;
        RECT 210.130 79.310 210.300 79.780 ;
        RECT 210.470 79.540 210.715 79.950 ;
        RECT 210.995 80.850 211.200 81.640 ;
        RECT 211.370 81.520 214.980 81.690 ;
        RECT 211.370 81.020 211.620 81.520 ;
        RECT 211.790 80.850 212.040 81.350 ;
        RECT 212.210 81.020 212.460 81.520 ;
        RECT 212.630 80.850 212.880 81.350 ;
        RECT 213.050 81.020 213.300 81.520 ;
        RECT 213.890 81.360 214.140 81.520 ;
        RECT 214.730 81.360 214.980 81.520 ;
        RECT 215.250 81.360 215.500 81.860 ;
        RECT 213.470 81.190 213.720 81.350 ;
        RECT 214.310 81.190 214.560 81.350 ;
        RECT 215.670 81.190 215.920 81.690 ;
        RECT 216.090 81.360 216.340 81.860 ;
        RECT 216.510 81.190 216.760 81.690 ;
        RECT 213.470 81.020 216.760 81.190 ;
        RECT 216.930 81.020 217.180 81.860 ;
        RECT 217.350 80.850 217.645 81.690 ;
        RECT 217.840 81.425 223.185 81.860 ;
        RECT 210.995 80.680 212.880 80.850 ;
        RECT 213.050 80.680 217.645 80.850 ;
        RECT 210.995 80.130 211.335 80.680 ;
        RECT 213.050 80.510 213.220 80.680 ;
        RECT 211.630 80.300 213.220 80.510 ;
        RECT 213.455 80.300 214.720 80.510 ;
        RECT 215.065 80.300 216.720 80.510 ;
        RECT 216.970 80.130 217.140 80.680 ;
        RECT 217.310 80.300 217.645 80.510 ;
        RECT 210.995 79.950 216.800 80.130 ;
        RECT 216.970 79.960 217.645 80.130 ;
        RECT 210.995 79.540 211.240 79.950 ;
        RECT 211.410 79.310 211.580 79.780 ;
        RECT 211.750 79.480 212.080 79.950 ;
        RECT 212.250 79.310 212.420 79.780 ;
        RECT 212.590 79.480 212.920 79.950 ;
        RECT 213.090 79.310 213.260 79.780 ;
        RECT 213.430 79.480 213.760 79.950 ;
        RECT 213.930 79.310 214.100 79.780 ;
        RECT 214.270 79.480 214.600 79.950 ;
        RECT 214.770 79.310 215.460 79.780 ;
        RECT 215.630 79.480 215.960 79.950 ;
        RECT 216.130 79.310 216.300 79.780 ;
        RECT 216.470 79.480 216.800 79.950 ;
        RECT 216.970 79.310 217.140 79.780 ;
        RECT 217.310 79.480 217.645 79.960 ;
        RECT 219.425 79.855 219.765 80.685 ;
        RECT 221.245 80.175 221.595 81.425 ;
        RECT 223.820 81.355 224.450 81.860 ;
        RECT 223.835 80.820 224.090 81.185 ;
        RECT 224.260 81.180 224.450 81.355 ;
        RECT 224.630 81.350 225.105 81.690 ;
        RECT 224.260 80.990 224.590 81.180 ;
        RECT 224.815 80.820 225.065 81.115 ;
        RECT 225.290 81.015 225.505 81.860 ;
        RECT 225.705 81.020 225.980 81.690 ;
        RECT 225.720 81.010 225.980 81.020 ;
        RECT 223.835 80.650 225.625 80.820 ;
        RECT 225.810 80.670 225.980 81.010 ;
        RECT 226.150 80.850 226.410 81.860 ;
        RECT 226.580 80.695 226.870 81.860 ;
        RECT 227.040 80.770 228.250 81.860 ;
        RECT 223.820 79.990 224.205 80.470 ;
        RECT 217.840 79.310 223.185 79.855 ;
        RECT 224.375 79.795 224.630 80.650 ;
        RECT 223.840 79.530 224.630 79.795 ;
        RECT 224.800 79.975 225.210 80.470 ;
        RECT 225.395 80.220 225.625 80.650 ;
        RECT 225.795 80.150 226.410 80.670 ;
        RECT 224.800 79.530 225.030 79.975 ;
        RECT 225.795 79.940 225.965 80.150 ;
        RECT 227.040 80.060 227.560 80.600 ;
        RECT 227.730 80.230 228.250 80.770 ;
        RECT 228.440 81.020 228.695 81.690 ;
        RECT 228.865 81.100 229.195 81.860 ;
        RECT 229.365 81.260 229.615 81.690 ;
        RECT 229.785 81.440 230.140 81.860 ;
        RECT 230.330 81.520 231.500 81.690 ;
        RECT 230.330 81.480 230.660 81.520 ;
        RECT 230.770 81.260 231.000 81.350 ;
        RECT 229.365 81.020 231.000 81.260 ;
        RECT 231.170 81.020 231.500 81.520 ;
        RECT 225.210 79.310 225.540 79.805 ;
        RECT 225.715 79.480 225.965 79.940 ;
        RECT 226.135 79.310 226.410 79.970 ;
        RECT 226.580 79.310 226.870 80.035 ;
        RECT 227.040 79.310 228.250 80.060 ;
        RECT 228.440 79.890 228.610 81.020 ;
        RECT 231.670 80.850 231.840 81.690 ;
        RECT 228.780 80.680 231.840 80.850 ;
        RECT 228.780 80.130 228.950 80.680 ;
        RECT 229.170 80.330 229.545 80.500 ;
        RECT 229.180 80.300 229.545 80.330 ;
        RECT 229.715 80.300 230.045 80.500 ;
        RECT 228.780 79.960 229.580 80.130 ;
        RECT 228.440 79.820 228.625 79.890 ;
        RECT 228.440 79.810 228.650 79.820 ;
        RECT 228.440 79.480 228.695 79.810 ;
        RECT 228.910 79.310 229.240 79.790 ;
        RECT 229.410 79.730 229.580 79.960 ;
        RECT 229.760 79.900 230.045 80.300 ;
        RECT 230.315 80.300 230.790 80.500 ;
        RECT 230.960 80.300 231.405 80.500 ;
        RECT 231.575 80.300 231.925 80.510 ;
        RECT 230.315 79.900 230.595 80.300 ;
        RECT 230.775 79.960 231.840 80.130 ;
        RECT 230.775 79.730 230.945 79.960 ;
        RECT 229.410 79.480 230.945 79.730 ;
        RECT 231.170 79.310 231.500 79.790 ;
        RECT 231.670 79.480 231.840 79.960 ;
        RECT 232.110 79.490 232.370 81.680 ;
        RECT 232.540 81.130 232.880 81.860 ;
        RECT 233.060 80.950 233.330 81.680 ;
        RECT 232.560 80.730 233.330 80.950 ;
        RECT 233.510 80.970 233.740 81.680 ;
        RECT 233.910 81.150 234.240 81.860 ;
        RECT 234.410 80.970 234.670 81.680 ;
        RECT 233.510 80.730 234.670 80.970 ;
        RECT 234.860 80.770 238.370 81.860 ;
        RECT 232.560 80.060 232.850 80.730 ;
        RECT 233.030 80.240 233.495 80.550 ;
        RECT 233.675 80.240 234.200 80.550 ;
        RECT 232.560 79.860 233.790 80.060 ;
        RECT 232.630 79.310 233.300 79.680 ;
        RECT 233.480 79.490 233.790 79.860 ;
        RECT 233.970 79.600 234.200 80.240 ;
        RECT 234.380 80.220 234.680 80.550 ;
        RECT 234.860 80.080 236.510 80.600 ;
        RECT 236.680 80.250 238.370 80.770 ;
        RECT 239.005 81.470 239.340 81.690 ;
        RECT 240.345 81.480 240.700 81.860 ;
        RECT 239.005 80.850 239.260 81.470 ;
        RECT 239.510 81.310 239.740 81.350 ;
        RECT 240.870 81.310 241.120 81.690 ;
        RECT 239.510 81.110 241.120 81.310 ;
        RECT 239.510 81.020 239.695 81.110 ;
        RECT 240.285 81.100 241.120 81.110 ;
        RECT 241.370 81.080 241.620 81.860 ;
        RECT 241.790 81.010 242.050 81.690 ;
        RECT 239.850 80.910 240.180 80.940 ;
        RECT 239.850 80.850 241.650 80.910 ;
        RECT 239.005 80.740 241.710 80.850 ;
        RECT 239.005 80.680 240.180 80.740 ;
        RECT 241.510 80.705 241.710 80.740 ;
        RECT 239.000 80.300 239.490 80.500 ;
        RECT 239.680 80.300 240.155 80.510 ;
        RECT 234.380 79.310 234.670 80.040 ;
        RECT 234.860 79.310 238.370 80.080 ;
        RECT 239.005 79.310 239.460 80.075 ;
        RECT 239.935 79.900 240.155 80.300 ;
        RECT 240.400 80.300 240.730 80.510 ;
        RECT 240.400 79.900 240.610 80.300 ;
        RECT 240.900 80.265 241.310 80.570 ;
        RECT 241.540 80.130 241.710 80.705 ;
        RECT 241.440 80.010 241.710 80.130 ;
        RECT 240.865 79.965 241.710 80.010 ;
        RECT 240.865 79.840 241.620 79.965 ;
        RECT 240.865 79.690 241.035 79.840 ;
        RECT 241.880 79.820 242.050 81.010 ;
        RECT 241.820 79.810 242.050 79.820 ;
        RECT 239.735 79.480 241.035 79.690 ;
        RECT 241.290 79.310 241.620 79.670 ;
        RECT 241.790 79.480 242.050 79.810 ;
        RECT 242.240 81.020 242.495 81.690 ;
        RECT 242.665 81.100 242.995 81.860 ;
        RECT 243.165 81.260 243.415 81.690 ;
        RECT 243.585 81.440 243.940 81.860 ;
        RECT 244.130 81.520 245.300 81.690 ;
        RECT 244.130 81.480 244.460 81.520 ;
        RECT 244.570 81.260 244.800 81.350 ;
        RECT 243.165 81.020 244.800 81.260 ;
        RECT 244.970 81.020 245.300 81.520 ;
        RECT 242.240 79.890 242.410 81.020 ;
        RECT 245.470 80.850 245.640 81.690 ;
        RECT 242.580 80.680 245.640 80.850 ;
        RECT 245.900 81.010 246.160 81.690 ;
        RECT 246.330 81.080 246.580 81.860 ;
        RECT 246.830 81.310 247.080 81.690 ;
        RECT 247.250 81.480 247.605 81.860 ;
        RECT 248.610 81.470 248.945 81.690 ;
        RECT 248.210 81.310 248.440 81.350 ;
        RECT 246.830 81.110 248.440 81.310 ;
        RECT 246.830 81.100 247.665 81.110 ;
        RECT 248.255 81.020 248.440 81.110 ;
        RECT 242.580 80.130 242.750 80.680 ;
        RECT 242.980 80.300 243.345 80.500 ;
        RECT 243.515 80.300 243.845 80.500 ;
        RECT 242.580 79.960 243.380 80.130 ;
        RECT 242.240 79.820 242.425 79.890 ;
        RECT 242.240 79.810 242.450 79.820 ;
        RECT 242.240 79.480 242.495 79.810 ;
        RECT 242.710 79.310 243.040 79.790 ;
        RECT 243.210 79.730 243.380 79.960 ;
        RECT 243.560 79.900 243.845 80.300 ;
        RECT 244.115 80.300 244.590 80.500 ;
        RECT 244.760 80.300 245.205 80.500 ;
        RECT 245.375 80.300 245.725 80.510 ;
        RECT 244.115 79.900 244.395 80.300 ;
        RECT 244.575 79.960 245.640 80.130 ;
        RECT 244.575 79.730 244.745 79.960 ;
        RECT 243.210 79.480 244.745 79.730 ;
        RECT 244.970 79.310 245.300 79.790 ;
        RECT 245.470 79.480 245.640 79.960 ;
        RECT 245.900 79.820 246.070 81.010 ;
        RECT 247.770 80.910 248.100 80.940 ;
        RECT 246.300 80.850 248.100 80.910 ;
        RECT 248.690 80.850 248.945 81.470 ;
        RECT 246.240 80.740 248.945 80.850 ;
        RECT 246.240 80.705 246.440 80.740 ;
        RECT 246.240 80.130 246.410 80.705 ;
        RECT 247.770 80.680 248.945 80.740 ;
        RECT 249.120 81.140 249.580 81.690 ;
        RECT 249.770 81.140 250.100 81.860 ;
        RECT 246.640 80.265 247.050 80.570 ;
        RECT 247.220 80.300 247.550 80.510 ;
        RECT 246.240 80.010 246.510 80.130 ;
        RECT 246.240 79.965 247.085 80.010 ;
        RECT 246.330 79.840 247.085 79.965 ;
        RECT 247.340 79.900 247.550 80.300 ;
        RECT 247.795 80.300 248.270 80.510 ;
        RECT 248.460 80.300 248.950 80.500 ;
        RECT 247.795 79.900 248.015 80.300 ;
        RECT 245.900 79.810 246.130 79.820 ;
        RECT 245.900 79.480 246.160 79.810 ;
        RECT 246.915 79.690 247.085 79.840 ;
        RECT 246.330 79.310 246.660 79.670 ;
        RECT 246.915 79.480 248.215 79.690 ;
        RECT 248.490 79.310 248.945 80.075 ;
        RECT 249.120 79.770 249.370 81.140 ;
        RECT 250.300 80.970 250.600 81.520 ;
        RECT 250.770 81.190 251.050 81.860 ;
        RECT 249.660 80.800 250.600 80.970 ;
        RECT 249.660 80.550 249.830 80.800 ;
        RECT 250.970 80.550 251.235 80.910 ;
        RECT 252.340 80.695 252.630 81.860 ;
        RECT 252.800 80.770 256.310 81.860 ;
        RECT 249.540 80.220 249.830 80.550 ;
        RECT 250.000 80.300 250.340 80.550 ;
        RECT 250.560 80.300 251.235 80.550 ;
        RECT 249.660 80.130 249.830 80.220 ;
        RECT 249.660 79.940 251.050 80.130 ;
        RECT 252.800 80.080 254.450 80.600 ;
        RECT 254.620 80.250 256.310 80.770 ;
        RECT 256.570 80.850 256.740 81.690 ;
        RECT 256.910 81.520 258.080 81.690 ;
        RECT 256.910 81.020 257.240 81.520 ;
        RECT 257.750 81.480 258.080 81.520 ;
        RECT 258.270 81.440 258.625 81.860 ;
        RECT 257.410 81.260 257.640 81.350 ;
        RECT 258.795 81.260 259.045 81.690 ;
        RECT 257.410 81.020 259.045 81.260 ;
        RECT 259.215 81.100 259.545 81.860 ;
        RECT 259.715 81.020 259.970 81.690 ;
        RECT 259.760 81.010 259.970 81.020 ;
        RECT 256.570 80.680 259.630 80.850 ;
        RECT 256.485 80.300 256.835 80.510 ;
        RECT 257.005 80.300 257.450 80.500 ;
        RECT 257.620 80.300 258.095 80.500 ;
        RECT 249.120 79.480 249.680 79.770 ;
        RECT 249.850 79.310 250.100 79.770 ;
        RECT 250.720 79.580 251.050 79.940 ;
        RECT 252.340 79.310 252.630 80.035 ;
        RECT 252.800 79.310 256.310 80.080 ;
        RECT 256.570 79.960 257.635 80.130 ;
        RECT 256.570 79.480 256.740 79.960 ;
        RECT 256.910 79.310 257.240 79.790 ;
        RECT 257.465 79.730 257.635 79.960 ;
        RECT 257.815 79.900 258.095 80.300 ;
        RECT 258.365 80.300 258.695 80.500 ;
        RECT 258.865 80.300 259.230 80.500 ;
        RECT 258.365 79.900 258.650 80.300 ;
        RECT 259.460 80.130 259.630 80.680 ;
        RECT 258.830 79.960 259.630 80.130 ;
        RECT 258.830 79.730 259.000 79.960 ;
        RECT 259.800 79.890 259.970 81.010 ;
        RECT 260.250 80.850 260.420 81.690 ;
        RECT 260.590 81.520 261.760 81.690 ;
        RECT 260.590 81.020 260.920 81.520 ;
        RECT 261.430 81.480 261.760 81.520 ;
        RECT 261.950 81.440 262.305 81.860 ;
        RECT 261.090 81.260 261.320 81.350 ;
        RECT 262.475 81.260 262.725 81.690 ;
        RECT 261.090 81.020 262.725 81.260 ;
        RECT 262.895 81.100 263.225 81.860 ;
        RECT 263.395 81.020 263.650 81.690 ;
        RECT 260.250 80.680 263.310 80.850 ;
        RECT 260.165 80.300 260.515 80.510 ;
        RECT 260.685 80.300 261.130 80.500 ;
        RECT 261.300 80.300 261.775 80.500 ;
        RECT 259.785 79.810 259.970 79.890 ;
        RECT 257.465 79.480 259.000 79.730 ;
        RECT 259.170 79.310 259.500 79.790 ;
        RECT 259.715 79.480 259.970 79.810 ;
        RECT 260.250 79.960 261.315 80.130 ;
        RECT 260.250 79.480 260.420 79.960 ;
        RECT 260.590 79.310 260.920 79.790 ;
        RECT 261.145 79.730 261.315 79.960 ;
        RECT 261.495 79.900 261.775 80.300 ;
        RECT 262.045 80.300 262.375 80.500 ;
        RECT 262.545 80.300 262.910 80.500 ;
        RECT 262.045 79.900 262.330 80.300 ;
        RECT 263.140 80.130 263.310 80.680 ;
        RECT 262.510 79.960 263.310 80.130 ;
        RECT 262.510 79.730 262.680 79.960 ;
        RECT 263.480 79.890 263.650 81.020 ;
        RECT 263.845 81.470 264.180 81.690 ;
        RECT 265.185 81.480 265.540 81.860 ;
        RECT 263.845 80.850 264.100 81.470 ;
        RECT 264.350 81.310 264.580 81.350 ;
        RECT 265.710 81.310 265.960 81.690 ;
        RECT 264.350 81.110 265.960 81.310 ;
        RECT 264.350 81.020 264.535 81.110 ;
        RECT 265.125 81.100 265.960 81.110 ;
        RECT 266.210 81.080 266.460 81.860 ;
        RECT 266.630 81.010 266.890 81.690 ;
        RECT 267.065 81.350 268.720 81.640 ;
        RECT 264.690 80.910 265.020 80.940 ;
        RECT 264.690 80.850 266.490 80.910 ;
        RECT 263.845 80.740 266.550 80.850 ;
        RECT 263.845 80.680 265.020 80.740 ;
        RECT 266.350 80.705 266.550 80.740 ;
        RECT 263.840 80.300 264.330 80.500 ;
        RECT 264.520 80.300 264.995 80.510 ;
        RECT 263.465 79.810 263.650 79.890 ;
        RECT 261.145 79.480 262.680 79.730 ;
        RECT 262.850 79.310 263.180 79.790 ;
        RECT 263.395 79.480 263.650 79.810 ;
        RECT 263.845 79.310 264.300 80.075 ;
        RECT 264.775 79.900 264.995 80.300 ;
        RECT 265.240 80.300 265.570 80.510 ;
        RECT 265.240 79.900 265.450 80.300 ;
        RECT 265.740 80.265 266.150 80.570 ;
        RECT 266.380 80.130 266.550 80.705 ;
        RECT 266.280 80.010 266.550 80.130 ;
        RECT 265.705 79.965 266.550 80.010 ;
        RECT 265.705 79.840 266.460 79.965 ;
        RECT 265.705 79.690 265.875 79.840 ;
        RECT 266.720 79.810 266.890 81.010 ;
        RECT 267.065 81.010 268.655 81.180 ;
        RECT 268.890 81.060 269.170 81.860 ;
        RECT 267.065 80.720 267.385 81.010 ;
        RECT 268.485 80.890 268.655 81.010 ;
        RECT 267.580 80.670 268.295 80.840 ;
        RECT 268.485 80.720 269.210 80.890 ;
        RECT 269.380 80.720 269.650 81.690 ;
        RECT 269.820 81.425 275.165 81.860 ;
        RECT 267.065 79.980 267.415 80.550 ;
        RECT 267.585 80.220 268.295 80.670 ;
        RECT 269.040 80.550 269.210 80.720 ;
        RECT 268.465 80.220 268.870 80.550 ;
        RECT 269.040 80.220 269.310 80.550 ;
        RECT 269.040 80.050 269.210 80.220 ;
        RECT 267.600 79.880 269.210 80.050 ;
        RECT 269.480 79.985 269.650 80.720 ;
        RECT 264.575 79.480 265.875 79.690 ;
        RECT 266.130 79.310 266.460 79.670 ;
        RECT 266.630 79.480 266.890 79.810 ;
        RECT 267.070 79.310 267.400 79.810 ;
        RECT 267.600 79.530 267.770 79.880 ;
        RECT 267.970 79.310 268.300 79.710 ;
        RECT 268.470 79.530 268.640 79.880 ;
        RECT 268.810 79.310 269.190 79.710 ;
        RECT 269.380 79.640 269.650 79.985 ;
        RECT 271.405 79.855 271.745 80.685 ;
        RECT 273.225 80.175 273.575 81.425 ;
        RECT 275.540 81.190 275.820 81.860 ;
        RECT 275.340 80.550 275.655 80.990 ;
        RECT 275.990 80.970 276.290 81.520 ;
        RECT 276.500 81.140 276.830 81.860 ;
        RECT 277.020 81.140 277.470 81.690 ;
        RECT 275.990 80.800 276.930 80.970 ;
        RECT 276.760 80.550 276.930 80.800 ;
        RECT 275.340 80.300 276.030 80.550 ;
        RECT 276.260 80.300 276.590 80.550 ;
        RECT 276.760 80.220 277.050 80.550 ;
        RECT 276.760 80.130 276.930 80.220 ;
        RECT 275.540 79.940 276.930 80.130 ;
        RECT 269.820 79.310 275.165 79.855 ;
        RECT 275.540 79.580 275.870 79.940 ;
        RECT 277.220 79.770 277.470 81.140 ;
        RECT 277.640 80.720 277.930 81.860 ;
        RECT 278.100 80.695 278.390 81.860 ;
        RECT 278.560 80.770 280.230 81.860 ;
        RECT 276.500 79.310 276.750 79.770 ;
        RECT 276.920 79.480 277.470 79.770 ;
        RECT 277.640 79.310 277.930 80.110 ;
        RECT 278.560 80.080 279.310 80.600 ;
        RECT 279.480 80.250 280.230 80.770 ;
        RECT 280.405 80.720 280.740 81.690 ;
        RECT 280.910 80.720 281.080 81.860 ;
        RECT 281.250 81.520 283.280 81.690 ;
        RECT 278.100 79.310 278.390 80.035 ;
        RECT 278.560 79.310 280.230 80.080 ;
        RECT 280.405 80.050 280.575 80.720 ;
        RECT 281.250 80.550 281.420 81.520 ;
        RECT 280.745 80.220 281.000 80.550 ;
        RECT 281.225 80.220 281.420 80.550 ;
        RECT 281.590 81.180 282.715 81.350 ;
        RECT 280.830 80.050 281.000 80.220 ;
        RECT 281.590 80.050 281.760 81.180 ;
        RECT 280.405 79.480 280.660 80.050 ;
        RECT 280.830 79.880 281.760 80.050 ;
        RECT 281.930 80.840 282.940 81.010 ;
        RECT 281.930 80.040 282.100 80.840 ;
        RECT 282.305 80.160 282.580 80.640 ;
        RECT 282.300 79.990 282.580 80.160 ;
        RECT 281.585 79.845 281.760 79.880 ;
        RECT 280.830 79.310 281.160 79.710 ;
        RECT 281.585 79.480 282.115 79.845 ;
        RECT 282.305 79.480 282.580 79.990 ;
        RECT 282.750 79.480 282.940 80.840 ;
        RECT 283.110 80.855 283.280 81.520 ;
        RECT 283.450 81.100 283.620 81.860 ;
        RECT 283.855 81.100 284.370 81.510 ;
        RECT 283.110 80.665 283.860 80.855 ;
        RECT 284.030 80.290 284.370 81.100 ;
        RECT 284.540 80.770 287.130 81.860 ;
        RECT 283.140 80.120 284.370 80.290 ;
        RECT 283.120 79.310 283.630 79.845 ;
        RECT 283.850 79.515 284.095 80.120 ;
        RECT 284.540 80.080 285.750 80.600 ;
        RECT 285.920 80.250 287.130 80.770 ;
        RECT 287.770 80.750 288.065 81.860 ;
        RECT 288.245 80.550 288.495 81.685 ;
        RECT 288.665 80.750 288.925 81.860 ;
        RECT 289.095 80.960 289.355 81.685 ;
        RECT 289.525 81.130 289.785 81.860 ;
        RECT 289.955 80.960 290.215 81.685 ;
        RECT 290.385 81.130 290.645 81.860 ;
        RECT 290.815 80.960 291.075 81.685 ;
        RECT 291.245 81.130 291.505 81.860 ;
        RECT 291.675 80.960 291.935 81.685 ;
        RECT 292.105 81.130 292.400 81.860 ;
        RECT 289.095 80.720 292.405 80.960 ;
        RECT 292.820 80.770 294.030 81.860 ;
        RECT 294.205 81.190 294.460 81.690 ;
        RECT 294.630 81.360 294.960 81.860 ;
        RECT 294.205 81.020 294.955 81.190 ;
        RECT 284.540 79.310 287.130 80.080 ;
        RECT 287.760 79.940 288.075 80.550 ;
        RECT 288.245 80.300 291.265 80.550 ;
        RECT 287.820 79.310 288.065 79.770 ;
        RECT 288.245 79.490 288.495 80.300 ;
        RECT 291.435 80.130 292.405 80.720 ;
        RECT 289.095 79.960 292.405 80.130 ;
        RECT 292.820 80.060 293.340 80.600 ;
        RECT 293.510 80.230 294.030 80.770 ;
        RECT 294.205 80.200 294.555 80.850 ;
        RECT 288.665 79.310 288.925 79.835 ;
        RECT 289.095 79.505 289.355 79.960 ;
        RECT 289.525 79.310 289.785 79.790 ;
        RECT 289.955 79.505 290.215 79.960 ;
        RECT 290.385 79.310 290.645 79.790 ;
        RECT 290.815 79.505 291.075 79.960 ;
        RECT 291.245 79.310 291.505 79.790 ;
        RECT 291.675 79.505 291.935 79.960 ;
        RECT 292.105 79.310 292.405 79.790 ;
        RECT 292.820 79.310 294.030 80.060 ;
        RECT 294.725 80.030 294.955 81.020 ;
        RECT 294.205 79.860 294.955 80.030 ;
        RECT 294.205 79.570 294.460 79.860 ;
        RECT 294.630 79.310 294.960 79.690 ;
        RECT 295.130 79.570 295.300 81.690 ;
        RECT 295.470 80.890 295.795 81.675 ;
        RECT 295.965 81.400 296.215 81.860 ;
        RECT 296.385 81.360 296.635 81.690 ;
        RECT 296.850 81.360 297.530 81.690 ;
        RECT 296.385 81.230 296.555 81.360 ;
        RECT 296.160 81.060 296.555 81.230 ;
        RECT 295.530 79.840 295.990 80.890 ;
        RECT 296.160 79.700 296.330 81.060 ;
        RECT 296.725 80.800 297.190 81.190 ;
        RECT 296.500 79.990 296.850 80.610 ;
        RECT 297.020 80.210 297.190 80.800 ;
        RECT 297.360 80.580 297.530 81.360 ;
        RECT 297.700 81.260 297.870 81.600 ;
        RECT 298.105 81.430 298.435 81.860 ;
        RECT 298.605 81.260 298.775 81.600 ;
        RECT 299.070 81.400 299.440 81.860 ;
        RECT 297.700 81.090 298.775 81.260 ;
        RECT 299.610 81.230 299.780 81.690 ;
        RECT 300.015 81.350 300.885 81.690 ;
        RECT 301.055 81.400 301.305 81.860 ;
        RECT 299.220 81.060 299.780 81.230 ;
        RECT 299.220 80.920 299.390 81.060 ;
        RECT 297.890 80.750 299.390 80.920 ;
        RECT 300.085 80.890 300.545 81.180 ;
        RECT 297.360 80.410 299.050 80.580 ;
        RECT 297.020 79.990 297.375 80.210 ;
        RECT 297.545 79.700 297.715 80.410 ;
        RECT 297.920 79.990 298.710 80.240 ;
        RECT 298.880 80.230 299.050 80.410 ;
        RECT 299.220 80.060 299.390 80.750 ;
        RECT 295.660 79.310 295.990 79.670 ;
        RECT 296.160 79.530 296.655 79.700 ;
        RECT 296.860 79.530 297.715 79.700 ;
        RECT 298.590 79.310 298.920 79.770 ;
        RECT 299.130 79.670 299.390 80.060 ;
        RECT 299.580 80.880 300.545 80.890 ;
        RECT 300.715 80.970 300.885 81.350 ;
        RECT 301.475 81.310 301.645 81.600 ;
        RECT 301.825 81.480 302.155 81.860 ;
        RECT 301.475 81.140 302.275 81.310 ;
        RECT 299.580 80.720 300.255 80.880 ;
        RECT 300.715 80.800 301.935 80.970 ;
        RECT 299.580 79.930 299.790 80.720 ;
        RECT 300.715 80.710 300.885 80.800 ;
        RECT 299.960 79.930 300.310 80.550 ;
        RECT 300.480 80.540 300.885 80.710 ;
        RECT 300.480 79.760 300.650 80.540 ;
        RECT 300.820 80.090 301.040 80.370 ;
        RECT 301.220 80.260 301.760 80.630 ;
        RECT 302.105 80.550 302.275 81.140 ;
        RECT 302.495 80.720 302.800 81.860 ;
        RECT 302.970 80.670 303.225 81.550 ;
        RECT 303.860 80.695 304.150 81.860 ;
        RECT 304.320 81.425 309.665 81.860 ;
        RECT 302.105 80.520 302.845 80.550 ;
        RECT 300.820 79.920 301.350 80.090 ;
        RECT 299.130 79.500 299.480 79.670 ;
        RECT 299.700 79.480 300.650 79.760 ;
        RECT 300.820 79.310 301.010 79.750 ;
        RECT 301.180 79.690 301.350 79.920 ;
        RECT 301.520 79.860 301.760 80.260 ;
        RECT 301.930 80.220 302.845 80.520 ;
        RECT 301.930 80.045 302.255 80.220 ;
        RECT 301.930 79.690 302.250 80.045 ;
        RECT 303.015 80.020 303.225 80.670 ;
        RECT 301.180 79.520 302.250 79.690 ;
        RECT 302.495 79.310 302.800 79.770 ;
        RECT 302.970 79.490 303.225 80.020 ;
        RECT 303.860 79.310 304.150 80.035 ;
        RECT 305.905 79.855 306.245 80.685 ;
        RECT 307.725 80.175 308.075 81.425 ;
        RECT 309.840 80.770 311.050 81.860 ;
        RECT 309.840 80.230 310.360 80.770 ;
        RECT 310.530 80.060 311.050 80.600 ;
        RECT 304.320 79.310 309.665 79.855 ;
        RECT 309.840 79.310 311.050 80.060 ;
        RECT 162.095 79.140 311.135 79.310 ;
        RECT 162.180 78.390 163.390 79.140 ;
        RECT 163.560 78.595 168.905 79.140 ;
        RECT 162.180 77.850 162.700 78.390 ;
        RECT 162.870 77.680 163.390 78.220 ;
        RECT 165.145 77.765 165.485 78.595 ;
        RECT 169.080 78.370 172.590 79.140 ;
        RECT 172.765 78.400 173.020 78.970 ;
        RECT 173.190 78.740 173.520 79.140 ;
        RECT 173.945 78.605 174.475 78.970 ;
        RECT 173.945 78.570 174.120 78.605 ;
        RECT 173.190 78.400 174.120 78.570 ;
        RECT 162.180 76.590 163.390 77.680 ;
        RECT 166.965 77.025 167.315 78.275 ;
        RECT 169.080 77.850 170.730 78.370 ;
        RECT 170.900 77.680 172.590 78.200 ;
        RECT 163.560 76.590 168.905 77.025 ;
        RECT 169.080 76.590 172.590 77.680 ;
        RECT 172.765 77.730 172.935 78.400 ;
        RECT 173.190 78.230 173.360 78.400 ;
        RECT 173.105 77.900 173.360 78.230 ;
        RECT 173.585 77.900 173.780 78.230 ;
        RECT 172.765 76.760 173.100 77.730 ;
        RECT 173.270 76.590 173.440 77.730 ;
        RECT 173.610 76.930 173.780 77.900 ;
        RECT 173.950 77.270 174.120 78.400 ;
        RECT 174.290 77.610 174.460 78.410 ;
        RECT 174.665 78.120 174.940 78.970 ;
        RECT 174.660 77.950 174.940 78.120 ;
        RECT 174.665 77.810 174.940 77.950 ;
        RECT 175.110 77.610 175.300 78.970 ;
        RECT 175.480 78.605 175.990 79.140 ;
        RECT 176.210 78.330 176.455 78.935 ;
        RECT 176.905 78.590 177.160 78.880 ;
        RECT 177.330 78.760 177.660 79.140 ;
        RECT 176.905 78.420 177.655 78.590 ;
        RECT 175.500 78.160 176.730 78.330 ;
        RECT 174.290 77.440 175.300 77.610 ;
        RECT 175.470 77.595 176.220 77.785 ;
        RECT 173.950 77.100 175.075 77.270 ;
        RECT 175.470 76.930 175.640 77.595 ;
        RECT 176.390 77.350 176.730 78.160 ;
        RECT 176.905 77.600 177.255 78.250 ;
        RECT 177.425 77.430 177.655 78.420 ;
        RECT 173.610 76.760 175.640 76.930 ;
        RECT 175.810 76.590 175.980 77.350 ;
        RECT 176.215 76.940 176.730 77.350 ;
        RECT 176.905 77.260 177.655 77.430 ;
        RECT 176.905 76.760 177.160 77.260 ;
        RECT 177.330 76.590 177.660 77.090 ;
        RECT 177.830 76.760 178.000 78.880 ;
        RECT 178.360 78.780 178.690 79.140 ;
        RECT 178.860 78.750 179.355 78.920 ;
        RECT 179.560 78.750 180.415 78.920 ;
        RECT 178.230 77.560 178.690 78.610 ;
        RECT 178.170 76.775 178.495 77.560 ;
        RECT 178.860 77.390 179.030 78.750 ;
        RECT 179.200 77.840 179.550 78.460 ;
        RECT 179.720 78.240 180.075 78.460 ;
        RECT 179.720 77.650 179.890 78.240 ;
        RECT 180.245 78.040 180.415 78.750 ;
        RECT 181.290 78.680 181.620 79.140 ;
        RECT 181.830 78.780 182.180 78.950 ;
        RECT 180.620 78.210 181.410 78.460 ;
        RECT 181.830 78.390 182.090 78.780 ;
        RECT 182.400 78.690 183.350 78.970 ;
        RECT 183.520 78.700 183.710 79.140 ;
        RECT 183.880 78.760 184.950 78.930 ;
        RECT 181.580 78.040 181.750 78.220 ;
        RECT 178.860 77.220 179.255 77.390 ;
        RECT 179.425 77.260 179.890 77.650 ;
        RECT 180.060 77.870 181.750 78.040 ;
        RECT 179.085 77.090 179.255 77.220 ;
        RECT 180.060 77.090 180.230 77.870 ;
        RECT 181.920 77.700 182.090 78.390 ;
        RECT 180.590 77.530 182.090 77.700 ;
        RECT 182.280 77.730 182.490 78.520 ;
        RECT 182.660 77.900 183.010 78.520 ;
        RECT 183.180 77.910 183.350 78.690 ;
        RECT 183.880 78.530 184.050 78.760 ;
        RECT 183.520 78.360 184.050 78.530 ;
        RECT 183.520 78.080 183.740 78.360 ;
        RECT 184.220 78.190 184.460 78.590 ;
        RECT 183.180 77.740 183.585 77.910 ;
        RECT 183.920 77.820 184.460 78.190 ;
        RECT 184.630 78.405 184.950 78.760 ;
        RECT 185.195 78.680 185.500 79.140 ;
        RECT 185.670 78.430 185.920 78.960 ;
        RECT 184.630 78.230 184.955 78.405 ;
        RECT 184.630 77.930 185.545 78.230 ;
        RECT 184.805 77.900 185.545 77.930 ;
        RECT 182.280 77.570 182.955 77.730 ;
        RECT 183.415 77.650 183.585 77.740 ;
        RECT 182.280 77.560 183.245 77.570 ;
        RECT 181.920 77.390 182.090 77.530 ;
        RECT 178.665 76.590 178.915 77.050 ;
        RECT 179.085 76.760 179.335 77.090 ;
        RECT 179.550 76.760 180.230 77.090 ;
        RECT 180.400 77.190 181.475 77.360 ;
        RECT 181.920 77.220 182.480 77.390 ;
        RECT 182.785 77.270 183.245 77.560 ;
        RECT 183.415 77.480 184.635 77.650 ;
        RECT 180.400 76.850 180.570 77.190 ;
        RECT 180.805 76.590 181.135 77.020 ;
        RECT 181.305 76.850 181.475 77.190 ;
        RECT 181.770 76.590 182.140 77.050 ;
        RECT 182.310 76.760 182.480 77.220 ;
        RECT 183.415 77.100 183.585 77.480 ;
        RECT 184.805 77.310 184.975 77.900 ;
        RECT 185.715 77.780 185.920 78.430 ;
        RECT 186.090 78.385 186.340 79.140 ;
        RECT 186.560 78.390 187.770 79.140 ;
        RECT 187.940 78.415 188.230 79.140 ;
        RECT 188.410 78.650 188.740 79.140 ;
        RECT 188.910 78.545 189.530 78.970 ;
        RECT 186.560 77.850 187.080 78.390 ;
        RECT 182.715 76.760 183.585 77.100 ;
        RECT 184.175 77.140 184.975 77.310 ;
        RECT 183.755 76.590 184.005 77.050 ;
        RECT 184.175 76.850 184.345 77.140 ;
        RECT 184.525 76.590 184.855 76.970 ;
        RECT 185.195 76.590 185.500 77.730 ;
        RECT 185.670 76.900 185.920 77.780 ;
        RECT 186.090 76.590 186.340 77.730 ;
        RECT 187.250 77.680 187.770 78.220 ;
        RECT 188.400 77.900 188.740 78.480 ;
        RECT 188.910 78.210 189.270 78.545 ;
        RECT 189.990 78.450 190.320 79.140 ;
        RECT 192.095 78.615 192.390 79.140 ;
        RECT 192.560 78.500 192.785 78.945 ;
        RECT 192.955 78.670 193.285 79.140 ;
        RECT 193.705 78.660 194.005 79.140 ;
        RECT 192.560 78.330 193.290 78.500 ;
        RECT 194.175 78.490 194.435 78.945 ;
        RECT 194.605 78.660 194.865 79.140 ;
        RECT 195.035 78.490 195.295 78.945 ;
        RECT 195.465 78.660 195.725 79.140 ;
        RECT 195.895 78.490 196.155 78.945 ;
        RECT 196.325 78.660 196.585 79.140 ;
        RECT 196.755 78.490 197.015 78.945 ;
        RECT 197.185 78.615 197.445 79.140 ;
        RECT 188.910 77.930 190.330 78.210 ;
        RECT 191.620 77.935 192.840 78.160 ;
        RECT 186.560 76.590 187.770 77.680 ;
        RECT 187.940 76.590 188.230 77.755 ;
        RECT 188.410 76.590 188.740 77.730 ;
        RECT 188.910 76.760 189.270 77.930 ;
        RECT 189.470 76.590 189.800 77.760 ;
        RECT 190.000 76.760 190.330 77.930 ;
        RECT 193.010 77.765 193.290 78.330 ;
        RECT 190.530 76.590 190.860 77.760 ;
        RECT 191.690 77.595 193.290 77.765 ;
        RECT 193.705 78.320 197.015 78.490 ;
        RECT 193.705 77.730 194.675 78.320 ;
        RECT 197.615 78.150 197.865 78.960 ;
        RECT 198.045 78.680 198.290 79.140 ;
        RECT 194.845 77.900 197.865 78.150 ;
        RECT 198.035 77.900 198.350 78.510 ;
        RECT 198.725 78.360 199.225 78.970 ;
        RECT 198.520 77.900 198.870 78.150 ;
        RECT 191.690 76.790 191.945 77.595 ;
        RECT 192.115 76.590 192.375 77.425 ;
        RECT 192.545 76.790 192.805 77.595 ;
        RECT 193.705 77.490 197.015 77.730 ;
        RECT 192.975 76.590 193.230 77.425 ;
        RECT 193.710 76.590 194.005 77.320 ;
        RECT 194.175 76.765 194.435 77.490 ;
        RECT 194.605 76.590 194.865 77.320 ;
        RECT 195.035 76.765 195.295 77.490 ;
        RECT 195.465 76.590 195.725 77.320 ;
        RECT 195.895 76.765 196.155 77.490 ;
        RECT 196.325 76.590 196.585 77.320 ;
        RECT 196.755 76.765 197.015 77.490 ;
        RECT 197.185 76.590 197.445 77.700 ;
        RECT 197.615 76.765 197.865 77.900 ;
        RECT 199.055 77.730 199.225 78.360 ;
        RECT 199.855 78.490 200.185 78.970 ;
        RECT 200.355 78.680 200.580 79.140 ;
        RECT 200.750 78.490 201.080 78.970 ;
        RECT 199.855 78.320 201.080 78.490 ;
        RECT 201.270 78.340 201.520 79.140 ;
        RECT 201.690 78.340 202.030 78.970 ;
        RECT 203.120 78.650 203.390 79.140 ;
        RECT 199.395 77.950 199.725 78.150 ;
        RECT 199.895 77.950 200.225 78.150 ;
        RECT 200.395 77.950 200.815 78.150 ;
        RECT 200.990 77.980 201.685 78.150 ;
        RECT 200.990 77.730 201.160 77.980 ;
        RECT 201.855 77.730 202.030 78.340 ;
        RECT 203.180 77.900 203.445 78.480 ;
        RECT 203.615 78.210 203.890 78.920 ;
        RECT 204.090 78.655 204.875 78.920 ;
        RECT 203.615 77.980 204.450 78.210 ;
        RECT 198.045 76.590 198.340 77.700 ;
        RECT 198.725 77.560 201.160 77.730 ;
        RECT 198.725 76.760 199.055 77.560 ;
        RECT 199.225 76.590 199.555 77.390 ;
        RECT 199.855 76.760 200.185 77.560 ;
        RECT 200.830 76.590 201.080 77.390 ;
        RECT 201.350 76.590 201.520 77.730 ;
        RECT 201.690 76.760 202.030 77.730 ;
        RECT 203.120 76.590 203.435 77.650 ;
        RECT 203.615 77.320 203.890 77.980 ;
        RECT 204.620 77.800 204.875 78.655 ;
        RECT 205.045 78.460 205.255 78.920 ;
        RECT 205.445 78.645 205.775 79.140 ;
        RECT 205.950 78.510 206.195 78.970 ;
        RECT 205.045 77.980 205.455 78.460 ;
        RECT 206.025 78.300 206.195 78.510 ;
        RECT 206.365 78.480 206.630 79.140 ;
        RECT 206.860 78.680 207.105 79.140 ;
        RECT 205.625 77.800 205.855 78.230 ;
        RECT 204.085 77.630 205.855 77.800 ;
        RECT 206.025 77.780 206.630 78.300 ;
        RECT 206.800 77.900 207.115 78.510 ;
        RECT 207.285 78.150 207.535 78.960 ;
        RECT 207.705 78.615 207.965 79.140 ;
        RECT 208.135 78.490 208.395 78.945 ;
        RECT 208.565 78.660 208.825 79.140 ;
        RECT 208.995 78.490 209.255 78.945 ;
        RECT 209.425 78.660 209.685 79.140 ;
        RECT 209.855 78.490 210.115 78.945 ;
        RECT 210.285 78.660 210.545 79.140 ;
        RECT 210.715 78.490 210.975 78.945 ;
        RECT 211.145 78.660 211.445 79.140 ;
        RECT 208.135 78.320 211.445 78.490 ;
        RECT 207.285 77.900 210.305 78.150 ;
        RECT 204.085 77.265 204.320 77.630 ;
        RECT 204.490 77.270 204.820 77.460 ;
        RECT 205.045 77.335 205.235 77.630 ;
        RECT 206.025 77.440 206.195 77.780 ;
        RECT 204.490 77.095 204.680 77.270 ;
        RECT 204.065 76.590 204.680 77.095 ;
        RECT 204.850 76.760 205.325 77.100 ;
        RECT 205.495 76.590 205.710 77.435 ;
        RECT 205.940 77.430 206.195 77.440 ;
        RECT 205.910 76.760 206.195 77.430 ;
        RECT 206.365 76.590 206.630 77.600 ;
        RECT 206.810 76.590 207.105 77.700 ;
        RECT 207.285 76.765 207.535 77.900 ;
        RECT 210.475 77.730 211.445 78.320 ;
        RECT 211.860 78.370 213.530 79.140 ;
        RECT 213.700 78.415 213.990 79.140 ;
        RECT 215.085 78.400 215.340 78.970 ;
        RECT 215.510 78.740 215.840 79.140 ;
        RECT 216.265 78.605 216.795 78.970 ;
        RECT 216.265 78.570 216.440 78.605 ;
        RECT 215.510 78.400 216.440 78.570 ;
        RECT 216.985 78.460 217.260 78.970 ;
        RECT 211.860 77.850 212.610 78.370 ;
        RECT 207.705 76.590 207.965 77.700 ;
        RECT 208.135 77.490 211.445 77.730 ;
        RECT 212.780 77.680 213.530 78.200 ;
        RECT 208.135 76.765 208.395 77.490 ;
        RECT 208.565 76.590 208.825 77.320 ;
        RECT 208.995 76.765 209.255 77.490 ;
        RECT 209.425 76.590 209.685 77.320 ;
        RECT 209.855 76.765 210.115 77.490 ;
        RECT 210.285 76.590 210.545 77.320 ;
        RECT 210.715 76.765 210.975 77.490 ;
        RECT 211.145 76.590 211.440 77.320 ;
        RECT 211.860 76.590 213.530 77.680 ;
        RECT 213.700 76.590 213.990 77.755 ;
        RECT 215.085 77.730 215.255 78.400 ;
        RECT 215.510 78.230 215.680 78.400 ;
        RECT 215.425 77.900 215.680 78.230 ;
        RECT 215.905 77.900 216.100 78.230 ;
        RECT 215.085 76.760 215.420 77.730 ;
        RECT 215.590 76.590 215.760 77.730 ;
        RECT 215.930 76.930 216.100 77.900 ;
        RECT 216.270 77.270 216.440 78.400 ;
        RECT 216.610 77.610 216.780 78.410 ;
        RECT 216.980 78.290 217.260 78.460 ;
        RECT 216.985 77.810 217.260 78.290 ;
        RECT 217.430 77.610 217.620 78.970 ;
        RECT 217.800 78.605 218.310 79.140 ;
        RECT 218.530 78.330 218.775 78.935 ;
        RECT 219.385 78.630 219.625 79.140 ;
        RECT 219.805 78.630 220.085 78.960 ;
        RECT 220.315 78.630 220.530 79.140 ;
        RECT 217.820 78.160 219.050 78.330 ;
        RECT 216.610 77.440 217.620 77.610 ;
        RECT 217.790 77.595 218.540 77.785 ;
        RECT 216.270 77.100 217.395 77.270 ;
        RECT 217.790 76.930 217.960 77.595 ;
        RECT 218.710 77.350 219.050 78.160 ;
        RECT 219.280 77.900 219.635 78.460 ;
        RECT 219.805 77.730 219.975 78.630 ;
        RECT 220.145 77.900 220.410 78.460 ;
        RECT 220.700 78.400 221.315 78.970 ;
        RECT 220.660 77.730 220.830 78.230 ;
        RECT 219.405 77.560 220.830 77.730 ;
        RECT 219.405 77.385 219.795 77.560 ;
        RECT 215.930 76.760 217.960 76.930 ;
        RECT 218.130 76.590 218.300 77.350 ;
        RECT 218.535 76.940 219.050 77.350 ;
        RECT 220.280 76.590 220.610 77.390 ;
        RECT 221.000 77.380 221.315 78.400 ;
        RECT 221.520 78.370 223.190 79.140 ;
        RECT 221.520 77.850 222.270 78.370 ;
        RECT 222.440 77.680 223.190 78.200 ;
        RECT 220.780 76.760 221.315 77.380 ;
        RECT 221.520 76.590 223.190 77.680 ;
        RECT 223.820 78.195 224.160 78.970 ;
        RECT 224.330 78.680 224.500 79.140 ;
        RECT 224.740 78.705 225.100 78.970 ;
        RECT 224.740 78.700 225.095 78.705 ;
        RECT 224.740 78.690 225.090 78.700 ;
        RECT 224.740 78.685 225.085 78.690 ;
        RECT 224.740 78.675 225.080 78.685 ;
        RECT 225.730 78.680 225.900 79.140 ;
        RECT 224.740 78.670 225.075 78.675 ;
        RECT 224.740 78.660 225.065 78.670 ;
        RECT 224.740 78.650 225.055 78.660 ;
        RECT 224.740 78.510 225.040 78.650 ;
        RECT 224.330 78.320 225.040 78.510 ;
        RECT 225.230 78.510 225.560 78.590 ;
        RECT 226.070 78.510 226.410 78.970 ;
        RECT 226.580 78.650 226.850 79.140 ;
        RECT 225.230 78.320 226.410 78.510 ;
        RECT 223.820 76.760 224.100 78.195 ;
        RECT 224.330 77.750 224.615 78.320 ;
        RECT 224.800 77.920 225.270 78.150 ;
        RECT 225.440 78.130 225.770 78.150 ;
        RECT 225.440 77.950 225.890 78.130 ;
        RECT 226.080 77.950 226.410 78.150 ;
        RECT 224.330 77.535 225.480 77.750 ;
        RECT 224.270 76.590 224.980 77.365 ;
        RECT 225.150 76.760 225.480 77.535 ;
        RECT 225.675 76.835 225.890 77.950 ;
        RECT 226.180 77.610 226.410 77.950 ;
        RECT 226.640 77.900 226.905 78.480 ;
        RECT 227.075 78.210 227.350 78.920 ;
        RECT 227.550 78.655 228.335 78.920 ;
        RECT 227.075 77.980 227.910 78.210 ;
        RECT 226.070 76.590 226.400 77.310 ;
        RECT 226.580 76.590 226.895 77.650 ;
        RECT 227.075 77.320 227.350 77.980 ;
        RECT 228.080 77.800 228.335 78.655 ;
        RECT 228.505 78.460 228.715 78.920 ;
        RECT 228.905 78.645 229.235 79.140 ;
        RECT 229.410 78.510 229.655 78.970 ;
        RECT 228.505 77.980 228.915 78.460 ;
        RECT 229.485 78.300 229.655 78.510 ;
        RECT 229.825 78.480 230.090 79.140 ;
        RECT 230.260 78.595 235.605 79.140 ;
        RECT 229.085 77.800 229.315 78.230 ;
        RECT 227.545 77.630 229.315 77.800 ;
        RECT 229.485 77.780 230.090 78.300 ;
        RECT 227.545 77.265 227.780 77.630 ;
        RECT 227.950 77.270 228.280 77.460 ;
        RECT 228.505 77.335 228.695 77.630 ;
        RECT 227.950 77.095 228.140 77.270 ;
        RECT 227.525 76.590 228.140 77.095 ;
        RECT 228.310 76.760 228.785 77.100 ;
        RECT 228.955 76.590 229.170 77.435 ;
        RECT 229.485 77.430 229.655 77.780 ;
        RECT 231.845 77.765 232.185 78.595 ;
        RECT 235.780 78.370 239.290 79.140 ;
        RECT 239.460 78.415 239.750 79.140 ;
        RECT 239.920 78.370 242.510 79.140 ;
        RECT 243.150 78.640 243.480 79.140 ;
        RECT 243.680 78.570 243.850 78.920 ;
        RECT 244.050 78.740 244.380 79.140 ;
        RECT 244.550 78.570 244.720 78.920 ;
        RECT 244.890 78.740 245.270 79.140 ;
        RECT 229.370 76.760 229.655 77.430 ;
        RECT 229.825 76.590 230.090 77.600 ;
        RECT 233.665 77.025 234.015 78.275 ;
        RECT 235.780 77.850 237.430 78.370 ;
        RECT 237.600 77.680 239.290 78.200 ;
        RECT 239.920 77.850 241.130 78.370 ;
        RECT 230.260 76.590 235.605 77.025 ;
        RECT 235.780 76.590 239.290 77.680 ;
        RECT 239.460 76.590 239.750 77.755 ;
        RECT 241.300 77.680 242.510 78.200 ;
        RECT 243.145 77.900 243.495 78.470 ;
        RECT 243.680 78.400 245.290 78.570 ;
        RECT 245.460 78.465 245.730 78.810 ;
        RECT 245.900 78.595 251.245 79.140 ;
        RECT 251.420 78.595 256.765 79.140 ;
        RECT 245.120 78.230 245.290 78.400 ;
        RECT 243.665 77.780 244.375 78.230 ;
        RECT 244.545 77.900 244.950 78.230 ;
        RECT 245.120 77.900 245.390 78.230 ;
        RECT 239.920 76.590 242.510 77.680 ;
        RECT 243.145 77.440 243.465 77.730 ;
        RECT 243.660 77.610 244.375 77.780 ;
        RECT 245.120 77.730 245.290 77.900 ;
        RECT 245.560 77.730 245.730 78.465 ;
        RECT 247.485 77.765 247.825 78.595 ;
        RECT 244.565 77.560 245.290 77.730 ;
        RECT 244.565 77.440 244.735 77.560 ;
        RECT 243.145 77.270 244.735 77.440 ;
        RECT 243.145 76.810 244.800 77.100 ;
        RECT 244.970 76.590 245.250 77.390 ;
        RECT 245.460 76.760 245.730 77.730 ;
        RECT 249.305 77.025 249.655 78.275 ;
        RECT 253.005 77.765 253.345 78.595 ;
        RECT 257.405 78.375 257.860 79.140 ;
        RECT 258.135 78.760 259.435 78.970 ;
        RECT 259.690 78.780 260.020 79.140 ;
        RECT 259.265 78.610 259.435 78.760 ;
        RECT 260.190 78.640 260.450 78.970 ;
        RECT 260.220 78.630 260.450 78.640 ;
        RECT 254.825 77.025 255.175 78.275 ;
        RECT 258.335 78.150 258.555 78.550 ;
        RECT 257.400 77.950 257.890 78.150 ;
        RECT 258.080 77.940 258.555 78.150 ;
        RECT 258.800 78.150 259.010 78.550 ;
        RECT 259.265 78.485 260.020 78.610 ;
        RECT 259.265 78.440 260.110 78.485 ;
        RECT 259.840 78.320 260.110 78.440 ;
        RECT 258.800 77.940 259.130 78.150 ;
        RECT 259.300 77.880 259.710 78.185 ;
        RECT 257.405 77.710 258.580 77.770 ;
        RECT 259.940 77.745 260.110 78.320 ;
        RECT 259.910 77.710 260.110 77.745 ;
        RECT 257.405 77.600 260.110 77.710 ;
        RECT 245.900 76.590 251.245 77.025 ;
        RECT 251.420 76.590 256.765 77.025 ;
        RECT 257.405 76.980 257.660 77.600 ;
        RECT 258.250 77.540 260.050 77.600 ;
        RECT 258.250 77.510 258.580 77.540 ;
        RECT 260.280 77.440 260.450 78.630 ;
        RECT 260.625 78.375 261.080 79.140 ;
        RECT 261.355 78.760 262.655 78.970 ;
        RECT 262.910 78.780 263.240 79.140 ;
        RECT 262.485 78.610 262.655 78.760 ;
        RECT 263.410 78.640 263.670 78.970 ;
        RECT 263.440 78.630 263.670 78.640 ;
        RECT 261.555 78.150 261.775 78.550 ;
        RECT 260.620 77.950 261.110 78.150 ;
        RECT 261.300 77.940 261.775 78.150 ;
        RECT 262.020 78.150 262.230 78.550 ;
        RECT 262.485 78.485 263.240 78.610 ;
        RECT 262.485 78.440 263.330 78.485 ;
        RECT 263.060 78.320 263.330 78.440 ;
        RECT 262.020 77.940 262.350 78.150 ;
        RECT 262.520 77.880 262.930 78.185 ;
        RECT 257.910 77.340 258.095 77.430 ;
        RECT 258.685 77.340 259.520 77.350 ;
        RECT 257.910 77.140 259.520 77.340 ;
        RECT 257.910 77.100 258.140 77.140 ;
        RECT 257.405 76.760 257.740 76.980 ;
        RECT 258.745 76.590 259.100 76.970 ;
        RECT 259.270 76.760 259.520 77.140 ;
        RECT 259.770 76.590 260.020 77.370 ;
        RECT 260.190 76.760 260.450 77.440 ;
        RECT 260.625 77.710 261.800 77.770 ;
        RECT 263.160 77.745 263.330 78.320 ;
        RECT 263.130 77.710 263.330 77.745 ;
        RECT 260.625 77.600 263.330 77.710 ;
        RECT 260.625 76.980 260.880 77.600 ;
        RECT 261.470 77.540 263.270 77.600 ;
        RECT 261.470 77.510 261.800 77.540 ;
        RECT 263.500 77.440 263.670 78.630 ;
        RECT 263.840 78.390 265.050 79.140 ;
        RECT 265.220 78.415 265.510 79.140 ;
        RECT 265.880 78.510 266.210 78.870 ;
        RECT 266.830 78.680 267.080 79.140 ;
        RECT 267.250 78.680 267.810 78.970 ;
        RECT 263.840 77.850 264.360 78.390 ;
        RECT 265.880 78.320 267.270 78.510 ;
        RECT 267.100 78.230 267.270 78.320 ;
        RECT 264.530 77.680 265.050 78.220 ;
        RECT 265.695 77.900 266.370 78.150 ;
        RECT 266.590 77.900 266.930 78.150 ;
        RECT 267.100 77.900 267.390 78.230 ;
        RECT 261.130 77.340 261.315 77.430 ;
        RECT 261.905 77.340 262.740 77.350 ;
        RECT 261.130 77.140 262.740 77.340 ;
        RECT 261.130 77.100 261.360 77.140 ;
        RECT 260.625 76.760 260.960 76.980 ;
        RECT 261.965 76.590 262.320 76.970 ;
        RECT 262.490 76.760 262.740 77.140 ;
        RECT 262.990 76.590 263.240 77.370 ;
        RECT 263.410 76.760 263.670 77.440 ;
        RECT 263.840 76.590 265.050 77.680 ;
        RECT 265.220 76.590 265.510 77.755 ;
        RECT 265.695 77.540 265.960 77.900 ;
        RECT 267.100 77.650 267.270 77.900 ;
        RECT 266.330 77.480 267.270 77.650 ;
        RECT 265.880 76.590 266.160 77.260 ;
        RECT 266.330 76.930 266.630 77.480 ;
        RECT 267.560 77.310 267.810 78.680 ;
        RECT 267.980 78.595 273.325 79.140 ;
        RECT 269.565 77.765 269.905 78.595 ;
        RECT 273.500 78.370 276.090 79.140 ;
        RECT 276.725 78.590 276.980 78.880 ;
        RECT 277.150 78.760 277.480 79.140 ;
        RECT 276.725 78.420 277.475 78.590 ;
        RECT 266.830 76.590 267.160 77.310 ;
        RECT 267.350 76.760 267.810 77.310 ;
        RECT 271.385 77.025 271.735 78.275 ;
        RECT 273.500 77.850 274.710 78.370 ;
        RECT 274.880 77.680 276.090 78.200 ;
        RECT 267.980 76.590 273.325 77.025 ;
        RECT 273.500 76.590 276.090 77.680 ;
        RECT 276.725 77.600 277.075 78.250 ;
        RECT 277.245 77.430 277.475 78.420 ;
        RECT 276.725 77.260 277.475 77.430 ;
        RECT 276.725 76.760 276.980 77.260 ;
        RECT 277.150 76.590 277.480 77.090 ;
        RECT 277.650 76.760 277.820 78.880 ;
        RECT 278.180 78.780 278.510 79.140 ;
        RECT 278.680 78.750 279.175 78.920 ;
        RECT 279.380 78.750 280.235 78.920 ;
        RECT 278.050 77.560 278.510 78.610 ;
        RECT 277.990 76.775 278.315 77.560 ;
        RECT 278.680 77.390 278.850 78.750 ;
        RECT 279.020 77.840 279.370 78.460 ;
        RECT 279.540 78.240 279.895 78.460 ;
        RECT 279.540 77.650 279.710 78.240 ;
        RECT 280.065 78.040 280.235 78.750 ;
        RECT 281.110 78.680 281.440 79.140 ;
        RECT 281.650 78.780 282.000 78.950 ;
        RECT 280.440 78.210 281.230 78.460 ;
        RECT 281.650 78.390 281.910 78.780 ;
        RECT 282.220 78.690 283.170 78.970 ;
        RECT 283.340 78.700 283.530 79.140 ;
        RECT 283.700 78.760 284.770 78.930 ;
        RECT 281.400 78.040 281.570 78.220 ;
        RECT 278.680 77.220 279.075 77.390 ;
        RECT 279.245 77.260 279.710 77.650 ;
        RECT 279.880 77.870 281.570 78.040 ;
        RECT 278.905 77.090 279.075 77.220 ;
        RECT 279.880 77.090 280.050 77.870 ;
        RECT 281.740 77.700 281.910 78.390 ;
        RECT 280.410 77.530 281.910 77.700 ;
        RECT 282.100 77.730 282.310 78.520 ;
        RECT 282.480 77.900 282.830 78.520 ;
        RECT 283.000 77.910 283.170 78.690 ;
        RECT 283.700 78.530 283.870 78.760 ;
        RECT 283.340 78.360 283.870 78.530 ;
        RECT 283.340 78.080 283.560 78.360 ;
        RECT 284.040 78.190 284.280 78.590 ;
        RECT 283.000 77.740 283.405 77.910 ;
        RECT 283.740 77.820 284.280 78.190 ;
        RECT 284.450 78.405 284.770 78.760 ;
        RECT 285.015 78.680 285.320 79.140 ;
        RECT 285.490 78.430 285.745 78.960 ;
        RECT 285.980 78.680 286.225 79.140 ;
        RECT 284.450 78.230 284.775 78.405 ;
        RECT 284.450 77.930 285.365 78.230 ;
        RECT 284.625 77.900 285.365 77.930 ;
        RECT 282.100 77.570 282.775 77.730 ;
        RECT 283.235 77.650 283.405 77.740 ;
        RECT 282.100 77.560 283.065 77.570 ;
        RECT 281.740 77.390 281.910 77.530 ;
        RECT 278.485 76.590 278.735 77.050 ;
        RECT 278.905 76.760 279.155 77.090 ;
        RECT 279.370 76.760 280.050 77.090 ;
        RECT 280.220 77.190 281.295 77.360 ;
        RECT 281.740 77.220 282.300 77.390 ;
        RECT 282.605 77.270 283.065 77.560 ;
        RECT 283.235 77.480 284.455 77.650 ;
        RECT 280.220 76.850 280.390 77.190 ;
        RECT 280.625 76.590 280.955 77.020 ;
        RECT 281.125 76.850 281.295 77.190 ;
        RECT 281.590 76.590 281.960 77.050 ;
        RECT 282.130 76.760 282.300 77.220 ;
        RECT 283.235 77.100 283.405 77.480 ;
        RECT 284.625 77.310 284.795 77.900 ;
        RECT 285.535 77.780 285.745 78.430 ;
        RECT 285.920 77.900 286.235 78.510 ;
        RECT 286.405 78.150 286.655 78.960 ;
        RECT 286.825 78.615 287.085 79.140 ;
        RECT 287.255 78.490 287.515 78.945 ;
        RECT 287.685 78.660 287.945 79.140 ;
        RECT 288.115 78.490 288.375 78.945 ;
        RECT 288.545 78.660 288.805 79.140 ;
        RECT 288.975 78.490 289.235 78.945 ;
        RECT 289.405 78.660 289.665 79.140 ;
        RECT 289.835 78.490 290.095 78.945 ;
        RECT 290.265 78.660 290.565 79.140 ;
        RECT 287.255 78.320 290.565 78.490 ;
        RECT 290.980 78.415 291.270 79.140 ;
        RECT 291.450 78.490 291.780 78.965 ;
        RECT 291.950 78.660 292.120 79.140 ;
        RECT 292.290 78.490 292.620 78.965 ;
        RECT 292.790 78.660 292.960 79.140 ;
        RECT 293.130 78.490 293.460 78.965 ;
        RECT 293.630 78.660 293.800 79.140 ;
        RECT 293.970 78.490 294.300 78.965 ;
        RECT 294.470 78.660 294.640 79.140 ;
        RECT 294.810 78.490 295.140 78.965 ;
        RECT 295.310 78.660 295.480 79.140 ;
        RECT 295.650 78.965 295.900 78.970 ;
        RECT 295.650 78.490 295.980 78.965 ;
        RECT 296.150 78.660 296.320 79.140 ;
        RECT 296.570 78.965 296.740 78.970 ;
        RECT 296.490 78.490 296.820 78.965 ;
        RECT 296.990 78.660 297.160 79.140 ;
        RECT 297.410 78.965 297.580 78.970 ;
        RECT 297.330 78.490 297.660 78.965 ;
        RECT 297.830 78.660 298.000 79.140 ;
        RECT 298.170 78.490 298.500 78.965 ;
        RECT 298.670 78.660 298.840 79.140 ;
        RECT 299.010 78.490 299.340 78.965 ;
        RECT 299.510 78.660 299.680 79.140 ;
        RECT 299.850 78.490 300.180 78.965 ;
        RECT 300.350 78.660 300.520 79.140 ;
        RECT 300.690 78.490 301.020 78.965 ;
        RECT 301.190 78.660 301.360 79.140 ;
        RECT 301.530 78.490 301.860 78.965 ;
        RECT 302.030 78.660 302.200 79.140 ;
        RECT 302.480 78.595 307.825 79.140 ;
        RECT 291.450 78.320 292.960 78.490 ;
        RECT 293.130 78.320 295.480 78.490 ;
        RECT 295.650 78.320 302.310 78.490 ;
        RECT 286.405 77.900 289.425 78.150 ;
        RECT 282.535 76.760 283.405 77.100 ;
        RECT 283.995 77.140 284.795 77.310 ;
        RECT 283.575 76.590 283.825 77.050 ;
        RECT 283.995 76.850 284.165 77.140 ;
        RECT 284.345 76.590 284.675 76.970 ;
        RECT 285.015 76.590 285.320 77.730 ;
        RECT 285.490 76.900 285.745 77.780 ;
        RECT 285.930 76.590 286.225 77.700 ;
        RECT 286.405 76.765 286.655 77.900 ;
        RECT 289.595 77.730 290.565 78.320 ;
        RECT 292.790 78.150 292.960 78.320 ;
        RECT 295.305 78.150 295.480 78.320 ;
        RECT 291.445 77.950 292.620 78.150 ;
        RECT 292.790 77.950 295.100 78.150 ;
        RECT 295.305 77.950 301.865 78.150 ;
        RECT 292.790 77.780 292.960 77.950 ;
        RECT 295.305 77.780 295.480 77.950 ;
        RECT 302.035 77.780 302.310 78.320 ;
        RECT 286.825 76.590 287.085 77.700 ;
        RECT 287.255 77.490 290.565 77.730 ;
        RECT 287.255 76.765 287.515 77.490 ;
        RECT 287.685 76.590 287.945 77.320 ;
        RECT 288.115 76.765 288.375 77.490 ;
        RECT 288.545 76.590 288.805 77.320 ;
        RECT 288.975 76.765 289.235 77.490 ;
        RECT 289.405 76.590 289.665 77.320 ;
        RECT 289.835 76.765 290.095 77.490 ;
        RECT 290.265 76.590 290.560 77.320 ;
        RECT 290.980 76.590 291.270 77.755 ;
        RECT 291.450 77.610 292.960 77.780 ;
        RECT 293.130 77.610 295.480 77.780 ;
        RECT 295.650 77.610 302.310 77.780 ;
        RECT 304.065 77.765 304.405 78.595 ;
        RECT 308.000 78.370 309.670 79.140 ;
        RECT 309.840 78.390 311.050 79.140 ;
        RECT 291.450 76.760 291.780 77.610 ;
        RECT 291.950 76.590 292.120 77.440 ;
        RECT 292.290 76.760 292.620 77.610 ;
        RECT 292.790 76.590 292.960 77.440 ;
        RECT 293.130 76.760 293.460 77.610 ;
        RECT 293.630 76.590 293.800 77.390 ;
        RECT 293.970 76.760 294.300 77.610 ;
        RECT 294.470 76.590 294.640 77.390 ;
        RECT 294.810 76.760 295.140 77.610 ;
        RECT 295.310 76.590 295.480 77.390 ;
        RECT 295.650 76.760 295.980 77.610 ;
        RECT 296.150 76.590 296.320 77.390 ;
        RECT 296.490 76.760 296.820 77.610 ;
        RECT 296.990 76.590 297.160 77.390 ;
        RECT 297.330 76.760 297.660 77.610 ;
        RECT 297.830 76.590 298.000 77.390 ;
        RECT 298.170 76.760 298.500 77.610 ;
        RECT 298.670 76.590 298.840 77.390 ;
        RECT 299.010 76.760 299.340 77.610 ;
        RECT 299.510 76.590 299.680 77.390 ;
        RECT 299.850 76.760 300.180 77.610 ;
        RECT 300.350 76.590 300.520 77.390 ;
        RECT 300.690 76.760 301.020 77.610 ;
        RECT 301.190 76.590 301.360 77.390 ;
        RECT 301.530 76.760 301.860 77.610 ;
        RECT 302.030 76.590 302.200 77.390 ;
        RECT 305.885 77.025 306.235 78.275 ;
        RECT 308.000 77.850 308.750 78.370 ;
        RECT 308.920 77.680 309.670 78.200 ;
        RECT 302.480 76.590 307.825 77.025 ;
        RECT 308.000 76.590 309.670 77.680 ;
        RECT 309.840 77.680 310.360 78.220 ;
        RECT 310.530 77.850 311.050 78.390 ;
        RECT 309.840 76.590 311.050 77.680 ;
        RECT 162.095 76.420 311.135 76.590 ;
        RECT 162.180 75.330 163.390 76.420 ;
        RECT 163.560 75.330 165.230 76.420 ;
        RECT 165.865 75.750 166.120 76.250 ;
        RECT 166.290 75.920 166.620 76.420 ;
        RECT 165.865 75.580 166.615 75.750 ;
        RECT 162.180 74.620 162.700 75.160 ;
        RECT 162.870 74.790 163.390 75.330 ;
        RECT 163.560 74.640 164.310 75.160 ;
        RECT 164.480 74.810 165.230 75.330 ;
        RECT 165.865 74.760 166.215 75.410 ;
        RECT 162.180 73.870 163.390 74.620 ;
        RECT 163.560 73.870 165.230 74.640 ;
        RECT 166.385 74.590 166.615 75.580 ;
        RECT 165.865 74.420 166.615 74.590 ;
        RECT 165.865 74.130 166.120 74.420 ;
        RECT 166.290 73.870 166.620 74.250 ;
        RECT 166.790 74.130 166.960 76.250 ;
        RECT 167.130 75.450 167.455 76.235 ;
        RECT 167.625 75.960 167.875 76.420 ;
        RECT 168.045 75.920 168.295 76.250 ;
        RECT 168.510 75.920 169.190 76.250 ;
        RECT 168.045 75.790 168.215 75.920 ;
        RECT 167.820 75.620 168.215 75.790 ;
        RECT 167.190 74.400 167.650 75.450 ;
        RECT 167.820 74.260 167.990 75.620 ;
        RECT 168.385 75.360 168.850 75.750 ;
        RECT 168.160 74.550 168.510 75.170 ;
        RECT 168.680 74.770 168.850 75.360 ;
        RECT 169.020 75.140 169.190 75.920 ;
        RECT 169.360 75.820 169.530 76.160 ;
        RECT 169.765 75.990 170.095 76.420 ;
        RECT 170.265 75.820 170.435 76.160 ;
        RECT 170.730 75.960 171.100 76.420 ;
        RECT 169.360 75.650 170.435 75.820 ;
        RECT 171.270 75.790 171.440 76.250 ;
        RECT 171.675 75.910 172.545 76.250 ;
        RECT 172.715 75.960 172.965 76.420 ;
        RECT 170.880 75.620 171.440 75.790 ;
        RECT 170.880 75.480 171.050 75.620 ;
        RECT 169.550 75.310 171.050 75.480 ;
        RECT 171.745 75.450 172.205 75.740 ;
        RECT 169.020 74.970 170.710 75.140 ;
        RECT 168.680 74.550 169.035 74.770 ;
        RECT 169.205 74.260 169.375 74.970 ;
        RECT 169.580 74.550 170.370 74.800 ;
        RECT 170.540 74.790 170.710 74.970 ;
        RECT 170.880 74.620 171.050 75.310 ;
        RECT 167.320 73.870 167.650 74.230 ;
        RECT 167.820 74.090 168.315 74.260 ;
        RECT 168.520 74.090 169.375 74.260 ;
        RECT 170.250 73.870 170.580 74.330 ;
        RECT 170.790 74.230 171.050 74.620 ;
        RECT 171.240 75.440 172.205 75.450 ;
        RECT 172.375 75.530 172.545 75.910 ;
        RECT 173.135 75.870 173.305 76.160 ;
        RECT 173.485 76.040 173.815 76.420 ;
        RECT 173.135 75.700 173.935 75.870 ;
        RECT 171.240 75.280 171.915 75.440 ;
        RECT 172.375 75.360 173.595 75.530 ;
        RECT 171.240 74.490 171.450 75.280 ;
        RECT 172.375 75.270 172.545 75.360 ;
        RECT 171.620 74.490 171.970 75.110 ;
        RECT 172.140 75.100 172.545 75.270 ;
        RECT 172.140 74.320 172.310 75.100 ;
        RECT 172.480 74.650 172.700 74.930 ;
        RECT 172.880 74.820 173.420 75.190 ;
        RECT 173.765 75.110 173.935 75.700 ;
        RECT 174.155 75.280 174.460 76.420 ;
        RECT 174.630 75.230 174.885 76.110 ;
        RECT 175.060 75.255 175.350 76.420 ;
        RECT 175.520 75.330 179.030 76.420 ;
        RECT 179.205 75.750 179.460 76.250 ;
        RECT 179.630 75.920 179.960 76.420 ;
        RECT 179.205 75.580 179.955 75.750 ;
        RECT 173.765 75.080 174.505 75.110 ;
        RECT 172.480 74.480 173.010 74.650 ;
        RECT 170.790 74.060 171.140 74.230 ;
        RECT 171.360 74.040 172.310 74.320 ;
        RECT 172.480 73.870 172.670 74.310 ;
        RECT 172.840 74.250 173.010 74.480 ;
        RECT 173.180 74.420 173.420 74.820 ;
        RECT 173.590 74.780 174.505 75.080 ;
        RECT 173.590 74.605 173.915 74.780 ;
        RECT 173.590 74.250 173.910 74.605 ;
        RECT 174.675 74.580 174.885 75.230 ;
        RECT 175.520 74.640 177.170 75.160 ;
        RECT 177.340 74.810 179.030 75.330 ;
        RECT 179.205 74.760 179.555 75.410 ;
        RECT 172.840 74.080 173.910 74.250 ;
        RECT 174.155 73.870 174.460 74.330 ;
        RECT 174.630 74.050 174.885 74.580 ;
        RECT 175.060 73.870 175.350 74.595 ;
        RECT 175.520 73.870 179.030 74.640 ;
        RECT 179.725 74.590 179.955 75.580 ;
        RECT 179.205 74.420 179.955 74.590 ;
        RECT 179.205 74.130 179.460 74.420 ;
        RECT 179.630 73.870 179.960 74.250 ;
        RECT 180.130 74.130 180.300 76.250 ;
        RECT 180.470 75.450 180.795 76.235 ;
        RECT 180.965 75.960 181.215 76.420 ;
        RECT 181.385 75.920 181.635 76.250 ;
        RECT 181.850 75.920 182.530 76.250 ;
        RECT 181.385 75.790 181.555 75.920 ;
        RECT 181.160 75.620 181.555 75.790 ;
        RECT 180.530 74.400 180.990 75.450 ;
        RECT 181.160 74.260 181.330 75.620 ;
        RECT 181.725 75.360 182.190 75.750 ;
        RECT 181.500 74.550 181.850 75.170 ;
        RECT 182.020 74.770 182.190 75.360 ;
        RECT 182.360 75.140 182.530 75.920 ;
        RECT 182.700 75.820 182.870 76.160 ;
        RECT 183.105 75.990 183.435 76.420 ;
        RECT 183.605 75.820 183.775 76.160 ;
        RECT 184.070 75.960 184.440 76.420 ;
        RECT 182.700 75.650 183.775 75.820 ;
        RECT 184.610 75.790 184.780 76.250 ;
        RECT 185.015 75.910 185.885 76.250 ;
        RECT 186.055 75.960 186.305 76.420 ;
        RECT 184.220 75.620 184.780 75.790 ;
        RECT 184.220 75.480 184.390 75.620 ;
        RECT 182.890 75.310 184.390 75.480 ;
        RECT 185.085 75.450 185.545 75.740 ;
        RECT 182.360 74.970 184.050 75.140 ;
        RECT 182.020 74.550 182.375 74.770 ;
        RECT 182.545 74.260 182.715 74.970 ;
        RECT 182.920 74.550 183.710 74.800 ;
        RECT 183.880 74.790 184.050 74.970 ;
        RECT 184.220 74.620 184.390 75.310 ;
        RECT 180.660 73.870 180.990 74.230 ;
        RECT 181.160 74.090 181.655 74.260 ;
        RECT 181.860 74.090 182.715 74.260 ;
        RECT 183.590 73.870 183.920 74.330 ;
        RECT 184.130 74.230 184.390 74.620 ;
        RECT 184.580 75.440 185.545 75.450 ;
        RECT 185.715 75.530 185.885 75.910 ;
        RECT 186.475 75.870 186.645 76.160 ;
        RECT 186.825 76.040 187.155 76.420 ;
        RECT 186.475 75.700 187.275 75.870 ;
        RECT 184.580 75.280 185.255 75.440 ;
        RECT 185.715 75.360 186.935 75.530 ;
        RECT 184.580 74.490 184.790 75.280 ;
        RECT 185.715 75.270 185.885 75.360 ;
        RECT 184.960 74.490 185.310 75.110 ;
        RECT 185.480 75.100 185.885 75.270 ;
        RECT 185.480 74.320 185.650 75.100 ;
        RECT 185.820 74.650 186.040 74.930 ;
        RECT 186.220 74.820 186.760 75.190 ;
        RECT 187.105 75.110 187.275 75.700 ;
        RECT 187.495 75.280 187.800 76.420 ;
        RECT 187.970 75.230 188.225 76.110 ;
        RECT 188.410 75.355 188.720 76.420 ;
        RECT 188.890 75.750 189.125 76.250 ;
        RECT 189.295 75.960 189.625 76.420 ;
        RECT 189.820 76.080 190.930 76.250 ;
        RECT 189.820 75.920 190.010 76.080 ;
        RECT 190.240 75.750 190.540 75.910 ;
        RECT 188.890 75.570 190.540 75.750 ;
        RECT 190.710 75.570 190.930 76.080 ;
        RECT 191.100 75.570 191.430 76.420 ;
        RECT 187.105 75.080 187.845 75.110 ;
        RECT 185.820 74.480 186.350 74.650 ;
        RECT 184.130 74.060 184.480 74.230 ;
        RECT 184.700 74.040 185.650 74.320 ;
        RECT 185.820 73.870 186.010 74.310 ;
        RECT 186.180 74.250 186.350 74.480 ;
        RECT 186.520 74.420 186.760 74.820 ;
        RECT 186.930 74.780 187.845 75.080 ;
        RECT 186.930 74.605 187.255 74.780 ;
        RECT 186.930 74.250 187.250 74.605 ;
        RECT 188.015 74.580 188.225 75.230 ;
        RECT 186.180 74.080 187.250 74.250 ;
        RECT 187.495 73.870 187.800 74.330 ;
        RECT 187.970 74.050 188.225 74.580 ;
        RECT 188.405 74.550 188.720 75.185 ;
        RECT 188.890 74.380 189.100 75.570 ;
        RECT 189.440 75.230 191.415 75.400 ;
        RECT 189.440 74.860 189.935 75.230 ;
        RECT 190.115 74.860 190.915 75.060 ;
        RECT 191.085 74.840 191.415 75.230 ;
        RECT 191.625 75.230 191.880 76.110 ;
        RECT 192.050 75.280 192.355 76.420 ;
        RECT 192.695 76.040 193.025 76.420 ;
        RECT 193.205 75.870 193.375 76.160 ;
        RECT 193.545 75.960 193.795 76.420 ;
        RECT 192.575 75.700 193.375 75.870 ;
        RECT 193.965 75.910 194.835 76.250 ;
        RECT 189.270 74.500 191.430 74.670 ;
        RECT 188.410 74.210 188.720 74.380 ;
        RECT 189.270 74.210 189.600 74.500 ;
        RECT 188.410 74.040 189.600 74.210 ;
        RECT 189.840 73.870 190.010 74.330 ;
        RECT 190.240 74.040 190.570 74.500 ;
        RECT 190.750 73.870 190.920 74.330 ;
        RECT 191.100 74.040 191.430 74.500 ;
        RECT 191.625 74.580 191.835 75.230 ;
        RECT 192.575 75.110 192.745 75.700 ;
        RECT 193.965 75.530 194.135 75.910 ;
        RECT 195.070 75.790 195.240 76.250 ;
        RECT 195.410 75.960 195.780 76.420 ;
        RECT 196.075 75.820 196.245 76.160 ;
        RECT 196.415 75.990 196.745 76.420 ;
        RECT 196.980 75.820 197.150 76.160 ;
        RECT 192.915 75.360 194.135 75.530 ;
        RECT 194.305 75.450 194.765 75.740 ;
        RECT 195.070 75.620 195.630 75.790 ;
        RECT 196.075 75.650 197.150 75.820 ;
        RECT 197.320 75.920 198.000 76.250 ;
        RECT 198.215 75.920 198.465 76.250 ;
        RECT 198.635 75.960 198.885 76.420 ;
        RECT 195.460 75.480 195.630 75.620 ;
        RECT 194.305 75.440 195.270 75.450 ;
        RECT 193.965 75.270 194.135 75.360 ;
        RECT 194.595 75.280 195.270 75.440 ;
        RECT 192.005 75.080 192.745 75.110 ;
        RECT 192.005 74.780 192.920 75.080 ;
        RECT 192.595 74.605 192.920 74.780 ;
        RECT 191.625 74.050 191.880 74.580 ;
        RECT 192.050 73.870 192.355 74.330 ;
        RECT 192.600 74.250 192.920 74.605 ;
        RECT 193.090 74.820 193.630 75.190 ;
        RECT 193.965 75.100 194.370 75.270 ;
        RECT 193.090 74.420 193.330 74.820 ;
        RECT 193.810 74.650 194.030 74.930 ;
        RECT 193.500 74.480 194.030 74.650 ;
        RECT 193.500 74.250 193.670 74.480 ;
        RECT 194.200 74.320 194.370 75.100 ;
        RECT 194.540 74.490 194.890 75.110 ;
        RECT 195.060 74.490 195.270 75.280 ;
        RECT 195.460 75.310 196.960 75.480 ;
        RECT 195.460 74.620 195.630 75.310 ;
        RECT 197.320 75.140 197.490 75.920 ;
        RECT 198.295 75.790 198.465 75.920 ;
        RECT 195.800 74.970 197.490 75.140 ;
        RECT 197.660 75.360 198.125 75.750 ;
        RECT 198.295 75.620 198.690 75.790 ;
        RECT 195.800 74.790 195.970 74.970 ;
        RECT 192.600 74.080 193.670 74.250 ;
        RECT 193.840 73.870 194.030 74.310 ;
        RECT 194.200 74.040 195.150 74.320 ;
        RECT 195.460 74.230 195.720 74.620 ;
        RECT 196.140 74.550 196.930 74.800 ;
        RECT 195.370 74.060 195.720 74.230 ;
        RECT 195.930 73.870 196.260 74.330 ;
        RECT 197.135 74.260 197.305 74.970 ;
        RECT 197.660 74.770 197.830 75.360 ;
        RECT 197.475 74.550 197.830 74.770 ;
        RECT 198.000 74.550 198.350 75.170 ;
        RECT 198.520 74.260 198.690 75.620 ;
        RECT 199.055 75.450 199.380 76.235 ;
        RECT 198.860 74.400 199.320 75.450 ;
        RECT 197.135 74.090 197.990 74.260 ;
        RECT 198.195 74.090 198.690 74.260 ;
        RECT 198.860 73.870 199.190 74.230 ;
        RECT 199.550 74.130 199.720 76.250 ;
        RECT 199.890 75.920 200.220 76.420 ;
        RECT 200.390 75.750 200.645 76.250 ;
        RECT 199.895 75.580 200.645 75.750 ;
        RECT 199.895 74.590 200.125 75.580 ;
        RECT 200.295 74.760 200.645 75.410 ;
        RECT 200.820 75.255 201.110 76.420 ;
        RECT 201.285 75.280 201.620 76.250 ;
        RECT 201.790 75.280 201.960 76.420 ;
        RECT 202.130 76.080 204.160 76.250 ;
        RECT 201.285 74.610 201.455 75.280 ;
        RECT 202.130 75.110 202.300 76.080 ;
        RECT 201.625 74.780 201.880 75.110 ;
        RECT 202.105 74.780 202.300 75.110 ;
        RECT 202.470 75.740 203.595 75.910 ;
        RECT 201.710 74.610 201.880 74.780 ;
        RECT 202.470 74.610 202.640 75.740 ;
        RECT 199.895 74.420 200.645 74.590 ;
        RECT 199.890 73.870 200.220 74.250 ;
        RECT 200.390 74.130 200.645 74.420 ;
        RECT 200.820 73.870 201.110 74.595 ;
        RECT 201.285 74.040 201.540 74.610 ;
        RECT 201.710 74.440 202.640 74.610 ;
        RECT 202.810 75.400 203.820 75.570 ;
        RECT 202.810 74.600 202.980 75.400 ;
        RECT 202.465 74.405 202.640 74.440 ;
        RECT 201.710 73.870 202.040 74.270 ;
        RECT 202.465 74.040 202.995 74.405 ;
        RECT 203.185 74.380 203.460 75.200 ;
        RECT 203.180 74.210 203.460 74.380 ;
        RECT 203.185 74.040 203.460 74.210 ;
        RECT 203.630 74.040 203.820 75.400 ;
        RECT 203.990 75.415 204.160 76.080 ;
        RECT 204.330 75.660 204.500 76.420 ;
        RECT 204.735 75.660 205.250 76.070 ;
        RECT 203.990 75.225 204.740 75.415 ;
        RECT 204.910 74.850 205.250 75.660 ;
        RECT 205.475 75.550 205.760 76.420 ;
        RECT 205.930 75.790 206.190 76.250 ;
        RECT 206.365 75.960 206.620 76.420 ;
        RECT 206.790 75.790 207.050 76.250 ;
        RECT 205.930 75.620 207.050 75.790 ;
        RECT 207.220 75.620 207.530 76.420 ;
        RECT 205.930 75.370 206.190 75.620 ;
        RECT 207.700 75.450 208.010 76.250 ;
        RECT 204.020 74.680 205.250 74.850 ;
        RECT 205.435 75.200 206.190 75.370 ;
        RECT 206.980 75.280 208.010 75.450 ;
        RECT 208.180 75.330 209.850 76.420 ;
        RECT 205.435 74.690 205.840 75.200 ;
        RECT 206.980 75.030 207.150 75.280 ;
        RECT 206.010 74.860 207.150 75.030 ;
        RECT 204.000 73.870 204.510 74.405 ;
        RECT 204.730 74.075 204.975 74.680 ;
        RECT 205.435 74.520 207.085 74.690 ;
        RECT 207.320 74.540 207.670 75.110 ;
        RECT 205.480 73.870 205.760 74.350 ;
        RECT 205.930 74.130 206.190 74.520 ;
        RECT 206.365 73.870 206.620 74.350 ;
        RECT 206.790 74.130 207.085 74.520 ;
        RECT 207.840 74.370 208.010 75.280 ;
        RECT 207.265 73.870 207.540 74.350 ;
        RECT 207.710 74.040 208.010 74.370 ;
        RECT 208.180 74.640 208.930 75.160 ;
        RECT 209.100 74.810 209.850 75.330 ;
        RECT 210.480 75.660 210.995 76.070 ;
        RECT 211.230 75.660 211.400 76.420 ;
        RECT 211.570 76.080 213.600 76.250 ;
        RECT 210.480 74.850 210.820 75.660 ;
        RECT 211.570 75.415 211.740 76.080 ;
        RECT 212.135 75.740 213.260 75.910 ;
        RECT 210.990 75.225 211.740 75.415 ;
        RECT 211.910 75.400 212.920 75.570 ;
        RECT 210.480 74.680 211.710 74.850 ;
        RECT 208.180 73.870 209.850 74.640 ;
        RECT 210.755 74.075 211.000 74.680 ;
        RECT 211.220 73.870 211.730 74.405 ;
        RECT 211.910 74.040 212.100 75.400 ;
        RECT 212.270 74.720 212.545 75.200 ;
        RECT 212.270 74.550 212.550 74.720 ;
        RECT 212.750 74.600 212.920 75.400 ;
        RECT 213.090 74.610 213.260 75.740 ;
        RECT 213.430 75.110 213.600 76.080 ;
        RECT 213.770 75.280 213.940 76.420 ;
        RECT 214.110 75.280 214.445 76.250 ;
        RECT 214.625 75.750 214.880 76.250 ;
        RECT 215.050 75.920 215.380 76.420 ;
        RECT 214.625 75.580 215.375 75.750 ;
        RECT 213.430 74.780 213.625 75.110 ;
        RECT 213.850 74.780 214.105 75.110 ;
        RECT 213.850 74.610 214.020 74.780 ;
        RECT 214.275 74.610 214.445 75.280 ;
        RECT 214.625 74.760 214.975 75.410 ;
        RECT 212.270 74.040 212.545 74.550 ;
        RECT 213.090 74.440 214.020 74.610 ;
        RECT 213.090 74.405 213.265 74.440 ;
        RECT 212.735 74.040 213.265 74.405 ;
        RECT 213.690 73.870 214.020 74.270 ;
        RECT 214.190 74.040 214.445 74.610 ;
        RECT 215.145 74.590 215.375 75.580 ;
        RECT 214.625 74.420 215.375 74.590 ;
        RECT 214.625 74.130 214.880 74.420 ;
        RECT 215.050 73.870 215.380 74.250 ;
        RECT 215.550 74.130 215.720 76.250 ;
        RECT 215.890 75.450 216.215 76.235 ;
        RECT 216.385 75.960 216.635 76.420 ;
        RECT 216.805 75.920 217.055 76.250 ;
        RECT 217.270 75.920 217.950 76.250 ;
        RECT 216.805 75.790 216.975 75.920 ;
        RECT 216.580 75.620 216.975 75.790 ;
        RECT 215.950 74.400 216.410 75.450 ;
        RECT 216.580 74.260 216.750 75.620 ;
        RECT 217.145 75.360 217.610 75.750 ;
        RECT 216.920 74.550 217.270 75.170 ;
        RECT 217.440 74.770 217.610 75.360 ;
        RECT 217.780 75.140 217.950 75.920 ;
        RECT 218.120 75.820 218.290 76.160 ;
        RECT 218.525 75.990 218.855 76.420 ;
        RECT 219.025 75.820 219.195 76.160 ;
        RECT 219.490 75.960 219.860 76.420 ;
        RECT 218.120 75.650 219.195 75.820 ;
        RECT 220.030 75.790 220.200 76.250 ;
        RECT 220.435 75.910 221.305 76.250 ;
        RECT 221.475 75.960 221.725 76.420 ;
        RECT 219.640 75.620 220.200 75.790 ;
        RECT 219.640 75.480 219.810 75.620 ;
        RECT 218.310 75.310 219.810 75.480 ;
        RECT 220.505 75.450 220.965 75.740 ;
        RECT 217.780 74.970 219.470 75.140 ;
        RECT 217.440 74.550 217.795 74.770 ;
        RECT 217.965 74.260 218.135 74.970 ;
        RECT 218.340 74.550 219.130 74.800 ;
        RECT 219.300 74.790 219.470 74.970 ;
        RECT 219.640 74.620 219.810 75.310 ;
        RECT 216.080 73.870 216.410 74.230 ;
        RECT 216.580 74.090 217.075 74.260 ;
        RECT 217.280 74.090 218.135 74.260 ;
        RECT 219.010 73.870 219.340 74.330 ;
        RECT 219.550 74.230 219.810 74.620 ;
        RECT 220.000 75.440 220.965 75.450 ;
        RECT 221.135 75.530 221.305 75.910 ;
        RECT 221.895 75.870 222.065 76.160 ;
        RECT 222.245 76.040 222.575 76.420 ;
        RECT 221.895 75.700 222.695 75.870 ;
        RECT 220.000 75.280 220.675 75.440 ;
        RECT 221.135 75.360 222.355 75.530 ;
        RECT 220.000 74.490 220.210 75.280 ;
        RECT 221.135 75.270 221.305 75.360 ;
        RECT 220.380 74.490 220.730 75.110 ;
        RECT 220.900 75.100 221.305 75.270 ;
        RECT 220.900 74.320 221.070 75.100 ;
        RECT 221.240 74.650 221.460 74.930 ;
        RECT 221.640 74.820 222.180 75.190 ;
        RECT 222.525 75.110 222.695 75.700 ;
        RECT 222.915 75.280 223.220 76.420 ;
        RECT 223.390 75.230 223.645 76.110 ;
        RECT 223.825 75.270 224.085 76.420 ;
        RECT 224.260 75.345 224.515 76.250 ;
        RECT 224.685 75.660 225.015 76.420 ;
        RECT 225.230 75.490 225.400 76.250 ;
        RECT 222.525 75.080 223.265 75.110 ;
        RECT 221.240 74.480 221.770 74.650 ;
        RECT 219.550 74.060 219.900 74.230 ;
        RECT 220.120 74.040 221.070 74.320 ;
        RECT 221.240 73.870 221.430 74.310 ;
        RECT 221.600 74.250 221.770 74.480 ;
        RECT 221.940 74.420 222.180 74.820 ;
        RECT 222.350 74.780 223.265 75.080 ;
        RECT 222.350 74.605 222.675 74.780 ;
        RECT 222.350 74.250 222.670 74.605 ;
        RECT 223.435 74.580 223.645 75.230 ;
        RECT 221.600 74.080 222.670 74.250 ;
        RECT 222.915 73.870 223.220 74.330 ;
        RECT 223.390 74.050 223.645 74.580 ;
        RECT 223.825 73.870 224.085 74.710 ;
        RECT 224.260 74.615 224.430 75.345 ;
        RECT 224.685 75.320 225.400 75.490 ;
        RECT 224.685 75.110 224.855 75.320 ;
        RECT 226.580 75.255 226.870 76.420 ;
        RECT 227.040 75.985 232.385 76.420 ;
        RECT 224.600 74.780 224.855 75.110 ;
        RECT 224.260 74.040 224.515 74.615 ;
        RECT 224.685 74.590 224.855 74.780 ;
        RECT 225.135 74.770 225.490 75.140 ;
        RECT 224.685 74.420 225.400 74.590 ;
        RECT 224.685 73.870 225.015 74.250 ;
        RECT 225.230 74.040 225.400 74.420 ;
        RECT 226.580 73.870 226.870 74.595 ;
        RECT 228.625 74.415 228.965 75.245 ;
        RECT 230.445 74.735 230.795 75.985 ;
        RECT 232.560 75.330 236.070 76.420 ;
        RECT 232.560 74.640 234.210 75.160 ;
        RECT 234.380 74.810 236.070 75.330 ;
        RECT 236.245 75.280 236.520 76.250 ;
        RECT 236.730 75.620 237.010 76.420 ;
        RECT 237.180 75.910 238.370 76.200 ;
        RECT 238.540 75.985 243.885 76.420 ;
        RECT 244.060 75.985 249.405 76.420 ;
        RECT 237.180 75.570 238.350 75.740 ;
        RECT 237.180 75.450 237.350 75.570 ;
        RECT 236.690 75.280 237.350 75.450 ;
        RECT 227.040 73.870 232.385 74.415 ;
        RECT 232.560 73.870 236.070 74.640 ;
        RECT 236.245 74.545 236.415 75.280 ;
        RECT 236.690 75.110 236.860 75.280 ;
        RECT 237.660 75.110 237.855 75.400 ;
        RECT 238.025 75.280 238.350 75.570 ;
        RECT 236.585 74.780 236.860 75.110 ;
        RECT 237.030 74.780 237.855 75.110 ;
        RECT 238.025 74.780 238.370 75.110 ;
        RECT 236.690 74.610 236.860 74.780 ;
        RECT 236.245 74.200 236.520 74.545 ;
        RECT 236.690 74.440 238.355 74.610 ;
        RECT 236.710 73.870 237.090 74.270 ;
        RECT 237.260 74.090 237.430 74.440 ;
        RECT 237.600 73.870 237.930 74.270 ;
        RECT 238.100 74.090 238.355 74.440 ;
        RECT 240.125 74.415 240.465 75.245 ;
        RECT 241.945 74.735 242.295 75.985 ;
        RECT 245.645 74.415 245.985 75.245 ;
        RECT 247.465 74.735 247.815 75.985 ;
        RECT 249.580 75.330 252.170 76.420 ;
        RECT 249.580 74.640 250.790 75.160 ;
        RECT 250.960 74.810 252.170 75.330 ;
        RECT 252.340 75.255 252.630 76.420 ;
        RECT 252.800 75.330 256.310 76.420 ;
        RECT 256.480 75.330 257.690 76.420 ;
        RECT 252.800 74.640 254.450 75.160 ;
        RECT 254.620 74.810 256.310 75.330 ;
        RECT 238.540 73.870 243.885 74.415 ;
        RECT 244.060 73.870 249.405 74.415 ;
        RECT 249.580 73.870 252.170 74.640 ;
        RECT 252.340 73.870 252.630 74.595 ;
        RECT 252.800 73.870 256.310 74.640 ;
        RECT 256.480 74.620 257.000 75.160 ;
        RECT 257.170 74.790 257.690 75.330 ;
        RECT 257.950 75.410 258.120 76.250 ;
        RECT 258.290 76.080 259.460 76.250 ;
        RECT 258.290 75.580 258.620 76.080 ;
        RECT 259.130 76.040 259.460 76.080 ;
        RECT 259.650 76.000 260.005 76.420 ;
        RECT 258.790 75.820 259.020 75.910 ;
        RECT 260.175 75.820 260.425 76.250 ;
        RECT 258.790 75.580 260.425 75.820 ;
        RECT 260.595 75.660 260.925 76.420 ;
        RECT 261.095 75.580 261.350 76.250 ;
        RECT 257.950 75.240 261.010 75.410 ;
        RECT 257.865 74.860 258.215 75.070 ;
        RECT 258.385 74.860 258.830 75.060 ;
        RECT 259.000 74.860 259.475 75.060 ;
        RECT 256.480 73.870 257.690 74.620 ;
        RECT 257.950 74.520 259.015 74.690 ;
        RECT 257.950 74.040 258.120 74.520 ;
        RECT 258.290 73.870 258.620 74.350 ;
        RECT 258.845 74.290 259.015 74.520 ;
        RECT 259.195 74.460 259.475 74.860 ;
        RECT 259.745 74.860 260.075 75.060 ;
        RECT 260.245 74.890 260.620 75.060 ;
        RECT 260.245 74.860 260.610 74.890 ;
        RECT 259.745 74.460 260.030 74.860 ;
        RECT 260.840 74.690 261.010 75.240 ;
        RECT 260.210 74.520 261.010 74.690 ;
        RECT 260.210 74.290 260.380 74.520 ;
        RECT 261.180 74.450 261.350 75.580 ;
        RECT 261.545 76.030 261.880 76.250 ;
        RECT 262.885 76.040 263.240 76.420 ;
        RECT 261.545 75.410 261.800 76.030 ;
        RECT 262.050 75.870 262.280 75.910 ;
        RECT 263.410 75.870 263.660 76.250 ;
        RECT 262.050 75.670 263.660 75.870 ;
        RECT 262.050 75.580 262.235 75.670 ;
        RECT 262.825 75.660 263.660 75.670 ;
        RECT 263.910 75.640 264.160 76.420 ;
        RECT 264.330 75.570 264.590 76.250 ;
        RECT 264.760 75.985 270.105 76.420 ;
        RECT 262.390 75.470 262.720 75.500 ;
        RECT 262.390 75.410 264.190 75.470 ;
        RECT 261.545 75.300 264.250 75.410 ;
        RECT 261.545 75.240 262.720 75.300 ;
        RECT 264.050 75.265 264.250 75.300 ;
        RECT 261.540 74.860 262.030 75.060 ;
        RECT 262.220 74.860 262.695 75.070 ;
        RECT 261.165 74.380 261.350 74.450 ;
        RECT 261.140 74.370 261.350 74.380 ;
        RECT 258.845 74.040 260.380 74.290 ;
        RECT 260.550 73.870 260.880 74.350 ;
        RECT 261.095 74.040 261.350 74.370 ;
        RECT 261.545 73.870 262.000 74.635 ;
        RECT 262.475 74.460 262.695 74.860 ;
        RECT 262.940 74.860 263.270 75.070 ;
        RECT 262.940 74.460 263.150 74.860 ;
        RECT 263.440 74.825 263.850 75.130 ;
        RECT 264.080 74.690 264.250 75.265 ;
        RECT 263.980 74.570 264.250 74.690 ;
        RECT 263.405 74.525 264.250 74.570 ;
        RECT 263.405 74.400 264.160 74.525 ;
        RECT 263.405 74.250 263.575 74.400 ;
        RECT 264.420 74.380 264.590 75.570 ;
        RECT 266.345 74.415 266.685 75.245 ;
        RECT 268.165 74.735 268.515 75.985 ;
        RECT 270.280 75.330 273.790 76.420 ;
        RECT 270.280 74.640 271.930 75.160 ;
        RECT 272.100 74.810 273.790 75.330 ;
        RECT 273.960 75.660 274.475 76.070 ;
        RECT 274.710 75.660 274.880 76.420 ;
        RECT 275.050 76.080 277.080 76.250 ;
        RECT 273.960 74.850 274.300 75.660 ;
        RECT 275.050 75.415 275.220 76.080 ;
        RECT 275.615 75.740 276.740 75.910 ;
        RECT 274.470 75.225 275.220 75.415 ;
        RECT 275.390 75.400 276.400 75.570 ;
        RECT 273.960 74.680 275.190 74.850 ;
        RECT 264.360 74.370 264.590 74.380 ;
        RECT 262.275 74.040 263.575 74.250 ;
        RECT 263.830 73.870 264.160 74.230 ;
        RECT 264.330 74.040 264.590 74.370 ;
        RECT 264.760 73.870 270.105 74.415 ;
        RECT 270.280 73.870 273.790 74.640 ;
        RECT 274.235 74.075 274.480 74.680 ;
        RECT 274.700 73.870 275.210 74.405 ;
        RECT 275.390 74.040 275.580 75.400 ;
        RECT 275.750 75.060 276.025 75.200 ;
        RECT 275.750 74.890 276.030 75.060 ;
        RECT 275.750 74.040 276.025 74.890 ;
        RECT 276.230 74.600 276.400 75.400 ;
        RECT 276.570 74.610 276.740 75.740 ;
        RECT 276.910 75.110 277.080 76.080 ;
        RECT 277.250 75.280 277.420 76.420 ;
        RECT 277.590 75.280 277.925 76.250 ;
        RECT 276.910 74.780 277.105 75.110 ;
        RECT 277.330 74.780 277.585 75.110 ;
        RECT 277.330 74.610 277.500 74.780 ;
        RECT 277.755 74.610 277.925 75.280 ;
        RECT 278.100 75.255 278.390 76.420 ;
        RECT 279.025 75.750 279.280 76.250 ;
        RECT 279.450 75.920 279.780 76.420 ;
        RECT 279.025 75.580 279.775 75.750 ;
        RECT 279.025 74.760 279.375 75.410 ;
        RECT 276.570 74.440 277.500 74.610 ;
        RECT 276.570 74.405 276.745 74.440 ;
        RECT 276.215 74.040 276.745 74.405 ;
        RECT 277.170 73.870 277.500 74.270 ;
        RECT 277.670 74.040 277.925 74.610 ;
        RECT 278.100 73.870 278.390 74.595 ;
        RECT 279.545 74.590 279.775 75.580 ;
        RECT 279.025 74.420 279.775 74.590 ;
        RECT 279.025 74.130 279.280 74.420 ;
        RECT 279.450 73.870 279.780 74.250 ;
        RECT 279.950 74.130 280.120 76.250 ;
        RECT 280.290 75.450 280.615 76.235 ;
        RECT 280.785 75.960 281.035 76.420 ;
        RECT 281.205 75.920 281.455 76.250 ;
        RECT 281.670 75.920 282.350 76.250 ;
        RECT 281.205 75.790 281.375 75.920 ;
        RECT 280.980 75.620 281.375 75.790 ;
        RECT 280.350 74.400 280.810 75.450 ;
        RECT 280.980 74.260 281.150 75.620 ;
        RECT 281.545 75.360 282.010 75.750 ;
        RECT 281.320 74.550 281.670 75.170 ;
        RECT 281.840 74.770 282.010 75.360 ;
        RECT 282.180 75.140 282.350 75.920 ;
        RECT 282.520 75.820 282.690 76.160 ;
        RECT 282.925 75.990 283.255 76.420 ;
        RECT 283.425 75.820 283.595 76.160 ;
        RECT 283.890 75.960 284.260 76.420 ;
        RECT 282.520 75.650 283.595 75.820 ;
        RECT 284.430 75.790 284.600 76.250 ;
        RECT 284.835 75.910 285.705 76.250 ;
        RECT 285.875 75.960 286.125 76.420 ;
        RECT 284.040 75.620 284.600 75.790 ;
        RECT 284.040 75.480 284.210 75.620 ;
        RECT 282.710 75.310 284.210 75.480 ;
        RECT 284.905 75.450 285.365 75.740 ;
        RECT 282.180 74.970 283.870 75.140 ;
        RECT 281.840 74.550 282.195 74.770 ;
        RECT 282.365 74.260 282.535 74.970 ;
        RECT 282.740 74.550 283.530 74.800 ;
        RECT 283.700 74.790 283.870 74.970 ;
        RECT 284.040 74.620 284.210 75.310 ;
        RECT 280.480 73.870 280.810 74.230 ;
        RECT 280.980 74.090 281.475 74.260 ;
        RECT 281.680 74.090 282.535 74.260 ;
        RECT 283.410 73.870 283.740 74.330 ;
        RECT 283.950 74.230 284.210 74.620 ;
        RECT 284.400 75.440 285.365 75.450 ;
        RECT 285.535 75.530 285.705 75.910 ;
        RECT 286.295 75.870 286.465 76.160 ;
        RECT 286.645 76.040 286.975 76.420 ;
        RECT 286.295 75.700 287.095 75.870 ;
        RECT 284.400 75.280 285.075 75.440 ;
        RECT 285.535 75.360 286.755 75.530 ;
        RECT 284.400 74.490 284.610 75.280 ;
        RECT 285.535 75.270 285.705 75.360 ;
        RECT 284.780 74.490 285.130 75.110 ;
        RECT 285.300 75.100 285.705 75.270 ;
        RECT 285.300 74.320 285.470 75.100 ;
        RECT 285.640 74.650 285.860 74.930 ;
        RECT 286.040 74.820 286.580 75.190 ;
        RECT 286.925 75.110 287.095 75.700 ;
        RECT 287.315 75.280 287.620 76.420 ;
        RECT 287.790 75.230 288.045 76.110 ;
        RECT 288.220 75.330 289.890 76.420 ;
        RECT 286.925 75.080 287.665 75.110 ;
        RECT 285.640 74.480 286.170 74.650 ;
        RECT 283.950 74.060 284.300 74.230 ;
        RECT 284.520 74.040 285.470 74.320 ;
        RECT 285.640 73.870 285.830 74.310 ;
        RECT 286.000 74.250 286.170 74.480 ;
        RECT 286.340 74.420 286.580 74.820 ;
        RECT 286.750 74.780 287.665 75.080 ;
        RECT 286.750 74.605 287.075 74.780 ;
        RECT 286.750 74.250 287.070 74.605 ;
        RECT 287.835 74.580 288.045 75.230 ;
        RECT 286.000 74.080 287.070 74.250 ;
        RECT 287.315 73.870 287.620 74.330 ;
        RECT 287.790 74.050 288.045 74.580 ;
        RECT 288.220 74.640 288.970 75.160 ;
        RECT 289.140 74.810 289.890 75.330 ;
        RECT 290.520 75.660 291.035 76.070 ;
        RECT 291.270 75.660 291.440 76.420 ;
        RECT 291.610 76.080 293.640 76.250 ;
        RECT 290.520 74.850 290.860 75.660 ;
        RECT 291.610 75.415 291.780 76.080 ;
        RECT 292.175 75.740 293.300 75.910 ;
        RECT 291.030 75.225 291.780 75.415 ;
        RECT 291.950 75.400 292.960 75.570 ;
        RECT 290.520 74.680 291.750 74.850 ;
        RECT 288.220 73.870 289.890 74.640 ;
        RECT 290.795 74.075 291.040 74.680 ;
        RECT 291.260 73.870 291.770 74.405 ;
        RECT 291.950 74.040 292.140 75.400 ;
        RECT 292.310 75.060 292.585 75.200 ;
        RECT 292.310 74.890 292.590 75.060 ;
        RECT 292.310 74.040 292.585 74.890 ;
        RECT 292.790 74.600 292.960 75.400 ;
        RECT 293.130 74.610 293.300 75.740 ;
        RECT 293.470 75.110 293.640 76.080 ;
        RECT 293.810 75.280 293.980 76.420 ;
        RECT 294.150 75.280 294.485 76.250 ;
        RECT 293.470 74.780 293.665 75.110 ;
        RECT 293.890 74.780 294.145 75.110 ;
        RECT 293.890 74.610 294.060 74.780 ;
        RECT 294.315 74.610 294.485 75.280 ;
        RECT 293.130 74.440 294.060 74.610 ;
        RECT 293.130 74.405 293.305 74.440 ;
        RECT 292.775 74.040 293.305 74.405 ;
        RECT 293.730 73.870 294.060 74.270 ;
        RECT 294.230 74.040 294.485 74.610 ;
        RECT 294.665 75.230 294.920 76.110 ;
        RECT 295.090 75.280 295.395 76.420 ;
        RECT 295.735 76.040 296.065 76.420 ;
        RECT 296.245 75.870 296.415 76.160 ;
        RECT 296.585 75.960 296.835 76.420 ;
        RECT 295.615 75.700 296.415 75.870 ;
        RECT 297.005 75.910 297.875 76.250 ;
        RECT 294.665 74.580 294.875 75.230 ;
        RECT 295.615 75.110 295.785 75.700 ;
        RECT 297.005 75.530 297.175 75.910 ;
        RECT 298.110 75.790 298.280 76.250 ;
        RECT 298.450 75.960 298.820 76.420 ;
        RECT 299.115 75.820 299.285 76.160 ;
        RECT 299.455 75.990 299.785 76.420 ;
        RECT 300.020 75.820 300.190 76.160 ;
        RECT 295.955 75.360 297.175 75.530 ;
        RECT 297.345 75.450 297.805 75.740 ;
        RECT 298.110 75.620 298.670 75.790 ;
        RECT 299.115 75.650 300.190 75.820 ;
        RECT 300.360 75.920 301.040 76.250 ;
        RECT 301.255 75.920 301.505 76.250 ;
        RECT 301.675 75.960 301.925 76.420 ;
        RECT 298.500 75.480 298.670 75.620 ;
        RECT 297.345 75.440 298.310 75.450 ;
        RECT 297.005 75.270 297.175 75.360 ;
        RECT 297.635 75.280 298.310 75.440 ;
        RECT 295.045 75.080 295.785 75.110 ;
        RECT 295.045 74.780 295.960 75.080 ;
        RECT 295.635 74.605 295.960 74.780 ;
        RECT 294.665 74.050 294.920 74.580 ;
        RECT 295.090 73.870 295.395 74.330 ;
        RECT 295.640 74.250 295.960 74.605 ;
        RECT 296.130 74.820 296.670 75.190 ;
        RECT 297.005 75.100 297.410 75.270 ;
        RECT 296.130 74.420 296.370 74.820 ;
        RECT 296.850 74.650 297.070 74.930 ;
        RECT 296.540 74.480 297.070 74.650 ;
        RECT 296.540 74.250 296.710 74.480 ;
        RECT 297.240 74.320 297.410 75.100 ;
        RECT 297.580 74.490 297.930 75.110 ;
        RECT 298.100 74.490 298.310 75.280 ;
        RECT 298.500 75.310 300.000 75.480 ;
        RECT 298.500 74.620 298.670 75.310 ;
        RECT 300.360 75.140 300.530 75.920 ;
        RECT 301.335 75.790 301.505 75.920 ;
        RECT 298.840 74.970 300.530 75.140 ;
        RECT 300.700 75.360 301.165 75.750 ;
        RECT 301.335 75.620 301.730 75.790 ;
        RECT 298.840 74.790 299.010 74.970 ;
        RECT 295.640 74.080 296.710 74.250 ;
        RECT 296.880 73.870 297.070 74.310 ;
        RECT 297.240 74.040 298.190 74.320 ;
        RECT 298.500 74.230 298.760 74.620 ;
        RECT 299.180 74.550 299.970 74.800 ;
        RECT 298.410 74.060 298.760 74.230 ;
        RECT 298.970 73.870 299.300 74.330 ;
        RECT 300.175 74.260 300.345 74.970 ;
        RECT 300.700 74.770 300.870 75.360 ;
        RECT 300.515 74.550 300.870 74.770 ;
        RECT 301.040 74.550 301.390 75.170 ;
        RECT 301.560 74.260 301.730 75.620 ;
        RECT 302.095 75.450 302.420 76.235 ;
        RECT 301.900 74.400 302.360 75.450 ;
        RECT 300.175 74.090 301.030 74.260 ;
        RECT 301.235 74.090 301.730 74.260 ;
        RECT 301.900 73.870 302.230 74.230 ;
        RECT 302.590 74.130 302.760 76.250 ;
        RECT 302.930 75.920 303.260 76.420 ;
        RECT 303.430 75.750 303.685 76.250 ;
        RECT 302.935 75.580 303.685 75.750 ;
        RECT 302.935 74.590 303.165 75.580 ;
        RECT 303.335 74.760 303.685 75.410 ;
        RECT 303.860 75.255 304.150 76.420 ;
        RECT 304.320 75.985 309.665 76.420 ;
        RECT 302.935 74.420 303.685 74.590 ;
        RECT 302.930 73.870 303.260 74.250 ;
        RECT 303.430 74.130 303.685 74.420 ;
        RECT 303.860 73.870 304.150 74.595 ;
        RECT 305.905 74.415 306.245 75.245 ;
        RECT 307.725 74.735 308.075 75.985 ;
        RECT 309.840 75.330 311.050 76.420 ;
        RECT 309.840 74.790 310.360 75.330 ;
        RECT 310.530 74.620 311.050 75.160 ;
        RECT 304.320 73.870 309.665 74.415 ;
        RECT 309.840 73.870 311.050 74.620 ;
        RECT 162.095 73.700 311.135 73.870 ;
        RECT 162.180 72.950 163.390 73.700 ;
        RECT 162.180 72.410 162.700 72.950 ;
        RECT 163.560 72.930 167.070 73.700 ;
        RECT 168.210 72.945 168.460 73.700 ;
        RECT 168.630 72.990 168.880 73.520 ;
        RECT 169.050 73.240 169.355 73.700 ;
        RECT 169.600 73.320 170.670 73.490 ;
        RECT 162.870 72.240 163.390 72.780 ;
        RECT 163.560 72.410 165.210 72.930 ;
        RECT 165.380 72.240 167.070 72.760 ;
        RECT 168.630 72.340 168.835 72.990 ;
        RECT 169.600 72.965 169.920 73.320 ;
        RECT 169.595 72.790 169.920 72.965 ;
        RECT 169.005 72.490 169.920 72.790 ;
        RECT 170.090 72.750 170.330 73.150 ;
        RECT 170.500 73.090 170.670 73.320 ;
        RECT 170.840 73.260 171.030 73.700 ;
        RECT 171.200 73.250 172.150 73.530 ;
        RECT 172.370 73.340 172.720 73.510 ;
        RECT 170.500 72.920 171.030 73.090 ;
        RECT 169.005 72.460 169.745 72.490 ;
        RECT 162.180 71.150 163.390 72.240 ;
        RECT 163.560 71.150 167.070 72.240 ;
        RECT 168.210 71.150 168.460 72.290 ;
        RECT 168.630 71.460 168.880 72.340 ;
        RECT 169.050 71.150 169.355 72.290 ;
        RECT 169.575 71.870 169.745 72.460 ;
        RECT 170.090 72.380 170.630 72.750 ;
        RECT 170.810 72.640 171.030 72.920 ;
        RECT 171.200 72.470 171.370 73.250 ;
        RECT 170.965 72.300 171.370 72.470 ;
        RECT 171.540 72.460 171.890 73.080 ;
        RECT 170.965 72.210 171.135 72.300 ;
        RECT 172.060 72.290 172.270 73.080 ;
        RECT 169.915 72.040 171.135 72.210 ;
        RECT 171.595 72.130 172.270 72.290 ;
        RECT 169.575 71.700 170.375 71.870 ;
        RECT 169.695 71.150 170.025 71.530 ;
        RECT 170.205 71.410 170.375 71.700 ;
        RECT 170.965 71.660 171.135 72.040 ;
        RECT 171.305 72.120 172.270 72.130 ;
        RECT 172.460 72.950 172.720 73.340 ;
        RECT 172.930 73.240 173.260 73.700 ;
        RECT 174.135 73.310 174.990 73.480 ;
        RECT 175.195 73.310 175.690 73.480 ;
        RECT 175.860 73.340 176.190 73.700 ;
        RECT 172.460 72.260 172.630 72.950 ;
        RECT 172.800 72.600 172.970 72.780 ;
        RECT 173.140 72.770 173.930 73.020 ;
        RECT 174.135 72.600 174.305 73.310 ;
        RECT 174.475 72.800 174.830 73.020 ;
        RECT 172.800 72.430 174.490 72.600 ;
        RECT 171.305 71.830 171.765 72.120 ;
        RECT 172.460 72.090 173.960 72.260 ;
        RECT 172.460 71.950 172.630 72.090 ;
        RECT 172.070 71.780 172.630 71.950 ;
        RECT 170.545 71.150 170.795 71.610 ;
        RECT 170.965 71.320 171.835 71.660 ;
        RECT 172.070 71.320 172.240 71.780 ;
        RECT 173.075 71.750 174.150 71.920 ;
        RECT 172.410 71.150 172.780 71.610 ;
        RECT 173.075 71.410 173.245 71.750 ;
        RECT 173.415 71.150 173.745 71.580 ;
        RECT 173.980 71.410 174.150 71.750 ;
        RECT 174.320 71.650 174.490 72.430 ;
        RECT 174.660 72.210 174.830 72.800 ;
        RECT 175.000 72.400 175.350 73.020 ;
        RECT 174.660 71.820 175.125 72.210 ;
        RECT 175.520 71.950 175.690 73.310 ;
        RECT 175.860 72.120 176.320 73.170 ;
        RECT 175.295 71.780 175.690 71.950 ;
        RECT 175.295 71.650 175.465 71.780 ;
        RECT 174.320 71.320 175.000 71.650 ;
        RECT 175.215 71.320 175.465 71.650 ;
        RECT 175.635 71.150 175.885 71.610 ;
        RECT 176.055 71.335 176.380 72.120 ;
        RECT 176.550 71.320 176.720 73.440 ;
        RECT 176.890 73.320 177.220 73.700 ;
        RECT 177.390 73.150 177.645 73.440 ;
        RECT 176.895 72.980 177.645 73.150 ;
        RECT 176.895 71.990 177.125 72.980 ;
        RECT 177.825 72.960 178.080 73.530 ;
        RECT 178.250 73.300 178.580 73.700 ;
        RECT 179.005 73.165 179.535 73.530 ;
        RECT 179.005 73.130 179.180 73.165 ;
        RECT 178.250 72.960 179.180 73.130 ;
        RECT 177.295 72.160 177.645 72.810 ;
        RECT 177.825 72.290 177.995 72.960 ;
        RECT 178.250 72.790 178.420 72.960 ;
        RECT 178.165 72.460 178.420 72.790 ;
        RECT 178.645 72.460 178.840 72.790 ;
        RECT 176.895 71.820 177.645 71.990 ;
        RECT 176.890 71.150 177.220 71.650 ;
        RECT 177.390 71.320 177.645 71.820 ;
        RECT 177.825 71.320 178.160 72.290 ;
        RECT 178.330 71.150 178.500 72.290 ;
        RECT 178.670 71.490 178.840 72.460 ;
        RECT 179.010 71.830 179.180 72.960 ;
        RECT 179.350 72.170 179.520 72.970 ;
        RECT 179.725 72.680 180.000 73.530 ;
        RECT 179.720 72.510 180.000 72.680 ;
        RECT 179.725 72.370 180.000 72.510 ;
        RECT 180.170 72.170 180.360 73.530 ;
        RECT 180.540 73.165 181.050 73.700 ;
        RECT 181.270 72.890 181.515 73.495 ;
        RECT 182.885 72.960 183.140 73.530 ;
        RECT 183.310 73.300 183.640 73.700 ;
        RECT 184.065 73.165 184.595 73.530 ;
        RECT 184.065 73.130 184.240 73.165 ;
        RECT 183.310 72.960 184.240 73.130 ;
        RECT 180.560 72.720 181.790 72.890 ;
        RECT 179.350 72.000 180.360 72.170 ;
        RECT 180.530 72.155 181.280 72.345 ;
        RECT 179.010 71.660 180.135 71.830 ;
        RECT 180.530 71.490 180.700 72.155 ;
        RECT 181.450 71.910 181.790 72.720 ;
        RECT 178.670 71.320 180.700 71.490 ;
        RECT 180.870 71.150 181.040 71.910 ;
        RECT 181.275 71.500 181.790 71.910 ;
        RECT 182.885 72.290 183.055 72.960 ;
        RECT 183.310 72.790 183.480 72.960 ;
        RECT 183.225 72.460 183.480 72.790 ;
        RECT 183.705 72.460 183.900 72.790 ;
        RECT 182.885 71.320 183.220 72.290 ;
        RECT 183.390 71.150 183.560 72.290 ;
        RECT 183.730 71.490 183.900 72.460 ;
        RECT 184.070 71.830 184.240 72.960 ;
        RECT 184.410 72.170 184.580 72.970 ;
        RECT 184.785 72.680 185.060 73.530 ;
        RECT 184.780 72.510 185.060 72.680 ;
        RECT 184.785 72.370 185.060 72.510 ;
        RECT 185.230 72.170 185.420 73.530 ;
        RECT 185.600 73.165 186.110 73.700 ;
        RECT 186.330 72.890 186.575 73.495 ;
        RECT 187.940 72.975 188.230 73.700 ;
        RECT 188.460 73.240 188.705 73.700 ;
        RECT 185.620 72.720 186.850 72.890 ;
        RECT 184.410 72.000 185.420 72.170 ;
        RECT 185.590 72.155 186.340 72.345 ;
        RECT 184.070 71.660 185.195 71.830 ;
        RECT 185.590 71.490 185.760 72.155 ;
        RECT 186.510 71.910 186.850 72.720 ;
        RECT 188.400 72.460 188.715 73.070 ;
        RECT 188.885 72.710 189.135 73.520 ;
        RECT 189.305 73.175 189.565 73.700 ;
        RECT 189.735 73.050 189.995 73.505 ;
        RECT 190.165 73.220 190.425 73.700 ;
        RECT 190.595 73.050 190.855 73.505 ;
        RECT 191.025 73.220 191.285 73.700 ;
        RECT 191.455 73.050 191.715 73.505 ;
        RECT 191.885 73.220 192.145 73.700 ;
        RECT 192.315 73.050 192.575 73.505 ;
        RECT 192.745 73.220 193.045 73.700 ;
        RECT 193.505 73.240 193.770 73.700 ;
        RECT 194.140 73.060 194.310 73.530 ;
        RECT 194.560 73.240 194.730 73.700 ;
        RECT 194.980 73.060 195.150 73.530 ;
        RECT 195.400 73.240 195.570 73.700 ;
        RECT 195.820 73.060 195.990 73.530 ;
        RECT 196.160 73.235 196.410 73.700 ;
        RECT 197.145 73.150 197.400 73.440 ;
        RECT 197.570 73.320 197.900 73.700 ;
        RECT 189.735 72.880 193.045 73.050 ;
        RECT 194.140 72.880 196.510 73.060 ;
        RECT 197.145 72.980 197.895 73.150 ;
        RECT 188.885 72.460 191.905 72.710 ;
        RECT 183.730 71.320 185.760 71.490 ;
        RECT 185.930 71.150 186.100 71.910 ;
        RECT 186.335 71.500 186.850 71.910 ;
        RECT 187.940 71.150 188.230 72.315 ;
        RECT 188.410 71.150 188.705 72.260 ;
        RECT 188.885 71.325 189.135 72.460 ;
        RECT 192.075 72.290 193.045 72.880 ;
        RECT 193.480 72.460 195.990 72.710 ;
        RECT 196.160 72.290 196.510 72.880 ;
        RECT 189.305 71.150 189.565 72.260 ;
        RECT 189.735 72.050 193.045 72.290 ;
        RECT 189.735 71.325 189.995 72.050 ;
        RECT 190.165 71.150 190.425 71.880 ;
        RECT 190.595 71.325 190.855 72.050 ;
        RECT 191.025 71.150 191.285 71.880 ;
        RECT 191.455 71.325 191.715 72.050 ;
        RECT 191.885 71.150 192.145 71.880 ;
        RECT 192.315 71.325 192.575 72.050 ;
        RECT 192.745 71.150 193.040 71.880 ;
        RECT 193.505 71.150 193.800 72.290 ;
        RECT 194.060 72.120 196.510 72.290 ;
        RECT 197.145 72.160 197.495 72.810 ;
        RECT 194.060 71.320 194.390 72.120 ;
        RECT 194.560 71.150 194.730 71.950 ;
        RECT 194.900 71.320 195.230 72.120 ;
        RECT 195.740 72.100 196.510 72.120 ;
        RECT 195.400 71.150 195.570 71.950 ;
        RECT 195.740 71.320 196.070 72.100 ;
        RECT 197.665 71.990 197.895 72.980 ;
        RECT 197.145 71.820 197.895 71.990 ;
        RECT 196.240 71.150 196.410 71.610 ;
        RECT 197.145 71.320 197.400 71.820 ;
        RECT 197.570 71.150 197.900 71.650 ;
        RECT 198.070 71.320 198.240 73.440 ;
        RECT 198.600 73.340 198.930 73.700 ;
        RECT 199.100 73.310 199.595 73.480 ;
        RECT 199.800 73.310 200.655 73.480 ;
        RECT 198.470 72.120 198.930 73.170 ;
        RECT 198.410 71.335 198.735 72.120 ;
        RECT 199.100 71.950 199.270 73.310 ;
        RECT 199.440 72.400 199.790 73.020 ;
        RECT 199.960 72.800 200.315 73.020 ;
        RECT 199.960 72.210 200.130 72.800 ;
        RECT 200.485 72.600 200.655 73.310 ;
        RECT 201.530 73.240 201.860 73.700 ;
        RECT 202.070 73.340 202.420 73.510 ;
        RECT 200.860 72.770 201.650 73.020 ;
        RECT 202.070 72.950 202.330 73.340 ;
        RECT 202.640 73.250 203.590 73.530 ;
        RECT 203.760 73.260 203.950 73.700 ;
        RECT 204.120 73.320 205.190 73.490 ;
        RECT 201.820 72.600 201.990 72.780 ;
        RECT 199.100 71.780 199.495 71.950 ;
        RECT 199.665 71.820 200.130 72.210 ;
        RECT 200.300 72.430 201.990 72.600 ;
        RECT 199.325 71.650 199.495 71.780 ;
        RECT 200.300 71.650 200.470 72.430 ;
        RECT 202.160 72.260 202.330 72.950 ;
        RECT 200.830 72.090 202.330 72.260 ;
        RECT 202.520 72.290 202.730 73.080 ;
        RECT 202.900 72.460 203.250 73.080 ;
        RECT 203.420 72.470 203.590 73.250 ;
        RECT 204.120 73.090 204.290 73.320 ;
        RECT 203.760 72.920 204.290 73.090 ;
        RECT 203.760 72.640 203.980 72.920 ;
        RECT 204.460 72.750 204.700 73.150 ;
        RECT 203.420 72.300 203.825 72.470 ;
        RECT 204.160 72.380 204.700 72.750 ;
        RECT 204.870 72.965 205.190 73.320 ;
        RECT 205.435 73.240 205.740 73.700 ;
        RECT 205.910 72.990 206.165 73.520 ;
        RECT 206.350 73.360 207.540 73.530 ;
        RECT 206.350 73.190 206.660 73.360 ;
        RECT 204.870 72.790 205.195 72.965 ;
        RECT 204.870 72.490 205.785 72.790 ;
        RECT 205.045 72.460 205.785 72.490 ;
        RECT 202.520 72.130 203.195 72.290 ;
        RECT 203.655 72.210 203.825 72.300 ;
        RECT 202.520 72.120 203.485 72.130 ;
        RECT 202.160 71.950 202.330 72.090 ;
        RECT 198.905 71.150 199.155 71.610 ;
        RECT 199.325 71.320 199.575 71.650 ;
        RECT 199.790 71.320 200.470 71.650 ;
        RECT 200.640 71.750 201.715 71.920 ;
        RECT 202.160 71.780 202.720 71.950 ;
        RECT 203.025 71.830 203.485 72.120 ;
        RECT 203.655 72.040 204.875 72.210 ;
        RECT 200.640 71.410 200.810 71.750 ;
        RECT 201.045 71.150 201.375 71.580 ;
        RECT 201.545 71.410 201.715 71.750 ;
        RECT 202.010 71.150 202.380 71.610 ;
        RECT 202.550 71.320 202.720 71.780 ;
        RECT 203.655 71.660 203.825 72.040 ;
        RECT 205.045 71.870 205.215 72.460 ;
        RECT 205.955 72.340 206.165 72.990 ;
        RECT 206.345 72.385 206.660 73.020 ;
        RECT 202.955 71.320 203.825 71.660 ;
        RECT 204.415 71.700 205.215 71.870 ;
        RECT 203.995 71.150 204.245 71.610 ;
        RECT 204.415 71.410 204.585 71.700 ;
        RECT 204.765 71.150 205.095 71.530 ;
        RECT 205.435 71.150 205.740 72.290 ;
        RECT 205.910 71.460 206.165 72.340 ;
        RECT 206.350 71.150 206.660 72.215 ;
        RECT 206.830 72.000 207.040 73.190 ;
        RECT 207.210 73.070 207.540 73.360 ;
        RECT 207.780 73.240 207.950 73.700 ;
        RECT 208.180 73.070 208.510 73.530 ;
        RECT 208.690 73.240 208.860 73.700 ;
        RECT 209.040 73.070 209.370 73.530 ;
        RECT 207.210 72.900 209.370 73.070 ;
        RECT 209.560 72.930 213.070 73.700 ;
        RECT 213.700 72.975 213.990 73.700 ;
        RECT 214.165 73.150 214.420 73.440 ;
        RECT 214.590 73.320 214.920 73.700 ;
        RECT 214.165 72.980 214.915 73.150 ;
        RECT 207.380 72.340 207.875 72.710 ;
        RECT 208.055 72.510 208.855 72.710 ;
        RECT 209.025 72.340 209.355 72.730 ;
        RECT 209.560 72.410 211.210 72.930 ;
        RECT 207.380 72.170 209.355 72.340 ;
        RECT 211.380 72.240 213.070 72.760 ;
        RECT 206.830 71.820 208.480 72.000 ;
        RECT 206.830 71.320 207.065 71.820 ;
        RECT 208.180 71.660 208.480 71.820 ;
        RECT 207.235 71.150 207.565 71.610 ;
        RECT 207.760 71.490 207.950 71.650 ;
        RECT 208.650 71.490 208.870 72.000 ;
        RECT 207.760 71.320 208.870 71.490 ;
        RECT 209.040 71.150 209.370 72.000 ;
        RECT 209.560 71.150 213.070 72.240 ;
        RECT 213.700 71.150 213.990 72.315 ;
        RECT 214.165 72.160 214.515 72.810 ;
        RECT 214.685 71.990 214.915 72.980 ;
        RECT 214.165 71.820 214.915 71.990 ;
        RECT 214.165 71.320 214.420 71.820 ;
        RECT 214.590 71.150 214.920 71.650 ;
        RECT 215.090 71.320 215.260 73.440 ;
        RECT 215.620 73.340 215.950 73.700 ;
        RECT 216.120 73.310 216.615 73.480 ;
        RECT 216.820 73.310 217.675 73.480 ;
        RECT 215.490 72.120 215.950 73.170 ;
        RECT 215.430 71.335 215.755 72.120 ;
        RECT 216.120 71.950 216.290 73.310 ;
        RECT 216.460 72.400 216.810 73.020 ;
        RECT 216.980 72.800 217.335 73.020 ;
        RECT 216.980 72.210 217.150 72.800 ;
        RECT 217.505 72.600 217.675 73.310 ;
        RECT 218.550 73.240 218.880 73.700 ;
        RECT 219.090 73.340 219.440 73.510 ;
        RECT 217.880 72.770 218.670 73.020 ;
        RECT 219.090 72.950 219.350 73.340 ;
        RECT 219.660 73.250 220.610 73.530 ;
        RECT 220.780 73.260 220.970 73.700 ;
        RECT 221.140 73.320 222.210 73.490 ;
        RECT 218.840 72.600 219.010 72.780 ;
        RECT 216.120 71.780 216.515 71.950 ;
        RECT 216.685 71.820 217.150 72.210 ;
        RECT 217.320 72.430 219.010 72.600 ;
        RECT 216.345 71.650 216.515 71.780 ;
        RECT 217.320 71.650 217.490 72.430 ;
        RECT 219.180 72.260 219.350 72.950 ;
        RECT 217.850 72.090 219.350 72.260 ;
        RECT 219.540 72.290 219.750 73.080 ;
        RECT 219.920 72.460 220.270 73.080 ;
        RECT 220.440 72.470 220.610 73.250 ;
        RECT 221.140 73.090 221.310 73.320 ;
        RECT 220.780 72.920 221.310 73.090 ;
        RECT 220.780 72.640 221.000 72.920 ;
        RECT 221.480 72.750 221.720 73.150 ;
        RECT 220.440 72.300 220.845 72.470 ;
        RECT 221.180 72.380 221.720 72.750 ;
        RECT 221.890 72.965 222.210 73.320 ;
        RECT 222.455 73.240 222.760 73.700 ;
        RECT 222.930 72.990 223.185 73.520 ;
        RECT 223.360 73.155 228.705 73.700 ;
        RECT 221.890 72.790 222.215 72.965 ;
        RECT 221.890 72.490 222.805 72.790 ;
        RECT 222.065 72.460 222.805 72.490 ;
        RECT 219.540 72.130 220.215 72.290 ;
        RECT 220.675 72.210 220.845 72.300 ;
        RECT 219.540 72.120 220.505 72.130 ;
        RECT 219.180 71.950 219.350 72.090 ;
        RECT 215.925 71.150 216.175 71.610 ;
        RECT 216.345 71.320 216.595 71.650 ;
        RECT 216.810 71.320 217.490 71.650 ;
        RECT 217.660 71.750 218.735 71.920 ;
        RECT 219.180 71.780 219.740 71.950 ;
        RECT 220.045 71.830 220.505 72.120 ;
        RECT 220.675 72.040 221.895 72.210 ;
        RECT 217.660 71.410 217.830 71.750 ;
        RECT 218.065 71.150 218.395 71.580 ;
        RECT 218.565 71.410 218.735 71.750 ;
        RECT 219.030 71.150 219.400 71.610 ;
        RECT 219.570 71.320 219.740 71.780 ;
        RECT 220.675 71.660 220.845 72.040 ;
        RECT 222.065 71.870 222.235 72.460 ;
        RECT 222.975 72.340 223.185 72.990 ;
        RECT 219.975 71.320 220.845 71.660 ;
        RECT 221.435 71.700 222.235 71.870 ;
        RECT 221.015 71.150 221.265 71.610 ;
        RECT 221.435 71.410 221.605 71.700 ;
        RECT 221.785 71.150 222.115 71.530 ;
        RECT 222.455 71.150 222.760 72.290 ;
        RECT 222.930 71.460 223.185 72.340 ;
        RECT 224.945 72.325 225.285 73.155 ;
        RECT 229.805 72.935 230.260 73.700 ;
        RECT 230.535 73.320 231.835 73.530 ;
        RECT 232.090 73.340 232.420 73.700 ;
        RECT 231.665 73.170 231.835 73.320 ;
        RECT 232.590 73.200 232.850 73.530 ;
        RECT 232.620 73.190 232.850 73.200 ;
        RECT 226.765 71.585 227.115 72.835 ;
        RECT 230.735 72.710 230.955 73.110 ;
        RECT 229.800 72.510 230.290 72.710 ;
        RECT 230.480 72.500 230.955 72.710 ;
        RECT 231.200 72.710 231.410 73.110 ;
        RECT 231.665 73.045 232.420 73.170 ;
        RECT 231.665 73.000 232.510 73.045 ;
        RECT 232.240 72.880 232.510 73.000 ;
        RECT 231.200 72.500 231.530 72.710 ;
        RECT 231.700 72.440 232.110 72.745 ;
        RECT 229.805 72.270 230.980 72.330 ;
        RECT 232.340 72.305 232.510 72.880 ;
        RECT 232.310 72.270 232.510 72.305 ;
        RECT 229.805 72.160 232.510 72.270 ;
        RECT 223.360 71.150 228.705 71.585 ;
        RECT 229.805 71.540 230.060 72.160 ;
        RECT 230.650 72.100 232.450 72.160 ;
        RECT 230.650 72.070 230.980 72.100 ;
        RECT 232.680 72.000 232.850 73.190 ;
        RECT 233.020 72.930 235.610 73.700 ;
        RECT 235.870 73.050 236.040 73.530 ;
        RECT 236.210 73.220 236.540 73.700 ;
        RECT 236.765 73.280 238.300 73.530 ;
        RECT 236.765 73.050 236.935 73.280 ;
        RECT 233.020 72.410 234.230 72.930 ;
        RECT 235.870 72.880 236.935 73.050 ;
        RECT 234.400 72.240 235.610 72.760 ;
        RECT 237.115 72.710 237.395 73.110 ;
        RECT 235.785 72.500 236.135 72.710 ;
        RECT 236.305 72.510 236.750 72.710 ;
        RECT 236.920 72.510 237.395 72.710 ;
        RECT 237.665 72.710 237.950 73.110 ;
        RECT 238.130 73.050 238.300 73.280 ;
        RECT 238.470 73.220 238.800 73.700 ;
        RECT 239.015 73.200 239.270 73.530 ;
        RECT 239.060 73.190 239.270 73.200 ;
        RECT 239.085 73.120 239.270 73.190 ;
        RECT 238.130 72.880 238.930 73.050 ;
        RECT 237.665 72.510 237.995 72.710 ;
        RECT 238.165 72.680 238.530 72.710 ;
        RECT 238.165 72.510 238.540 72.680 ;
        RECT 238.760 72.330 238.930 72.880 ;
        RECT 230.310 71.900 230.495 71.990 ;
        RECT 231.085 71.900 231.920 71.910 ;
        RECT 230.310 71.700 231.920 71.900 ;
        RECT 230.310 71.660 230.540 71.700 ;
        RECT 229.805 71.320 230.140 71.540 ;
        RECT 231.145 71.150 231.500 71.530 ;
        RECT 231.670 71.320 231.920 71.700 ;
        RECT 232.170 71.150 232.420 71.930 ;
        RECT 232.590 71.320 232.850 72.000 ;
        RECT 233.020 71.150 235.610 72.240 ;
        RECT 235.870 72.160 238.930 72.330 ;
        RECT 235.870 71.320 236.040 72.160 ;
        RECT 239.100 71.990 239.270 73.120 ;
        RECT 239.460 72.975 239.750 73.700 ;
        RECT 239.920 72.950 241.130 73.700 ;
        RECT 241.320 73.200 241.575 73.530 ;
        RECT 241.790 73.220 242.120 73.700 ;
        RECT 242.290 73.280 243.825 73.530 ;
        RECT 241.320 73.190 241.530 73.200 ;
        RECT 241.320 73.120 241.505 73.190 ;
        RECT 239.920 72.410 240.440 72.950 ;
        RECT 236.210 71.490 236.540 71.990 ;
        RECT 236.710 71.750 238.345 71.990 ;
        RECT 236.710 71.660 236.940 71.750 ;
        RECT 237.050 71.490 237.380 71.530 ;
        RECT 236.210 71.320 237.380 71.490 ;
        RECT 237.570 71.150 237.925 71.570 ;
        RECT 238.095 71.320 238.345 71.750 ;
        RECT 238.515 71.150 238.845 71.910 ;
        RECT 239.015 71.320 239.270 71.990 ;
        RECT 239.460 71.150 239.750 72.315 ;
        RECT 240.610 72.240 241.130 72.780 ;
        RECT 239.920 71.150 241.130 72.240 ;
        RECT 241.320 71.990 241.490 73.120 ;
        RECT 242.290 73.050 242.460 73.280 ;
        RECT 241.660 72.880 242.460 73.050 ;
        RECT 241.660 72.330 241.830 72.880 ;
        RECT 242.640 72.710 242.925 73.110 ;
        RECT 242.060 72.510 242.425 72.710 ;
        RECT 242.595 72.510 242.925 72.710 ;
        RECT 243.195 72.710 243.475 73.110 ;
        RECT 243.655 73.050 243.825 73.280 ;
        RECT 244.050 73.220 244.380 73.700 ;
        RECT 244.550 73.050 244.720 73.530 ;
        RECT 244.980 73.155 250.325 73.700 ;
        RECT 250.500 73.155 255.845 73.700 ;
        RECT 243.655 72.880 244.720 73.050 ;
        RECT 243.195 72.510 243.670 72.710 ;
        RECT 243.840 72.510 244.285 72.710 ;
        RECT 244.455 72.500 244.805 72.710 ;
        RECT 241.660 72.160 244.720 72.330 ;
        RECT 246.565 72.325 246.905 73.155 ;
        RECT 241.320 71.320 241.575 71.990 ;
        RECT 241.745 71.150 242.075 71.910 ;
        RECT 242.245 71.750 243.880 71.990 ;
        RECT 242.245 71.320 242.495 71.750 ;
        RECT 243.650 71.660 243.880 71.750 ;
        RECT 242.665 71.150 243.020 71.570 ;
        RECT 243.210 71.490 243.540 71.530 ;
        RECT 244.050 71.490 244.380 71.990 ;
        RECT 243.210 71.320 244.380 71.490 ;
        RECT 244.550 71.320 244.720 72.160 ;
        RECT 248.385 71.585 248.735 72.835 ;
        RECT 252.085 72.325 252.425 73.155 ;
        RECT 256.020 72.930 257.690 73.700 ;
        RECT 258.325 72.935 258.780 73.700 ;
        RECT 259.055 73.320 260.355 73.530 ;
        RECT 260.610 73.340 260.940 73.700 ;
        RECT 260.185 73.170 260.355 73.320 ;
        RECT 261.110 73.200 261.370 73.530 ;
        RECT 253.905 71.585 254.255 72.835 ;
        RECT 256.020 72.410 256.770 72.930 ;
        RECT 256.940 72.240 257.690 72.760 ;
        RECT 259.255 72.710 259.475 73.110 ;
        RECT 258.320 72.510 258.810 72.710 ;
        RECT 259.000 72.500 259.475 72.710 ;
        RECT 259.720 72.710 259.930 73.110 ;
        RECT 260.185 73.045 260.940 73.170 ;
        RECT 260.185 73.000 261.030 73.045 ;
        RECT 260.760 72.880 261.030 73.000 ;
        RECT 259.720 72.500 260.050 72.710 ;
        RECT 260.220 72.440 260.630 72.745 ;
        RECT 244.980 71.150 250.325 71.585 ;
        RECT 250.500 71.150 255.845 71.585 ;
        RECT 256.020 71.150 257.690 72.240 ;
        RECT 258.325 72.270 259.500 72.330 ;
        RECT 260.860 72.305 261.030 72.880 ;
        RECT 260.830 72.270 261.030 72.305 ;
        RECT 258.325 72.160 261.030 72.270 ;
        RECT 258.325 71.540 258.580 72.160 ;
        RECT 259.170 72.100 260.970 72.160 ;
        RECT 259.170 72.070 259.500 72.100 ;
        RECT 261.200 72.000 261.370 73.200 ;
        RECT 258.830 71.900 259.015 71.990 ;
        RECT 259.605 71.900 260.440 71.910 ;
        RECT 258.830 71.700 260.440 71.900 ;
        RECT 258.830 71.660 259.060 71.700 ;
        RECT 258.325 71.320 258.660 71.540 ;
        RECT 259.665 71.150 260.020 71.530 ;
        RECT 260.190 71.320 260.440 71.700 ;
        RECT 260.690 71.150 260.940 71.930 ;
        RECT 261.110 71.320 261.370 72.000 ;
        RECT 261.540 73.200 261.800 73.530 ;
        RECT 261.970 73.340 262.300 73.700 ;
        RECT 262.555 73.320 263.855 73.530 ;
        RECT 261.540 72.000 261.710 73.200 ;
        RECT 262.555 73.170 262.725 73.320 ;
        RECT 261.970 73.045 262.725 73.170 ;
        RECT 261.880 73.000 262.725 73.045 ;
        RECT 261.880 72.880 262.150 73.000 ;
        RECT 261.880 72.305 262.050 72.880 ;
        RECT 262.280 72.440 262.690 72.745 ;
        RECT 262.980 72.710 263.190 73.110 ;
        RECT 262.860 72.500 263.190 72.710 ;
        RECT 263.435 72.710 263.655 73.110 ;
        RECT 264.130 72.935 264.585 73.700 ;
        RECT 265.220 72.975 265.510 73.700 ;
        RECT 265.680 73.155 271.025 73.700 ;
        RECT 263.435 72.500 263.910 72.710 ;
        RECT 264.100 72.510 264.590 72.710 ;
        RECT 261.880 72.270 262.080 72.305 ;
        RECT 263.410 72.270 264.585 72.330 ;
        RECT 267.265 72.325 267.605 73.155 ;
        RECT 271.200 72.930 273.790 73.700 ;
        RECT 274.440 73.070 274.770 73.530 ;
        RECT 274.950 73.240 275.120 73.700 ;
        RECT 275.300 73.070 275.630 73.530 ;
        RECT 275.860 73.240 276.030 73.700 ;
        RECT 276.270 73.360 277.460 73.530 ;
        RECT 276.270 73.070 276.600 73.360 ;
        RECT 277.150 73.190 277.460 73.360 ;
        RECT 261.880 72.160 264.585 72.270 ;
        RECT 261.940 72.100 263.740 72.160 ;
        RECT 263.410 72.070 263.740 72.100 ;
        RECT 261.540 71.320 261.800 72.000 ;
        RECT 261.970 71.150 262.220 71.930 ;
        RECT 262.470 71.900 263.305 71.910 ;
        RECT 263.895 71.900 264.080 71.990 ;
        RECT 262.470 71.700 264.080 71.900 ;
        RECT 262.470 71.320 262.720 71.700 ;
        RECT 263.850 71.660 264.080 71.700 ;
        RECT 264.330 71.540 264.585 72.160 ;
        RECT 262.890 71.150 263.245 71.530 ;
        RECT 264.250 71.320 264.585 71.540 ;
        RECT 265.220 71.150 265.510 72.315 ;
        RECT 269.085 71.585 269.435 72.835 ;
        RECT 271.200 72.410 272.410 72.930 ;
        RECT 274.440 72.900 276.600 73.070 ;
        RECT 272.580 72.240 273.790 72.760 ;
        RECT 265.680 71.150 271.025 71.585 ;
        RECT 271.200 71.150 273.790 72.240 ;
        RECT 274.455 72.340 274.785 72.730 ;
        RECT 274.955 72.510 275.755 72.710 ;
        RECT 275.935 72.340 276.430 72.710 ;
        RECT 274.455 72.170 276.430 72.340 ;
        RECT 276.770 72.000 276.980 73.190 ;
        RECT 277.150 72.385 277.465 73.020 ;
        RECT 277.645 72.990 277.900 73.520 ;
        RECT 278.070 73.240 278.375 73.700 ;
        RECT 278.620 73.320 279.690 73.490 ;
        RECT 277.645 72.340 277.855 72.990 ;
        RECT 278.620 72.965 278.940 73.320 ;
        RECT 278.615 72.790 278.940 72.965 ;
        RECT 278.025 72.490 278.940 72.790 ;
        RECT 279.110 72.750 279.350 73.150 ;
        RECT 279.520 73.090 279.690 73.320 ;
        RECT 279.860 73.260 280.050 73.700 ;
        RECT 280.220 73.250 281.170 73.530 ;
        RECT 281.390 73.340 281.740 73.510 ;
        RECT 279.520 72.920 280.050 73.090 ;
        RECT 278.025 72.460 278.765 72.490 ;
        RECT 274.440 71.150 274.770 72.000 ;
        RECT 274.940 71.490 275.160 72.000 ;
        RECT 275.330 71.820 276.980 72.000 ;
        RECT 275.330 71.660 275.630 71.820 ;
        RECT 275.860 71.490 276.050 71.650 ;
        RECT 274.940 71.320 276.050 71.490 ;
        RECT 276.245 71.150 276.575 71.610 ;
        RECT 276.745 71.320 276.980 71.820 ;
        RECT 277.150 71.150 277.460 72.215 ;
        RECT 277.645 71.460 277.900 72.340 ;
        RECT 278.070 71.150 278.375 72.290 ;
        RECT 278.595 71.870 278.765 72.460 ;
        RECT 279.110 72.380 279.650 72.750 ;
        RECT 279.830 72.640 280.050 72.920 ;
        RECT 280.220 72.470 280.390 73.250 ;
        RECT 279.985 72.300 280.390 72.470 ;
        RECT 280.560 72.460 280.910 73.080 ;
        RECT 279.985 72.210 280.155 72.300 ;
        RECT 281.080 72.290 281.290 73.080 ;
        RECT 278.935 72.040 280.155 72.210 ;
        RECT 280.615 72.130 281.290 72.290 ;
        RECT 278.595 71.700 279.395 71.870 ;
        RECT 278.715 71.150 279.045 71.530 ;
        RECT 279.225 71.410 279.395 71.700 ;
        RECT 279.985 71.660 280.155 72.040 ;
        RECT 280.325 72.120 281.290 72.130 ;
        RECT 281.480 72.950 281.740 73.340 ;
        RECT 281.950 73.240 282.280 73.700 ;
        RECT 283.155 73.310 284.010 73.480 ;
        RECT 284.215 73.310 284.710 73.480 ;
        RECT 284.880 73.340 285.210 73.700 ;
        RECT 281.480 72.260 281.650 72.950 ;
        RECT 281.820 72.600 281.990 72.780 ;
        RECT 282.160 72.770 282.950 73.020 ;
        RECT 283.155 72.600 283.325 73.310 ;
        RECT 283.495 72.800 283.850 73.020 ;
        RECT 281.820 72.430 283.510 72.600 ;
        RECT 280.325 71.830 280.785 72.120 ;
        RECT 281.480 72.090 282.980 72.260 ;
        RECT 281.480 71.950 281.650 72.090 ;
        RECT 281.090 71.780 281.650 71.950 ;
        RECT 279.565 71.150 279.815 71.610 ;
        RECT 279.985 71.320 280.855 71.660 ;
        RECT 281.090 71.320 281.260 71.780 ;
        RECT 282.095 71.750 283.170 71.920 ;
        RECT 281.430 71.150 281.800 71.610 ;
        RECT 282.095 71.410 282.265 71.750 ;
        RECT 282.435 71.150 282.765 71.580 ;
        RECT 283.000 71.410 283.170 71.750 ;
        RECT 283.340 71.650 283.510 72.430 ;
        RECT 283.680 72.210 283.850 72.800 ;
        RECT 284.020 72.400 284.370 73.020 ;
        RECT 283.680 71.820 284.145 72.210 ;
        RECT 284.540 71.950 284.710 73.310 ;
        RECT 284.880 72.120 285.340 73.170 ;
        RECT 284.315 71.780 284.710 71.950 ;
        RECT 284.315 71.650 284.485 71.780 ;
        RECT 283.340 71.320 284.020 71.650 ;
        RECT 284.235 71.320 284.485 71.650 ;
        RECT 284.655 71.150 284.905 71.610 ;
        RECT 285.075 71.335 285.400 72.120 ;
        RECT 285.570 71.320 285.740 73.440 ;
        RECT 285.910 73.320 286.240 73.700 ;
        RECT 286.410 73.150 286.665 73.440 ;
        RECT 285.915 72.980 286.665 73.150 ;
        RECT 285.915 71.990 286.145 72.980 ;
        RECT 286.845 72.960 287.100 73.530 ;
        RECT 287.270 73.300 287.600 73.700 ;
        RECT 288.025 73.165 288.555 73.530 ;
        RECT 288.025 73.130 288.200 73.165 ;
        RECT 287.270 72.960 288.200 73.130 ;
        RECT 286.315 72.160 286.665 72.810 ;
        RECT 286.845 72.290 287.015 72.960 ;
        RECT 287.270 72.790 287.440 72.960 ;
        RECT 287.185 72.460 287.440 72.790 ;
        RECT 287.665 72.460 287.860 72.790 ;
        RECT 285.915 71.820 286.665 71.990 ;
        RECT 285.910 71.150 286.240 71.650 ;
        RECT 286.410 71.320 286.665 71.820 ;
        RECT 286.845 71.320 287.180 72.290 ;
        RECT 287.350 71.150 287.520 72.290 ;
        RECT 287.690 71.490 287.860 72.460 ;
        RECT 288.030 71.830 288.200 72.960 ;
        RECT 288.370 72.170 288.540 72.970 ;
        RECT 288.745 72.680 289.020 73.530 ;
        RECT 288.740 72.510 289.020 72.680 ;
        RECT 288.745 72.370 289.020 72.510 ;
        RECT 289.190 72.170 289.380 73.530 ;
        RECT 289.560 73.165 290.070 73.700 ;
        RECT 290.290 72.890 290.535 73.495 ;
        RECT 290.980 72.975 291.270 73.700 ;
        RECT 291.440 73.155 296.785 73.700 ;
        RECT 289.580 72.720 290.810 72.890 ;
        RECT 288.370 72.000 289.380 72.170 ;
        RECT 289.550 72.155 290.300 72.345 ;
        RECT 288.030 71.660 289.155 71.830 ;
        RECT 289.550 71.490 289.720 72.155 ;
        RECT 290.470 71.910 290.810 72.720 ;
        RECT 293.025 72.325 293.365 73.155 ;
        RECT 296.965 73.150 297.220 73.440 ;
        RECT 297.390 73.320 297.720 73.700 ;
        RECT 296.965 72.980 297.715 73.150 ;
        RECT 287.690 71.320 289.720 71.490 ;
        RECT 289.890 71.150 290.060 71.910 ;
        RECT 290.295 71.500 290.810 71.910 ;
        RECT 290.980 71.150 291.270 72.315 ;
        RECT 294.845 71.585 295.195 72.835 ;
        RECT 296.965 72.160 297.315 72.810 ;
        RECT 297.485 71.990 297.715 72.980 ;
        RECT 296.965 71.820 297.715 71.990 ;
        RECT 291.440 71.150 296.785 71.585 ;
        RECT 296.965 71.320 297.220 71.820 ;
        RECT 297.390 71.150 297.720 71.650 ;
        RECT 297.890 71.320 298.060 73.440 ;
        RECT 298.420 73.340 298.750 73.700 ;
        RECT 298.920 73.310 299.415 73.480 ;
        RECT 299.620 73.310 300.475 73.480 ;
        RECT 298.290 72.120 298.750 73.170 ;
        RECT 298.230 71.335 298.555 72.120 ;
        RECT 298.920 71.950 299.090 73.310 ;
        RECT 299.260 72.400 299.610 73.020 ;
        RECT 299.780 72.800 300.135 73.020 ;
        RECT 299.780 72.210 299.950 72.800 ;
        RECT 300.305 72.600 300.475 73.310 ;
        RECT 301.350 73.240 301.680 73.700 ;
        RECT 301.890 73.340 302.240 73.510 ;
        RECT 300.680 72.770 301.470 73.020 ;
        RECT 301.890 72.950 302.150 73.340 ;
        RECT 302.460 73.250 303.410 73.530 ;
        RECT 303.580 73.260 303.770 73.700 ;
        RECT 303.940 73.320 305.010 73.490 ;
        RECT 301.640 72.600 301.810 72.780 ;
        RECT 298.920 71.780 299.315 71.950 ;
        RECT 299.485 71.820 299.950 72.210 ;
        RECT 300.120 72.430 301.810 72.600 ;
        RECT 299.145 71.650 299.315 71.780 ;
        RECT 300.120 71.650 300.290 72.430 ;
        RECT 301.980 72.260 302.150 72.950 ;
        RECT 300.650 72.090 302.150 72.260 ;
        RECT 302.340 72.290 302.550 73.080 ;
        RECT 302.720 72.460 303.070 73.080 ;
        RECT 303.240 72.470 303.410 73.250 ;
        RECT 303.940 73.090 304.110 73.320 ;
        RECT 303.580 72.920 304.110 73.090 ;
        RECT 303.580 72.640 303.800 72.920 ;
        RECT 304.280 72.750 304.520 73.150 ;
        RECT 303.240 72.300 303.645 72.470 ;
        RECT 303.980 72.380 304.520 72.750 ;
        RECT 304.690 72.965 305.010 73.320 ;
        RECT 305.255 73.240 305.560 73.700 ;
        RECT 305.730 72.990 305.980 73.520 ;
        RECT 304.690 72.790 305.015 72.965 ;
        RECT 304.690 72.490 305.605 72.790 ;
        RECT 304.865 72.460 305.605 72.490 ;
        RECT 302.340 72.130 303.015 72.290 ;
        RECT 303.475 72.210 303.645 72.300 ;
        RECT 302.340 72.120 303.305 72.130 ;
        RECT 301.980 71.950 302.150 72.090 ;
        RECT 298.725 71.150 298.975 71.610 ;
        RECT 299.145 71.320 299.395 71.650 ;
        RECT 299.610 71.320 300.290 71.650 ;
        RECT 300.460 71.750 301.535 71.920 ;
        RECT 301.980 71.780 302.540 71.950 ;
        RECT 302.845 71.830 303.305 72.120 ;
        RECT 303.475 72.040 304.695 72.210 ;
        RECT 300.460 71.410 300.630 71.750 ;
        RECT 300.865 71.150 301.195 71.580 ;
        RECT 301.365 71.410 301.535 71.750 ;
        RECT 301.830 71.150 302.200 71.610 ;
        RECT 302.370 71.320 302.540 71.780 ;
        RECT 303.475 71.660 303.645 72.040 ;
        RECT 304.865 71.870 305.035 72.460 ;
        RECT 305.775 72.340 305.980 72.990 ;
        RECT 306.150 72.945 306.400 73.700 ;
        RECT 307.170 73.150 307.340 73.530 ;
        RECT 307.555 73.320 307.885 73.700 ;
        RECT 307.170 72.980 307.885 73.150 ;
        RECT 307.080 72.430 307.435 72.800 ;
        RECT 307.715 72.790 307.885 72.980 ;
        RECT 308.055 72.955 308.310 73.530 ;
        RECT 307.715 72.460 307.970 72.790 ;
        RECT 302.775 71.320 303.645 71.660 ;
        RECT 304.235 71.700 305.035 71.870 ;
        RECT 303.815 71.150 304.065 71.610 ;
        RECT 304.235 71.410 304.405 71.700 ;
        RECT 304.585 71.150 304.915 71.530 ;
        RECT 305.255 71.150 305.560 72.290 ;
        RECT 305.730 71.460 305.980 72.340 ;
        RECT 306.150 71.150 306.400 72.290 ;
        RECT 307.715 72.250 307.885 72.460 ;
        RECT 307.170 72.080 307.885 72.250 ;
        RECT 308.140 72.225 308.310 72.955 ;
        RECT 308.485 72.860 308.745 73.700 ;
        RECT 309.840 72.950 311.050 73.700 ;
        RECT 307.170 71.320 307.340 72.080 ;
        RECT 307.555 71.150 307.885 71.910 ;
        RECT 308.055 71.320 308.310 72.225 ;
        RECT 308.485 71.150 308.745 72.300 ;
        RECT 309.840 72.240 310.360 72.780 ;
        RECT 310.530 72.410 311.050 72.950 ;
        RECT 309.840 71.150 311.050 72.240 ;
        RECT 162.095 70.980 311.135 71.150 ;
        RECT 162.180 69.890 163.390 70.980 ;
        RECT 163.560 70.545 168.905 70.980 ;
        RECT 162.180 69.180 162.700 69.720 ;
        RECT 162.870 69.350 163.390 69.890 ;
        RECT 162.180 68.430 163.390 69.180 ;
        RECT 165.145 68.975 165.485 69.805 ;
        RECT 166.965 69.295 167.315 70.545 ;
        RECT 169.080 69.890 170.750 70.980 ;
        RECT 169.080 69.200 169.830 69.720 ;
        RECT 170.000 69.370 170.750 69.890 ;
        RECT 170.925 69.840 171.260 70.810 ;
        RECT 171.430 69.840 171.600 70.980 ;
        RECT 171.770 70.640 173.800 70.810 ;
        RECT 163.560 68.430 168.905 68.975 ;
        RECT 169.080 68.430 170.750 69.200 ;
        RECT 170.925 69.170 171.095 69.840 ;
        RECT 171.770 69.670 171.940 70.640 ;
        RECT 171.265 69.340 171.520 69.670 ;
        RECT 171.745 69.340 171.940 69.670 ;
        RECT 172.110 70.300 173.235 70.470 ;
        RECT 171.350 69.170 171.520 69.340 ;
        RECT 172.110 69.170 172.280 70.300 ;
        RECT 170.925 68.600 171.180 69.170 ;
        RECT 171.350 69.000 172.280 69.170 ;
        RECT 172.450 69.960 173.460 70.130 ;
        RECT 172.450 69.160 172.620 69.960 ;
        RECT 172.825 69.620 173.100 69.760 ;
        RECT 172.820 69.450 173.100 69.620 ;
        RECT 172.105 68.965 172.280 69.000 ;
        RECT 171.350 68.430 171.680 68.830 ;
        RECT 172.105 68.600 172.635 68.965 ;
        RECT 172.825 68.600 173.100 69.450 ;
        RECT 173.270 68.600 173.460 69.960 ;
        RECT 173.630 69.975 173.800 70.640 ;
        RECT 173.970 70.220 174.140 70.980 ;
        RECT 174.375 70.220 174.890 70.630 ;
        RECT 173.630 69.785 174.380 69.975 ;
        RECT 174.550 69.410 174.890 70.220 ;
        RECT 175.060 69.815 175.350 70.980 ;
        RECT 175.525 69.840 175.860 70.810 ;
        RECT 176.030 69.840 176.200 70.980 ;
        RECT 176.370 70.640 178.400 70.810 ;
        RECT 173.660 69.240 174.890 69.410 ;
        RECT 173.640 68.430 174.150 68.965 ;
        RECT 174.370 68.635 174.615 69.240 ;
        RECT 175.525 69.170 175.695 69.840 ;
        RECT 176.370 69.670 176.540 70.640 ;
        RECT 175.865 69.340 176.120 69.670 ;
        RECT 176.345 69.340 176.540 69.670 ;
        RECT 176.710 70.300 177.835 70.470 ;
        RECT 175.950 69.170 176.120 69.340 ;
        RECT 176.710 69.170 176.880 70.300 ;
        RECT 175.060 68.430 175.350 69.155 ;
        RECT 175.525 68.600 175.780 69.170 ;
        RECT 175.950 69.000 176.880 69.170 ;
        RECT 177.050 69.960 178.060 70.130 ;
        RECT 177.050 69.160 177.220 69.960 ;
        RECT 176.705 68.965 176.880 69.000 ;
        RECT 175.950 68.430 176.280 68.830 ;
        RECT 176.705 68.600 177.235 68.965 ;
        RECT 177.425 68.940 177.700 69.760 ;
        RECT 177.420 68.770 177.700 68.940 ;
        RECT 177.425 68.600 177.700 68.770 ;
        RECT 177.870 68.600 178.060 69.960 ;
        RECT 178.230 69.975 178.400 70.640 ;
        RECT 178.570 70.220 178.740 70.980 ;
        RECT 178.975 70.220 179.490 70.630 ;
        RECT 178.230 69.785 178.980 69.975 ;
        RECT 179.150 69.410 179.490 70.220 ;
        RECT 179.660 69.890 183.170 70.980 ;
        RECT 178.260 69.240 179.490 69.410 ;
        RECT 178.240 68.430 178.750 68.965 ;
        RECT 178.970 68.635 179.215 69.240 ;
        RECT 179.660 69.200 181.310 69.720 ;
        RECT 181.480 69.370 183.170 69.890 ;
        RECT 183.390 69.885 183.640 70.980 ;
        RECT 184.375 70.640 186.440 70.810 ;
        RECT 183.810 69.800 184.165 70.215 ;
        RECT 184.375 69.800 184.620 70.640 ;
        RECT 183.995 69.630 184.165 69.800 ;
        RECT 183.340 69.420 183.825 69.630 ;
        RECT 183.995 69.420 184.620 69.630 ;
        RECT 183.995 69.250 184.165 69.420 ;
        RECT 184.790 69.250 185.040 70.470 ;
        RECT 185.210 69.800 185.480 70.640 ;
        RECT 185.770 69.970 186.020 70.470 ;
        RECT 186.190 70.140 186.440 70.640 ;
        RECT 186.610 69.970 186.860 70.810 ;
        RECT 187.030 70.140 187.280 70.980 ;
        RECT 187.450 69.970 187.765 70.810 ;
        RECT 188.190 70.250 188.485 70.980 ;
        RECT 188.655 70.080 188.915 70.805 ;
        RECT 189.085 70.250 189.345 70.980 ;
        RECT 189.515 70.080 189.775 70.805 ;
        RECT 189.945 70.250 190.205 70.980 ;
        RECT 190.375 70.080 190.635 70.805 ;
        RECT 190.805 70.250 191.065 70.980 ;
        RECT 191.235 70.080 191.495 70.805 ;
        RECT 185.770 69.800 187.765 69.970 ;
        RECT 188.185 69.840 191.495 70.080 ;
        RECT 191.665 69.870 191.925 70.980 ;
        RECT 185.215 69.420 186.720 69.630 ;
        RECT 186.890 69.420 187.745 69.630 ;
        RECT 188.185 69.250 189.155 69.840 ;
        RECT 192.095 69.670 192.345 70.805 ;
        RECT 192.525 69.870 192.820 70.980 ;
        RECT 193.970 69.885 194.220 70.980 ;
        RECT 194.955 70.640 197.020 70.810 ;
        RECT 194.390 69.800 194.745 70.215 ;
        RECT 194.955 69.800 195.200 70.640 ;
        RECT 189.325 69.420 192.345 69.670 ;
        RECT 179.660 68.430 183.170 69.200 ;
        RECT 183.350 68.430 183.640 69.170 ;
        RECT 183.810 68.725 184.165 69.250 ;
        RECT 184.375 68.430 184.580 69.240 ;
        RECT 184.750 69.070 187.320 69.250 ;
        RECT 184.750 68.600 185.080 69.070 ;
        RECT 185.250 68.430 185.980 68.900 ;
        RECT 186.150 68.600 186.480 69.070 ;
        RECT 186.650 68.430 186.820 68.900 ;
        RECT 186.990 68.600 187.320 69.070 ;
        RECT 187.490 68.430 187.765 69.250 ;
        RECT 188.185 69.080 191.495 69.250 ;
        RECT 188.185 68.430 188.485 68.910 ;
        RECT 188.655 68.625 188.915 69.080 ;
        RECT 189.085 68.430 189.345 68.910 ;
        RECT 189.515 68.625 189.775 69.080 ;
        RECT 189.945 68.430 190.205 68.910 ;
        RECT 190.375 68.625 190.635 69.080 ;
        RECT 190.805 68.430 191.065 68.910 ;
        RECT 191.235 68.625 191.495 69.080 ;
        RECT 191.665 68.430 191.925 68.955 ;
        RECT 192.095 68.610 192.345 69.420 ;
        RECT 192.515 69.060 192.830 69.670 ;
        RECT 194.575 69.630 194.745 69.800 ;
        RECT 193.920 69.420 194.405 69.630 ;
        RECT 194.575 69.420 195.200 69.630 ;
        RECT 194.575 69.250 194.745 69.420 ;
        RECT 195.370 69.250 195.620 70.470 ;
        RECT 195.790 69.800 196.060 70.640 ;
        RECT 196.350 69.970 196.600 70.470 ;
        RECT 196.770 70.140 197.020 70.640 ;
        RECT 197.190 69.970 197.440 70.810 ;
        RECT 197.610 70.140 197.860 70.980 ;
        RECT 198.030 69.970 198.345 70.810 ;
        RECT 196.350 69.800 198.345 69.970 ;
        RECT 198.520 69.890 200.190 70.980 ;
        RECT 195.795 69.420 197.300 69.630 ;
        RECT 197.470 69.420 198.325 69.630 ;
        RECT 192.525 68.430 192.770 68.890 ;
        RECT 193.930 68.430 194.220 69.170 ;
        RECT 194.390 68.725 194.745 69.250 ;
        RECT 194.955 68.430 195.160 69.240 ;
        RECT 195.330 69.070 197.900 69.250 ;
        RECT 195.330 68.600 195.660 69.070 ;
        RECT 195.830 68.430 196.560 68.900 ;
        RECT 196.730 68.600 197.060 69.070 ;
        RECT 197.230 68.430 197.400 68.900 ;
        RECT 197.570 68.600 197.900 69.070 ;
        RECT 198.070 68.430 198.345 69.250 ;
        RECT 198.520 69.200 199.270 69.720 ;
        RECT 199.440 69.370 200.190 69.890 ;
        RECT 200.820 69.815 201.110 70.980 ;
        RECT 201.285 69.840 201.620 70.810 ;
        RECT 201.790 69.840 201.960 70.980 ;
        RECT 202.130 70.640 204.160 70.810 ;
        RECT 198.520 68.430 200.190 69.200 ;
        RECT 201.285 69.170 201.455 69.840 ;
        RECT 202.130 69.670 202.300 70.640 ;
        RECT 201.625 69.340 201.880 69.670 ;
        RECT 202.105 69.340 202.300 69.670 ;
        RECT 202.470 70.300 203.595 70.470 ;
        RECT 201.710 69.170 201.880 69.340 ;
        RECT 202.470 69.170 202.640 70.300 ;
        RECT 200.820 68.430 201.110 69.155 ;
        RECT 201.285 68.600 201.540 69.170 ;
        RECT 201.710 69.000 202.640 69.170 ;
        RECT 202.810 69.960 203.820 70.130 ;
        RECT 202.810 69.160 202.980 69.960 ;
        RECT 202.465 68.965 202.640 69.000 ;
        RECT 201.710 68.430 202.040 68.830 ;
        RECT 202.465 68.600 202.995 68.965 ;
        RECT 203.185 68.940 203.460 69.760 ;
        RECT 203.180 68.770 203.460 68.940 ;
        RECT 203.185 68.600 203.460 68.770 ;
        RECT 203.630 68.600 203.820 69.960 ;
        RECT 203.990 69.975 204.160 70.640 ;
        RECT 204.330 70.220 204.500 70.980 ;
        RECT 204.735 70.220 205.250 70.630 ;
        RECT 205.420 70.545 210.765 70.980 ;
        RECT 203.990 69.785 204.740 69.975 ;
        RECT 204.910 69.410 205.250 70.220 ;
        RECT 204.020 69.240 205.250 69.410 ;
        RECT 204.000 68.430 204.510 68.965 ;
        RECT 204.730 68.635 204.975 69.240 ;
        RECT 207.005 68.975 207.345 69.805 ;
        RECT 208.825 69.295 209.175 70.545 ;
        RECT 212.065 70.010 212.395 70.810 ;
        RECT 212.565 70.180 212.895 70.980 ;
        RECT 213.195 70.010 213.525 70.810 ;
        RECT 214.170 70.180 214.420 70.980 ;
        RECT 212.065 69.840 214.500 70.010 ;
        RECT 214.690 69.840 214.860 70.980 ;
        RECT 215.030 69.840 215.370 70.810 ;
        RECT 215.540 70.545 220.885 70.980 ;
        RECT 221.060 70.545 226.405 70.980 ;
        RECT 211.860 69.420 212.210 69.670 ;
        RECT 212.395 69.210 212.565 69.840 ;
        RECT 212.735 69.420 213.065 69.620 ;
        RECT 213.235 69.420 213.565 69.620 ;
        RECT 213.735 69.420 214.155 69.620 ;
        RECT 214.330 69.590 214.500 69.840 ;
        RECT 215.140 69.790 215.370 69.840 ;
        RECT 214.330 69.420 215.025 69.590 ;
        RECT 205.420 68.430 210.765 68.975 ;
        RECT 212.065 68.600 212.565 69.210 ;
        RECT 213.195 69.080 214.420 69.250 ;
        RECT 215.195 69.230 215.370 69.790 ;
        RECT 213.195 68.600 213.525 69.080 ;
        RECT 213.695 68.430 213.920 68.890 ;
        RECT 214.090 68.600 214.420 69.080 ;
        RECT 214.610 68.430 214.860 69.230 ;
        RECT 215.030 68.600 215.370 69.230 ;
        RECT 217.125 68.975 217.465 69.805 ;
        RECT 218.945 69.295 219.295 70.545 ;
        RECT 222.645 68.975 222.985 69.805 ;
        RECT 224.465 69.295 224.815 70.545 ;
        RECT 226.580 69.815 226.870 70.980 ;
        RECT 227.040 70.545 232.385 70.980 ;
        RECT 233.480 70.550 233.820 70.810 ;
        RECT 215.540 68.430 220.885 68.975 ;
        RECT 221.060 68.430 226.405 68.975 ;
        RECT 226.580 68.430 226.870 69.155 ;
        RECT 228.625 68.975 228.965 69.805 ;
        RECT 230.445 69.295 230.795 70.545 ;
        RECT 233.480 69.150 233.740 70.550 ;
        RECT 233.990 70.180 234.320 70.980 ;
        RECT 234.785 70.010 235.035 70.810 ;
        RECT 235.220 70.260 235.550 70.980 ;
        RECT 235.770 70.010 236.020 70.810 ;
        RECT 236.190 70.600 236.525 70.980 ;
        RECT 233.930 69.840 236.120 70.010 ;
        RECT 233.930 69.670 234.245 69.840 ;
        RECT 233.915 69.420 234.245 69.670 ;
        RECT 227.040 68.430 232.385 68.975 ;
        RECT 233.480 68.640 233.820 69.150 ;
        RECT 233.990 68.430 234.260 69.230 ;
        RECT 234.440 68.700 234.720 69.670 ;
        RECT 234.900 68.700 235.200 69.670 ;
        RECT 235.380 68.705 235.730 69.670 ;
        RECT 235.950 68.930 236.120 69.840 ;
        RECT 236.290 69.110 236.530 70.420 ;
        RECT 236.700 69.890 240.210 70.980 ;
        RECT 236.700 69.200 238.350 69.720 ;
        RECT 238.520 69.370 240.210 69.890 ;
        RECT 235.950 68.600 236.445 68.930 ;
        RECT 236.700 68.430 240.210 69.200 ;
        RECT 241.300 68.600 241.560 70.810 ;
        RECT 241.730 70.600 242.060 70.980 ;
        RECT 242.485 70.430 242.655 70.810 ;
        RECT 242.915 70.600 243.245 70.980 ;
        RECT 243.440 70.430 243.610 70.810 ;
        RECT 243.820 70.600 244.150 70.980 ;
        RECT 244.400 70.430 244.590 70.810 ;
        RECT 244.830 70.600 245.160 70.980 ;
        RECT 245.470 70.480 245.730 70.810 ;
        RECT 241.730 70.260 243.680 70.430 ;
        RECT 241.730 69.340 241.900 70.260 ;
        RECT 242.270 69.670 242.465 69.980 ;
        RECT 242.735 69.670 242.920 69.980 ;
        RECT 242.210 69.340 242.465 69.670 ;
        RECT 242.690 69.340 242.920 69.670 ;
        RECT 241.730 68.430 242.060 68.810 ;
        RECT 242.270 68.765 242.465 69.340 ;
        RECT 242.735 68.760 242.920 69.340 ;
        RECT 243.170 68.770 243.340 69.670 ;
        RECT 243.510 69.270 243.680 70.260 ;
        RECT 243.850 70.260 244.590 70.430 ;
        RECT 243.850 69.750 244.020 70.260 ;
        RECT 244.190 69.920 244.770 70.090 ;
        RECT 245.040 69.970 245.390 70.300 ;
        RECT 244.600 69.800 244.770 69.920 ;
        RECT 245.560 69.800 245.730 70.480 ;
        RECT 245.990 69.970 246.160 70.810 ;
        RECT 246.330 70.640 247.500 70.810 ;
        RECT 246.330 70.140 246.660 70.640 ;
        RECT 247.170 70.600 247.500 70.640 ;
        RECT 247.690 70.560 248.045 70.980 ;
        RECT 246.830 70.380 247.060 70.470 ;
        RECT 248.215 70.380 248.465 70.810 ;
        RECT 246.830 70.140 248.465 70.380 ;
        RECT 248.635 70.220 248.965 70.980 ;
        RECT 249.135 70.140 249.390 70.810 ;
        RECT 245.990 69.800 249.050 69.970 ;
        RECT 243.850 69.580 244.420 69.750 ;
        RECT 244.600 69.630 245.730 69.800 ;
        RECT 243.510 68.940 244.060 69.270 ;
        RECT 244.250 69.100 244.420 69.580 ;
        RECT 244.590 69.290 245.210 69.460 ;
        RECT 245.000 69.110 245.210 69.290 ;
        RECT 244.250 68.770 244.650 69.100 ;
        RECT 245.560 68.930 245.730 69.630 ;
        RECT 245.905 69.420 246.255 69.630 ;
        RECT 246.425 69.420 246.870 69.620 ;
        RECT 247.040 69.420 247.515 69.620 ;
        RECT 243.170 68.600 244.650 68.770 ;
        RECT 244.830 68.430 245.160 68.810 ;
        RECT 245.470 68.600 245.730 68.930 ;
        RECT 245.990 69.080 247.055 69.250 ;
        RECT 245.990 68.600 246.160 69.080 ;
        RECT 246.330 68.430 246.660 68.910 ;
        RECT 246.885 68.850 247.055 69.080 ;
        RECT 247.235 69.020 247.515 69.420 ;
        RECT 247.785 69.420 248.115 69.620 ;
        RECT 248.285 69.420 248.650 69.620 ;
        RECT 247.785 69.020 248.070 69.420 ;
        RECT 248.880 69.250 249.050 69.800 ;
        RECT 248.250 69.080 249.050 69.250 ;
        RECT 248.250 68.850 248.420 69.080 ;
        RECT 249.220 69.010 249.390 70.140 ;
        RECT 249.580 69.890 252.170 70.980 ;
        RECT 249.205 68.940 249.390 69.010 ;
        RECT 249.180 68.930 249.390 68.940 ;
        RECT 246.885 68.600 248.420 68.850 ;
        RECT 248.590 68.430 248.920 68.910 ;
        RECT 249.135 68.600 249.390 68.930 ;
        RECT 249.580 69.200 250.790 69.720 ;
        RECT 250.960 69.370 252.170 69.890 ;
        RECT 252.340 69.815 252.630 70.980 ;
        RECT 252.800 69.890 256.310 70.980 ;
        RECT 256.480 69.890 257.690 70.980 ;
        RECT 252.800 69.200 254.450 69.720 ;
        RECT 254.620 69.370 256.310 69.890 ;
        RECT 249.580 68.430 252.170 69.200 ;
        RECT 252.340 68.430 252.630 69.155 ;
        RECT 252.800 68.430 256.310 69.200 ;
        RECT 256.480 69.180 257.000 69.720 ;
        RECT 257.170 69.350 257.690 69.890 ;
        RECT 257.950 69.970 258.120 70.810 ;
        RECT 258.290 70.640 259.460 70.810 ;
        RECT 258.290 70.140 258.620 70.640 ;
        RECT 259.130 70.600 259.460 70.640 ;
        RECT 259.650 70.560 260.005 70.980 ;
        RECT 258.790 70.380 259.020 70.470 ;
        RECT 260.175 70.380 260.425 70.810 ;
        RECT 258.790 70.140 260.425 70.380 ;
        RECT 260.595 70.220 260.925 70.980 ;
        RECT 261.095 70.140 261.350 70.810 ;
        RECT 261.140 70.130 261.350 70.140 ;
        RECT 257.950 69.800 261.010 69.970 ;
        RECT 257.865 69.420 258.215 69.630 ;
        RECT 258.385 69.420 258.830 69.620 ;
        RECT 259.000 69.420 259.475 69.620 ;
        RECT 256.480 68.430 257.690 69.180 ;
        RECT 257.950 69.080 259.015 69.250 ;
        RECT 257.950 68.600 258.120 69.080 ;
        RECT 258.290 68.430 258.620 68.910 ;
        RECT 258.845 68.850 259.015 69.080 ;
        RECT 259.195 69.020 259.475 69.420 ;
        RECT 259.745 69.420 260.075 69.620 ;
        RECT 260.245 69.420 260.610 69.620 ;
        RECT 259.745 69.020 260.030 69.420 ;
        RECT 260.840 69.250 261.010 69.800 ;
        RECT 260.210 69.080 261.010 69.250 ;
        RECT 260.210 68.850 260.380 69.080 ;
        RECT 261.180 69.010 261.350 70.130 ;
        RECT 261.630 69.970 261.800 70.810 ;
        RECT 261.970 70.640 263.140 70.810 ;
        RECT 261.970 70.140 262.300 70.640 ;
        RECT 262.810 70.600 263.140 70.640 ;
        RECT 263.330 70.560 263.685 70.980 ;
        RECT 262.470 70.380 262.700 70.470 ;
        RECT 263.855 70.380 264.105 70.810 ;
        RECT 262.470 70.140 264.105 70.380 ;
        RECT 264.275 70.220 264.605 70.980 ;
        RECT 264.775 70.140 265.030 70.810 ;
        RECT 265.220 70.470 266.410 70.760 ;
        RECT 261.630 69.800 264.690 69.970 ;
        RECT 261.545 69.420 261.895 69.630 ;
        RECT 262.065 69.420 262.510 69.620 ;
        RECT 262.680 69.420 263.155 69.620 ;
        RECT 261.165 68.930 261.350 69.010 ;
        RECT 258.845 68.600 260.380 68.850 ;
        RECT 260.550 68.430 260.880 68.910 ;
        RECT 261.095 68.600 261.350 68.930 ;
        RECT 261.630 69.080 262.695 69.250 ;
        RECT 261.630 68.600 261.800 69.080 ;
        RECT 261.970 68.430 262.300 68.910 ;
        RECT 262.525 68.850 262.695 69.080 ;
        RECT 262.875 69.020 263.155 69.420 ;
        RECT 263.425 69.420 263.755 69.620 ;
        RECT 263.925 69.450 264.300 69.620 ;
        RECT 263.925 69.420 264.290 69.450 ;
        RECT 263.425 69.020 263.710 69.420 ;
        RECT 264.520 69.250 264.690 69.800 ;
        RECT 263.890 69.080 264.690 69.250 ;
        RECT 263.890 68.850 264.060 69.080 ;
        RECT 264.860 69.010 265.030 70.140 ;
        RECT 265.240 70.130 266.410 70.300 ;
        RECT 266.580 70.180 266.860 70.980 ;
        RECT 265.240 69.840 265.565 70.130 ;
        RECT 266.240 70.010 266.410 70.130 ;
        RECT 265.735 69.670 265.930 69.960 ;
        RECT 266.240 69.840 266.900 70.010 ;
        RECT 267.070 69.840 267.345 70.810 ;
        RECT 267.520 69.890 269.190 70.980 ;
        RECT 270.005 70.620 270.455 70.980 ;
        RECT 271.020 70.620 271.350 70.980 ;
        RECT 271.920 70.620 272.255 70.980 ;
        RECT 272.780 70.620 273.110 70.980 ;
        RECT 266.730 69.670 266.900 69.840 ;
        RECT 265.220 69.340 265.565 69.670 ;
        RECT 265.735 69.340 266.560 69.670 ;
        RECT 266.730 69.340 267.005 69.670 ;
        RECT 266.730 69.170 266.900 69.340 ;
        RECT 264.845 68.930 265.030 69.010 ;
        RECT 262.525 68.600 264.060 68.850 ;
        RECT 264.230 68.430 264.560 68.910 ;
        RECT 264.775 68.600 265.030 68.930 ;
        RECT 265.235 69.000 266.900 69.170 ;
        RECT 267.175 69.105 267.345 69.840 ;
        RECT 265.235 68.650 265.490 69.000 ;
        RECT 265.660 68.430 265.990 68.830 ;
        RECT 266.160 68.650 266.330 69.000 ;
        RECT 266.500 68.430 266.880 68.830 ;
        RECT 267.070 68.760 267.345 69.105 ;
        RECT 267.520 69.200 268.270 69.720 ;
        RECT 268.440 69.370 269.190 69.890 ;
        RECT 269.425 69.840 269.785 70.510 ;
        RECT 269.955 70.220 273.720 70.450 ;
        RECT 267.520 68.430 269.190 69.200 ;
        RECT 269.425 69.150 269.645 69.840 ;
        RECT 269.955 69.670 270.125 70.220 ;
        RECT 270.555 69.870 271.330 70.040 ;
        RECT 271.500 69.880 272.810 70.050 ;
        RECT 271.160 69.700 271.330 69.870 ;
        RECT 269.815 69.340 270.125 69.670 ;
        RECT 269.425 68.890 269.910 69.150 ;
        RECT 270.295 69.070 270.510 69.685 ;
        RECT 270.800 69.340 270.990 69.685 ;
        RECT 271.160 69.365 272.375 69.700 ;
        RECT 271.160 69.150 271.390 69.365 ;
        RECT 272.545 69.190 272.810 69.880 ;
        RECT 270.695 68.960 271.390 69.150 ;
        RECT 271.560 68.960 272.810 69.190 ;
        RECT 272.990 68.960 273.270 70.050 ;
        RECT 270.695 68.890 270.875 68.960 ;
        RECT 269.425 68.700 270.875 68.890 ;
        RECT 271.560 68.860 271.750 68.960 ;
        RECT 269.425 68.600 269.910 68.700 ;
        RECT 271.055 68.430 271.385 68.790 ;
        RECT 271.920 68.430 272.250 68.790 ;
        RECT 272.420 68.600 272.610 68.960 ;
        RECT 272.780 68.430 273.110 68.790 ;
        RECT 273.440 68.770 273.720 70.220 ;
        RECT 273.960 69.890 275.170 70.980 ;
        RECT 275.350 70.260 275.680 70.980 ;
        RECT 273.960 69.180 274.480 69.720 ;
        RECT 274.650 69.350 275.170 69.890 ;
        RECT 275.340 69.620 275.570 69.960 ;
        RECT 275.860 69.620 276.075 70.735 ;
        RECT 276.270 70.035 276.600 70.810 ;
        RECT 276.770 70.205 277.480 70.980 ;
        RECT 276.270 69.820 277.420 70.035 ;
        RECT 275.340 69.420 275.670 69.620 ;
        RECT 275.860 69.440 276.310 69.620 ;
        RECT 275.980 69.420 276.310 69.440 ;
        RECT 276.480 69.420 276.950 69.650 ;
        RECT 277.135 69.250 277.420 69.820 ;
        RECT 277.650 69.375 277.930 70.810 ;
        RECT 278.100 69.815 278.390 70.980 ;
        RECT 278.565 70.310 278.820 70.810 ;
        RECT 278.990 70.480 279.320 70.980 ;
        RECT 278.565 70.140 279.315 70.310 ;
        RECT 273.960 68.430 275.170 69.180 ;
        RECT 275.340 69.060 276.520 69.250 ;
        RECT 275.340 68.600 275.680 69.060 ;
        RECT 276.190 68.980 276.520 69.060 ;
        RECT 276.710 69.060 277.420 69.250 ;
        RECT 276.710 68.920 277.010 69.060 ;
        RECT 276.695 68.910 277.010 68.920 ;
        RECT 276.685 68.900 277.010 68.910 ;
        RECT 276.675 68.895 277.010 68.900 ;
        RECT 275.850 68.430 276.020 68.890 ;
        RECT 276.670 68.885 277.010 68.895 ;
        RECT 276.665 68.880 277.010 68.885 ;
        RECT 276.660 68.870 277.010 68.880 ;
        RECT 276.655 68.865 277.010 68.870 ;
        RECT 276.650 68.600 277.010 68.865 ;
        RECT 277.250 68.430 277.420 68.890 ;
        RECT 277.590 68.600 277.930 69.375 ;
        RECT 278.565 69.320 278.915 69.970 ;
        RECT 278.100 68.430 278.390 69.155 ;
        RECT 279.085 69.150 279.315 70.140 ;
        RECT 278.565 68.980 279.315 69.150 ;
        RECT 278.565 68.690 278.820 68.980 ;
        RECT 278.990 68.430 279.320 68.810 ;
        RECT 279.490 68.690 279.660 70.810 ;
        RECT 279.830 70.010 280.155 70.795 ;
        RECT 280.325 70.520 280.575 70.980 ;
        RECT 280.745 70.480 280.995 70.810 ;
        RECT 281.210 70.480 281.890 70.810 ;
        RECT 280.745 70.350 280.915 70.480 ;
        RECT 280.520 70.180 280.915 70.350 ;
        RECT 279.890 68.960 280.350 70.010 ;
        RECT 280.520 68.820 280.690 70.180 ;
        RECT 281.085 69.920 281.550 70.310 ;
        RECT 280.860 69.110 281.210 69.730 ;
        RECT 281.380 69.330 281.550 69.920 ;
        RECT 281.720 69.700 281.890 70.480 ;
        RECT 282.060 70.380 282.230 70.720 ;
        RECT 282.465 70.550 282.795 70.980 ;
        RECT 282.965 70.380 283.135 70.720 ;
        RECT 283.430 70.520 283.800 70.980 ;
        RECT 282.060 70.210 283.135 70.380 ;
        RECT 283.970 70.350 284.140 70.810 ;
        RECT 284.375 70.470 285.245 70.810 ;
        RECT 285.415 70.520 285.665 70.980 ;
        RECT 283.580 70.180 284.140 70.350 ;
        RECT 283.580 70.040 283.750 70.180 ;
        RECT 282.250 69.870 283.750 70.040 ;
        RECT 284.445 70.010 284.905 70.300 ;
        RECT 281.720 69.530 283.410 69.700 ;
        RECT 281.380 69.110 281.735 69.330 ;
        RECT 281.905 68.820 282.075 69.530 ;
        RECT 282.280 69.110 283.070 69.360 ;
        RECT 283.240 69.350 283.410 69.530 ;
        RECT 283.580 69.180 283.750 69.870 ;
        RECT 280.020 68.430 280.350 68.790 ;
        RECT 280.520 68.650 281.015 68.820 ;
        RECT 281.220 68.650 282.075 68.820 ;
        RECT 282.950 68.430 283.280 68.890 ;
        RECT 283.490 68.790 283.750 69.180 ;
        RECT 283.940 70.000 284.905 70.010 ;
        RECT 285.075 70.090 285.245 70.470 ;
        RECT 285.835 70.430 286.005 70.720 ;
        RECT 286.185 70.600 286.515 70.980 ;
        RECT 285.835 70.260 286.635 70.430 ;
        RECT 283.940 69.840 284.615 70.000 ;
        RECT 285.075 69.920 286.295 70.090 ;
        RECT 283.940 69.050 284.150 69.840 ;
        RECT 285.075 69.830 285.245 69.920 ;
        RECT 284.320 69.050 284.670 69.670 ;
        RECT 284.840 69.660 285.245 69.830 ;
        RECT 284.840 68.880 285.010 69.660 ;
        RECT 285.180 69.210 285.400 69.490 ;
        RECT 285.580 69.380 286.120 69.750 ;
        RECT 286.465 69.670 286.635 70.260 ;
        RECT 286.855 69.840 287.160 70.980 ;
        RECT 287.330 69.790 287.585 70.670 ;
        RECT 287.760 69.890 291.270 70.980 ;
        RECT 291.445 70.310 291.700 70.810 ;
        RECT 291.870 70.480 292.200 70.980 ;
        RECT 291.445 70.140 292.195 70.310 ;
        RECT 286.465 69.640 287.205 69.670 ;
        RECT 285.180 69.040 285.710 69.210 ;
        RECT 283.490 68.620 283.840 68.790 ;
        RECT 284.060 68.600 285.010 68.880 ;
        RECT 285.180 68.430 285.370 68.870 ;
        RECT 285.540 68.810 285.710 69.040 ;
        RECT 285.880 68.980 286.120 69.380 ;
        RECT 286.290 69.340 287.205 69.640 ;
        RECT 286.290 69.165 286.615 69.340 ;
        RECT 286.290 68.810 286.610 69.165 ;
        RECT 287.375 69.140 287.585 69.790 ;
        RECT 285.540 68.640 286.610 68.810 ;
        RECT 286.855 68.430 287.160 68.890 ;
        RECT 287.330 68.610 287.585 69.140 ;
        RECT 287.760 69.200 289.410 69.720 ;
        RECT 289.580 69.370 291.270 69.890 ;
        RECT 291.445 69.320 291.795 69.970 ;
        RECT 287.760 68.430 291.270 69.200 ;
        RECT 291.965 69.150 292.195 70.140 ;
        RECT 291.445 68.980 292.195 69.150 ;
        RECT 291.445 68.690 291.700 68.980 ;
        RECT 291.870 68.430 292.200 68.810 ;
        RECT 292.370 68.690 292.540 70.810 ;
        RECT 292.710 70.010 293.035 70.795 ;
        RECT 293.205 70.520 293.455 70.980 ;
        RECT 293.625 70.480 293.875 70.810 ;
        RECT 294.090 70.480 294.770 70.810 ;
        RECT 293.625 70.350 293.795 70.480 ;
        RECT 293.400 70.180 293.795 70.350 ;
        RECT 292.770 68.960 293.230 70.010 ;
        RECT 293.400 68.820 293.570 70.180 ;
        RECT 293.965 69.920 294.430 70.310 ;
        RECT 293.740 69.110 294.090 69.730 ;
        RECT 294.260 69.330 294.430 69.920 ;
        RECT 294.600 69.700 294.770 70.480 ;
        RECT 294.940 70.380 295.110 70.720 ;
        RECT 295.345 70.550 295.675 70.980 ;
        RECT 295.845 70.380 296.015 70.720 ;
        RECT 296.310 70.520 296.680 70.980 ;
        RECT 294.940 70.210 296.015 70.380 ;
        RECT 296.850 70.350 297.020 70.810 ;
        RECT 297.255 70.470 298.125 70.810 ;
        RECT 298.295 70.520 298.545 70.980 ;
        RECT 296.460 70.180 297.020 70.350 ;
        RECT 296.460 70.040 296.630 70.180 ;
        RECT 295.130 69.870 296.630 70.040 ;
        RECT 297.325 70.010 297.785 70.300 ;
        RECT 294.600 69.530 296.290 69.700 ;
        RECT 294.260 69.110 294.615 69.330 ;
        RECT 294.785 68.820 294.955 69.530 ;
        RECT 295.160 69.110 295.950 69.360 ;
        RECT 296.120 69.350 296.290 69.530 ;
        RECT 296.460 69.180 296.630 69.870 ;
        RECT 292.900 68.430 293.230 68.790 ;
        RECT 293.400 68.650 293.895 68.820 ;
        RECT 294.100 68.650 294.955 68.820 ;
        RECT 295.830 68.430 296.160 68.890 ;
        RECT 296.370 68.790 296.630 69.180 ;
        RECT 296.820 70.000 297.785 70.010 ;
        RECT 297.955 70.090 298.125 70.470 ;
        RECT 298.715 70.430 298.885 70.720 ;
        RECT 299.065 70.600 299.395 70.980 ;
        RECT 298.715 70.260 299.515 70.430 ;
        RECT 296.820 69.840 297.495 70.000 ;
        RECT 297.955 69.920 299.175 70.090 ;
        RECT 296.820 69.050 297.030 69.840 ;
        RECT 297.955 69.830 298.125 69.920 ;
        RECT 297.200 69.050 297.550 69.670 ;
        RECT 297.720 69.660 298.125 69.830 ;
        RECT 297.720 68.880 297.890 69.660 ;
        RECT 298.060 69.210 298.280 69.490 ;
        RECT 298.460 69.380 299.000 69.750 ;
        RECT 299.345 69.670 299.515 70.260 ;
        RECT 299.735 69.840 300.040 70.980 ;
        RECT 300.210 69.790 300.465 70.670 ;
        RECT 301.155 70.110 301.440 70.980 ;
        RECT 301.610 70.350 301.870 70.810 ;
        RECT 302.045 70.520 302.300 70.980 ;
        RECT 302.470 70.350 302.730 70.810 ;
        RECT 301.610 70.180 302.730 70.350 ;
        RECT 302.900 70.180 303.210 70.980 ;
        RECT 301.610 69.930 301.870 70.180 ;
        RECT 303.380 70.010 303.690 70.810 ;
        RECT 299.345 69.640 300.085 69.670 ;
        RECT 298.060 69.040 298.590 69.210 ;
        RECT 296.370 68.620 296.720 68.790 ;
        RECT 296.940 68.600 297.890 68.880 ;
        RECT 298.060 68.430 298.250 68.870 ;
        RECT 298.420 68.810 298.590 69.040 ;
        RECT 298.760 68.980 299.000 69.380 ;
        RECT 299.170 69.340 300.085 69.640 ;
        RECT 299.170 69.165 299.495 69.340 ;
        RECT 299.170 68.810 299.490 69.165 ;
        RECT 300.255 69.140 300.465 69.790 ;
        RECT 298.420 68.640 299.490 68.810 ;
        RECT 299.735 68.430 300.040 68.890 ;
        RECT 300.210 68.610 300.465 69.140 ;
        RECT 301.115 69.760 301.870 69.930 ;
        RECT 302.660 69.840 303.690 70.010 ;
        RECT 301.115 69.250 301.520 69.760 ;
        RECT 302.660 69.590 302.830 69.840 ;
        RECT 301.690 69.420 302.830 69.590 ;
        RECT 301.115 69.080 302.765 69.250 ;
        RECT 303.000 69.100 303.350 69.670 ;
        RECT 301.160 68.430 301.440 68.910 ;
        RECT 301.610 68.690 301.870 69.080 ;
        RECT 302.045 68.430 302.300 68.910 ;
        RECT 302.470 68.690 302.765 69.080 ;
        RECT 303.520 68.930 303.690 69.840 ;
        RECT 303.860 69.815 304.150 70.980 ;
        RECT 304.325 69.840 304.660 70.810 ;
        RECT 304.830 69.840 305.000 70.980 ;
        RECT 305.170 70.640 307.200 70.810 ;
        RECT 304.325 69.170 304.495 69.840 ;
        RECT 305.170 69.670 305.340 70.640 ;
        RECT 304.665 69.340 304.920 69.670 ;
        RECT 305.145 69.340 305.340 69.670 ;
        RECT 305.510 70.300 306.635 70.470 ;
        RECT 304.750 69.170 304.920 69.340 ;
        RECT 305.510 69.170 305.680 70.300 ;
        RECT 302.945 68.430 303.220 68.910 ;
        RECT 303.390 68.600 303.690 68.930 ;
        RECT 303.860 68.430 304.150 69.155 ;
        RECT 304.325 68.600 304.580 69.170 ;
        RECT 304.750 69.000 305.680 69.170 ;
        RECT 305.850 69.960 306.860 70.130 ;
        RECT 305.850 69.160 306.020 69.960 ;
        RECT 306.225 69.620 306.500 69.760 ;
        RECT 306.220 69.450 306.500 69.620 ;
        RECT 305.505 68.965 305.680 69.000 ;
        RECT 304.750 68.430 305.080 68.830 ;
        RECT 305.505 68.600 306.035 68.965 ;
        RECT 306.225 68.600 306.500 69.450 ;
        RECT 306.670 68.600 306.860 69.960 ;
        RECT 307.030 69.975 307.200 70.640 ;
        RECT 307.370 70.220 307.540 70.980 ;
        RECT 307.775 70.220 308.290 70.630 ;
        RECT 307.030 69.785 307.780 69.975 ;
        RECT 307.950 69.410 308.290 70.220 ;
        RECT 308.460 69.890 309.670 70.980 ;
        RECT 307.060 69.240 308.290 69.410 ;
        RECT 307.040 68.430 307.550 68.965 ;
        RECT 307.770 68.635 308.015 69.240 ;
        RECT 308.460 69.180 308.980 69.720 ;
        RECT 309.150 69.350 309.670 69.890 ;
        RECT 309.840 69.890 311.050 70.980 ;
        RECT 309.840 69.350 310.360 69.890 ;
        RECT 310.530 69.180 311.050 69.720 ;
        RECT 308.460 68.430 309.670 69.180 ;
        RECT 309.840 68.430 311.050 69.180 ;
        RECT 162.095 68.260 311.135 68.430 ;
        RECT 162.180 67.510 163.390 68.260 ;
        RECT 162.180 66.970 162.700 67.510 ;
        RECT 163.560 67.490 166.150 68.260 ;
        RECT 166.785 67.550 167.040 68.080 ;
        RECT 167.210 67.800 167.515 68.260 ;
        RECT 167.760 67.880 168.830 68.050 ;
        RECT 162.870 66.800 163.390 67.340 ;
        RECT 163.560 66.970 164.770 67.490 ;
        RECT 164.940 66.800 166.150 67.320 ;
        RECT 162.180 65.710 163.390 66.800 ;
        RECT 163.560 65.710 166.150 66.800 ;
        RECT 166.785 66.900 166.995 67.550 ;
        RECT 167.760 67.525 168.080 67.880 ;
        RECT 167.755 67.350 168.080 67.525 ;
        RECT 167.165 67.050 168.080 67.350 ;
        RECT 168.250 67.310 168.490 67.710 ;
        RECT 168.660 67.650 168.830 67.880 ;
        RECT 169.000 67.820 169.190 68.260 ;
        RECT 169.360 67.810 170.310 68.090 ;
        RECT 170.530 67.900 170.880 68.070 ;
        RECT 168.660 67.480 169.190 67.650 ;
        RECT 167.165 67.020 167.905 67.050 ;
        RECT 166.785 66.020 167.040 66.900 ;
        RECT 167.210 65.710 167.515 66.850 ;
        RECT 167.735 66.430 167.905 67.020 ;
        RECT 168.250 66.940 168.790 67.310 ;
        RECT 168.970 67.200 169.190 67.480 ;
        RECT 169.360 67.030 169.530 67.810 ;
        RECT 169.125 66.860 169.530 67.030 ;
        RECT 169.700 67.020 170.050 67.640 ;
        RECT 169.125 66.770 169.295 66.860 ;
        RECT 170.220 66.850 170.430 67.640 ;
        RECT 168.075 66.600 169.295 66.770 ;
        RECT 169.755 66.690 170.430 66.850 ;
        RECT 167.735 66.260 168.535 66.430 ;
        RECT 167.855 65.710 168.185 66.090 ;
        RECT 168.365 65.970 168.535 66.260 ;
        RECT 169.125 66.220 169.295 66.600 ;
        RECT 169.465 66.680 170.430 66.690 ;
        RECT 170.620 67.510 170.880 67.900 ;
        RECT 171.090 67.800 171.420 68.260 ;
        RECT 172.295 67.870 173.150 68.040 ;
        RECT 173.355 67.870 173.850 68.040 ;
        RECT 174.020 67.900 174.350 68.260 ;
        RECT 170.620 66.820 170.790 67.510 ;
        RECT 170.960 67.160 171.130 67.340 ;
        RECT 171.300 67.330 172.090 67.580 ;
        RECT 172.295 67.160 172.465 67.870 ;
        RECT 172.635 67.360 172.990 67.580 ;
        RECT 170.960 66.990 172.650 67.160 ;
        RECT 169.465 66.390 169.925 66.680 ;
        RECT 170.620 66.650 172.120 66.820 ;
        RECT 170.620 66.510 170.790 66.650 ;
        RECT 170.230 66.340 170.790 66.510 ;
        RECT 168.705 65.710 168.955 66.170 ;
        RECT 169.125 65.880 169.995 66.220 ;
        RECT 170.230 65.880 170.400 66.340 ;
        RECT 171.235 66.310 172.310 66.480 ;
        RECT 170.570 65.710 170.940 66.170 ;
        RECT 171.235 65.970 171.405 66.310 ;
        RECT 171.575 65.710 171.905 66.140 ;
        RECT 172.140 65.970 172.310 66.310 ;
        RECT 172.480 66.210 172.650 66.990 ;
        RECT 172.820 66.770 172.990 67.360 ;
        RECT 173.160 66.960 173.510 67.580 ;
        RECT 172.820 66.380 173.285 66.770 ;
        RECT 173.680 66.510 173.850 67.870 ;
        RECT 174.020 66.680 174.480 67.730 ;
        RECT 173.455 66.340 173.850 66.510 ;
        RECT 173.455 66.210 173.625 66.340 ;
        RECT 172.480 65.880 173.160 66.210 ;
        RECT 173.375 65.880 173.625 66.210 ;
        RECT 173.795 65.710 174.045 66.170 ;
        RECT 174.215 65.895 174.540 66.680 ;
        RECT 174.710 65.880 174.880 68.000 ;
        RECT 175.050 67.880 175.380 68.260 ;
        RECT 175.550 67.710 175.805 68.000 ;
        RECT 175.055 67.540 175.805 67.710 ;
        RECT 176.905 67.710 177.160 68.000 ;
        RECT 177.330 67.880 177.660 68.260 ;
        RECT 176.905 67.540 177.655 67.710 ;
        RECT 175.055 66.550 175.285 67.540 ;
        RECT 175.455 66.720 175.805 67.370 ;
        RECT 176.905 66.720 177.255 67.370 ;
        RECT 177.425 66.550 177.655 67.540 ;
        RECT 175.055 66.380 175.805 66.550 ;
        RECT 175.050 65.710 175.380 66.210 ;
        RECT 175.550 65.880 175.805 66.380 ;
        RECT 176.905 66.380 177.655 66.550 ;
        RECT 176.905 65.880 177.160 66.380 ;
        RECT 177.330 65.710 177.660 66.210 ;
        RECT 177.830 65.880 178.000 68.000 ;
        RECT 178.360 67.900 178.690 68.260 ;
        RECT 178.860 67.870 179.355 68.040 ;
        RECT 179.560 67.870 180.415 68.040 ;
        RECT 178.230 66.680 178.690 67.730 ;
        RECT 178.170 65.895 178.495 66.680 ;
        RECT 178.860 66.510 179.030 67.870 ;
        RECT 179.200 66.960 179.550 67.580 ;
        RECT 179.720 67.360 180.075 67.580 ;
        RECT 179.720 66.770 179.890 67.360 ;
        RECT 180.245 67.160 180.415 67.870 ;
        RECT 181.290 67.800 181.620 68.260 ;
        RECT 181.830 67.900 182.180 68.070 ;
        RECT 180.620 67.330 181.410 67.580 ;
        RECT 181.830 67.510 182.090 67.900 ;
        RECT 182.400 67.810 183.350 68.090 ;
        RECT 183.520 67.820 183.710 68.260 ;
        RECT 183.880 67.880 184.950 68.050 ;
        RECT 181.580 67.160 181.750 67.340 ;
        RECT 178.860 66.340 179.255 66.510 ;
        RECT 179.425 66.380 179.890 66.770 ;
        RECT 180.060 66.990 181.750 67.160 ;
        RECT 179.085 66.210 179.255 66.340 ;
        RECT 180.060 66.210 180.230 66.990 ;
        RECT 181.920 66.820 182.090 67.510 ;
        RECT 180.590 66.650 182.090 66.820 ;
        RECT 182.280 66.850 182.490 67.640 ;
        RECT 182.660 67.020 183.010 67.640 ;
        RECT 183.180 67.030 183.350 67.810 ;
        RECT 183.880 67.650 184.050 67.880 ;
        RECT 183.520 67.480 184.050 67.650 ;
        RECT 183.520 67.200 183.740 67.480 ;
        RECT 184.220 67.310 184.460 67.710 ;
        RECT 183.180 66.860 183.585 67.030 ;
        RECT 183.920 66.940 184.460 67.310 ;
        RECT 184.630 67.525 184.950 67.880 ;
        RECT 185.195 67.800 185.500 68.260 ;
        RECT 185.670 67.550 185.920 68.080 ;
        RECT 184.630 67.350 184.955 67.525 ;
        RECT 184.630 67.050 185.545 67.350 ;
        RECT 184.805 67.020 185.545 67.050 ;
        RECT 182.280 66.690 182.955 66.850 ;
        RECT 183.415 66.770 183.585 66.860 ;
        RECT 182.280 66.680 183.245 66.690 ;
        RECT 181.920 66.510 182.090 66.650 ;
        RECT 178.665 65.710 178.915 66.170 ;
        RECT 179.085 65.880 179.335 66.210 ;
        RECT 179.550 65.880 180.230 66.210 ;
        RECT 180.400 66.310 181.475 66.480 ;
        RECT 181.920 66.340 182.480 66.510 ;
        RECT 182.785 66.390 183.245 66.680 ;
        RECT 183.415 66.600 184.635 66.770 ;
        RECT 180.400 65.970 180.570 66.310 ;
        RECT 180.805 65.710 181.135 66.140 ;
        RECT 181.305 65.970 181.475 66.310 ;
        RECT 181.770 65.710 182.140 66.170 ;
        RECT 182.310 65.880 182.480 66.340 ;
        RECT 183.415 66.220 183.585 66.600 ;
        RECT 184.805 66.430 184.975 67.020 ;
        RECT 185.715 66.900 185.920 67.550 ;
        RECT 186.090 67.505 186.340 68.260 ;
        RECT 186.560 67.510 187.770 68.260 ;
        RECT 187.940 67.535 188.230 68.260 ;
        RECT 188.410 67.920 189.600 68.090 ;
        RECT 188.410 67.750 188.720 67.920 ;
        RECT 186.560 66.970 187.080 67.510 ;
        RECT 182.715 65.880 183.585 66.220 ;
        RECT 184.175 66.260 184.975 66.430 ;
        RECT 183.755 65.710 184.005 66.170 ;
        RECT 184.175 65.970 184.345 66.260 ;
        RECT 184.525 65.710 184.855 66.090 ;
        RECT 185.195 65.710 185.500 66.850 ;
        RECT 185.670 66.020 185.920 66.900 ;
        RECT 186.090 65.710 186.340 66.850 ;
        RECT 187.250 66.800 187.770 67.340 ;
        RECT 188.405 66.945 188.720 67.580 ;
        RECT 186.560 65.710 187.770 66.800 ;
        RECT 187.940 65.710 188.230 66.875 ;
        RECT 188.410 65.710 188.720 66.775 ;
        RECT 188.890 66.560 189.100 67.750 ;
        RECT 189.270 67.630 189.600 67.920 ;
        RECT 189.840 67.800 190.010 68.260 ;
        RECT 190.240 67.630 190.570 68.090 ;
        RECT 190.750 67.800 190.920 68.260 ;
        RECT 191.100 67.630 191.430 68.090 ;
        RECT 191.625 67.860 191.960 68.260 ;
        RECT 192.130 67.690 192.335 68.090 ;
        RECT 192.545 67.780 192.820 68.260 ;
        RECT 193.030 67.760 193.290 68.090 ;
        RECT 189.270 67.460 191.430 67.630 ;
        RECT 191.650 67.520 192.335 67.690 ;
        RECT 189.440 66.900 189.935 67.270 ;
        RECT 190.115 67.070 190.915 67.270 ;
        RECT 191.085 66.900 191.415 67.290 ;
        RECT 189.440 66.730 191.415 66.900 ;
        RECT 188.890 66.380 190.540 66.560 ;
        RECT 188.890 65.880 189.125 66.380 ;
        RECT 190.240 66.220 190.540 66.380 ;
        RECT 189.295 65.710 189.625 66.170 ;
        RECT 189.820 66.050 190.010 66.210 ;
        RECT 190.710 66.050 190.930 66.560 ;
        RECT 189.820 65.880 190.930 66.050 ;
        RECT 191.100 65.710 191.430 66.560 ;
        RECT 191.650 66.490 191.990 67.520 ;
        RECT 192.160 66.850 192.410 67.350 ;
        RECT 192.590 67.020 192.950 67.600 ;
        RECT 193.120 66.850 193.290 67.760 ;
        RECT 193.460 67.490 196.050 68.260 ;
        RECT 193.460 66.970 194.670 67.490 ;
        RECT 196.680 67.460 197.020 68.090 ;
        RECT 197.190 67.460 197.440 68.260 ;
        RECT 197.630 67.610 197.960 68.090 ;
        RECT 198.130 67.800 198.355 68.260 ;
        RECT 198.525 67.610 198.855 68.090 ;
        RECT 192.160 66.680 193.290 66.850 ;
        RECT 194.840 66.800 196.050 67.320 ;
        RECT 191.650 66.315 192.315 66.490 ;
        RECT 191.625 65.710 191.960 66.135 ;
        RECT 192.130 65.910 192.315 66.315 ;
        RECT 192.520 65.710 192.850 66.490 ;
        RECT 193.020 65.910 193.290 66.680 ;
        RECT 193.460 65.710 196.050 66.800 ;
        RECT 196.680 66.850 196.855 67.460 ;
        RECT 197.630 67.440 198.855 67.610 ;
        RECT 199.485 67.480 199.985 68.090 ;
        RECT 200.450 67.710 200.620 68.090 ;
        RECT 200.835 67.880 201.165 68.260 ;
        RECT 200.450 67.540 201.165 67.710 ;
        RECT 197.025 67.100 197.720 67.270 ;
        RECT 197.895 67.240 198.315 67.270 ;
        RECT 197.550 66.850 197.720 67.100 ;
        RECT 197.890 67.070 198.315 67.240 ;
        RECT 198.485 67.070 198.815 67.270 ;
        RECT 198.985 67.070 199.315 67.270 ;
        RECT 199.485 66.850 199.655 67.480 ;
        RECT 199.840 67.020 200.190 67.270 ;
        RECT 200.360 66.990 200.715 67.360 ;
        RECT 200.995 67.350 201.165 67.540 ;
        RECT 201.335 67.515 201.590 68.090 ;
        RECT 200.995 67.020 201.250 67.350 ;
        RECT 196.680 65.880 197.020 66.850 ;
        RECT 197.190 65.710 197.360 66.850 ;
        RECT 197.550 66.680 199.985 66.850 ;
        RECT 200.995 66.810 201.165 67.020 ;
        RECT 197.630 65.710 197.880 66.510 ;
        RECT 198.525 65.880 198.855 66.680 ;
        RECT 199.155 65.710 199.485 66.510 ;
        RECT 199.655 65.880 199.985 66.680 ;
        RECT 200.450 66.640 201.165 66.810 ;
        RECT 201.420 66.785 201.590 67.515 ;
        RECT 201.765 67.420 202.025 68.260 ;
        RECT 202.200 67.715 207.545 68.260 ;
        RECT 203.785 66.885 204.125 67.715 ;
        RECT 207.720 67.630 208.060 68.090 ;
        RECT 208.230 67.800 208.400 68.260 ;
        RECT 209.030 67.825 209.390 68.090 ;
        RECT 209.035 67.820 209.390 67.825 ;
        RECT 209.040 67.810 209.390 67.820 ;
        RECT 209.045 67.805 209.390 67.810 ;
        RECT 209.050 67.795 209.390 67.805 ;
        RECT 209.630 67.800 209.800 68.260 ;
        RECT 209.055 67.790 209.390 67.795 ;
        RECT 209.065 67.780 209.390 67.790 ;
        RECT 209.075 67.770 209.390 67.780 ;
        RECT 208.570 67.630 208.900 67.710 ;
        RECT 207.720 67.440 208.900 67.630 ;
        RECT 209.090 67.630 209.390 67.770 ;
        RECT 209.090 67.440 209.800 67.630 ;
        RECT 200.450 65.880 200.620 66.640 ;
        RECT 200.835 65.710 201.165 66.470 ;
        RECT 201.335 65.880 201.590 66.785 ;
        RECT 201.765 65.710 202.025 66.860 ;
        RECT 205.605 66.145 205.955 67.395 ;
        RECT 207.720 67.070 208.050 67.270 ;
        RECT 208.360 67.250 208.690 67.270 ;
        RECT 208.240 67.070 208.690 67.250 ;
        RECT 207.720 66.730 207.950 67.070 ;
        RECT 202.200 65.710 207.545 66.145 ;
        RECT 207.730 65.710 208.060 66.430 ;
        RECT 208.240 65.955 208.455 67.070 ;
        RECT 208.860 67.040 209.330 67.270 ;
        RECT 209.515 66.870 209.800 67.440 ;
        RECT 209.970 67.315 210.310 68.090 ;
        RECT 210.810 67.860 211.140 68.260 ;
        RECT 211.310 67.690 211.640 68.030 ;
        RECT 212.690 67.860 213.020 68.260 ;
        RECT 208.650 66.655 209.800 66.870 ;
        RECT 208.650 65.880 208.980 66.655 ;
        RECT 209.150 65.710 209.860 66.485 ;
        RECT 210.030 65.880 210.310 67.315 ;
        RECT 210.655 67.520 213.020 67.690 ;
        RECT 213.190 67.535 213.520 68.045 ;
        RECT 213.700 67.535 213.990 68.260 ;
        RECT 210.655 66.520 210.825 67.520 ;
        RECT 212.850 67.350 213.020 67.520 ;
        RECT 210.995 66.690 211.240 67.350 ;
        RECT 211.455 66.690 211.720 67.350 ;
        RECT 211.915 66.690 212.200 67.350 ;
        RECT 212.375 67.020 212.680 67.350 ;
        RECT 212.850 67.020 213.160 67.350 ;
        RECT 212.375 66.690 212.590 67.020 ;
        RECT 210.655 66.350 211.110 66.520 ;
        RECT 210.780 65.920 211.110 66.350 ;
        RECT 211.290 66.350 212.580 66.520 ;
        RECT 211.290 65.930 211.540 66.350 ;
        RECT 211.770 65.710 212.100 66.180 ;
        RECT 212.330 65.930 212.580 66.350 ;
        RECT 212.770 65.710 213.020 66.850 ;
        RECT 213.330 66.770 213.520 67.535 ;
        RECT 214.160 67.460 214.500 68.090 ;
        RECT 214.670 67.460 214.920 68.260 ;
        RECT 215.110 67.610 215.440 68.090 ;
        RECT 215.610 67.800 215.835 68.260 ;
        RECT 216.005 67.610 216.335 68.090 ;
        RECT 213.190 65.920 213.520 66.770 ;
        RECT 213.700 65.710 213.990 66.875 ;
        RECT 214.160 66.850 214.335 67.460 ;
        RECT 215.110 67.440 216.335 67.610 ;
        RECT 216.965 67.480 217.465 68.090 ;
        RECT 217.845 67.495 218.300 68.260 ;
        RECT 218.575 67.880 219.875 68.090 ;
        RECT 220.130 67.900 220.460 68.260 ;
        RECT 219.705 67.730 219.875 67.880 ;
        RECT 220.630 67.760 220.890 68.090 ;
        RECT 214.505 67.100 215.200 67.270 ;
        RECT 215.030 66.850 215.200 67.100 ;
        RECT 215.375 67.070 215.795 67.270 ;
        RECT 215.965 67.070 216.295 67.270 ;
        RECT 216.465 67.070 216.795 67.270 ;
        RECT 216.965 66.850 217.135 67.480 ;
        RECT 218.775 67.270 218.995 67.670 ;
        RECT 217.320 67.020 217.670 67.270 ;
        RECT 217.840 67.070 218.330 67.270 ;
        RECT 218.520 67.060 218.995 67.270 ;
        RECT 219.240 67.270 219.450 67.670 ;
        RECT 219.705 67.605 220.460 67.730 ;
        RECT 219.705 67.560 220.550 67.605 ;
        RECT 220.280 67.440 220.550 67.560 ;
        RECT 219.240 67.060 219.570 67.270 ;
        RECT 219.740 67.000 220.150 67.305 ;
        RECT 214.160 65.880 214.500 66.850 ;
        RECT 214.670 65.710 214.840 66.850 ;
        RECT 215.030 66.680 217.465 66.850 ;
        RECT 215.110 65.710 215.360 66.510 ;
        RECT 216.005 65.880 216.335 66.680 ;
        RECT 216.635 65.710 216.965 66.510 ;
        RECT 217.135 65.880 217.465 66.680 ;
        RECT 217.845 66.830 219.020 66.890 ;
        RECT 220.380 66.865 220.550 67.440 ;
        RECT 220.350 66.830 220.550 66.865 ;
        RECT 217.845 66.720 220.550 66.830 ;
        RECT 217.845 66.100 218.100 66.720 ;
        RECT 218.690 66.660 220.490 66.720 ;
        RECT 218.690 66.630 219.020 66.660 ;
        RECT 220.720 66.560 220.890 67.760 ;
        RECT 221.060 67.490 222.730 68.260 ;
        RECT 222.900 67.880 224.285 68.090 ;
        RECT 222.900 67.610 223.190 67.880 ;
        RECT 223.360 67.520 223.785 67.710 ;
        RECT 223.955 67.690 224.285 67.880 ;
        RECT 224.520 67.860 224.850 68.260 ;
        RECT 225.025 67.690 225.355 68.090 ;
        RECT 225.560 67.700 225.730 68.260 ;
        RECT 223.955 67.520 225.355 67.690 ;
        RECT 225.900 67.520 226.410 68.090 ;
        RECT 221.060 66.970 221.810 67.490 ;
        RECT 221.980 66.800 222.730 67.320 ;
        RECT 222.900 67.020 223.175 67.350 ;
        RECT 218.350 66.460 218.535 66.550 ;
        RECT 219.125 66.460 219.960 66.470 ;
        RECT 218.350 66.260 219.960 66.460 ;
        RECT 218.350 66.220 218.580 66.260 ;
        RECT 217.845 65.880 218.180 66.100 ;
        RECT 219.185 65.710 219.540 66.090 ;
        RECT 219.710 65.880 219.960 66.260 ;
        RECT 220.210 65.710 220.460 66.490 ;
        RECT 220.630 65.880 220.890 66.560 ;
        RECT 221.060 65.710 222.730 66.800 ;
        RECT 222.900 65.710 223.190 66.850 ;
        RECT 223.360 66.510 223.530 67.520 ;
        RECT 223.700 66.685 224.055 67.350 ;
        RECT 224.240 66.685 224.515 67.350 ;
        RECT 224.685 67.020 225.030 67.350 ;
        RECT 225.320 67.270 225.490 67.350 ;
        RECT 225.860 67.270 226.050 67.350 ;
        RECT 225.240 67.020 225.490 67.270 ;
        RECT 225.685 67.020 226.050 67.270 ;
        RECT 223.360 66.260 224.315 66.510 ;
        RECT 223.985 66.050 224.315 66.260 ;
        RECT 224.685 66.220 225.010 67.020 ;
        RECT 225.685 66.850 225.855 67.020 ;
        RECT 226.235 66.850 226.410 67.520 ;
        RECT 225.180 66.680 225.855 66.850 ;
        RECT 225.180 66.050 225.350 66.680 ;
        RECT 223.985 65.880 225.350 66.050 ;
        RECT 225.520 65.710 225.810 66.510 ;
        RECT 226.025 65.890 226.410 66.850 ;
        RECT 227.040 67.800 227.600 68.090 ;
        RECT 227.770 67.800 228.020 68.260 ;
        RECT 227.040 66.430 227.290 67.800 ;
        RECT 228.640 67.630 228.970 67.990 ;
        RECT 229.340 67.715 234.685 68.260 ;
        RECT 227.580 67.440 228.970 67.630 ;
        RECT 227.580 67.350 227.750 67.440 ;
        RECT 227.460 67.020 227.750 67.350 ;
        RECT 227.920 67.020 228.260 67.270 ;
        RECT 228.480 67.020 229.155 67.270 ;
        RECT 227.580 66.770 227.750 67.020 ;
        RECT 227.580 66.600 228.520 66.770 ;
        RECT 228.890 66.660 229.155 67.020 ;
        RECT 230.925 66.885 231.265 67.715 ;
        RECT 234.860 67.490 238.370 68.260 ;
        RECT 239.460 67.535 239.750 68.260 ;
        RECT 240.010 67.780 240.310 68.260 ;
        RECT 240.480 67.610 240.740 68.065 ;
        RECT 240.910 67.780 241.170 68.260 ;
        RECT 241.350 67.610 241.610 68.065 ;
        RECT 241.780 67.780 242.030 68.260 ;
        RECT 242.210 67.610 242.470 68.065 ;
        RECT 242.640 67.780 242.890 68.260 ;
        RECT 243.070 67.610 243.330 68.065 ;
        RECT 243.500 67.780 243.745 68.260 ;
        RECT 243.915 67.610 244.190 68.065 ;
        RECT 244.360 67.780 244.605 68.260 ;
        RECT 244.775 67.610 245.035 68.065 ;
        RECT 245.205 67.780 245.465 68.260 ;
        RECT 245.635 67.610 245.895 68.065 ;
        RECT 246.065 67.780 246.325 68.260 ;
        RECT 246.495 67.610 246.755 68.065 ;
        RECT 246.925 67.700 247.185 68.260 ;
        RECT 227.040 65.880 227.500 66.430 ;
        RECT 227.690 65.710 228.020 66.430 ;
        RECT 228.220 66.050 228.520 66.600 ;
        RECT 228.690 65.710 228.970 66.380 ;
        RECT 232.745 66.145 233.095 67.395 ;
        RECT 234.860 66.970 236.510 67.490 ;
        RECT 240.010 67.440 246.755 67.610 ;
        RECT 236.680 66.800 238.370 67.320 ;
        RECT 229.340 65.710 234.685 66.145 ;
        RECT 234.860 65.710 238.370 66.800 ;
        RECT 239.460 65.710 239.750 66.875 ;
        RECT 240.010 66.850 241.175 67.440 ;
        RECT 247.355 67.270 247.605 68.080 ;
        RECT 247.785 67.735 248.045 68.260 ;
        RECT 248.215 67.270 248.465 68.080 ;
        RECT 248.645 67.750 248.950 68.260 ;
        RECT 249.120 67.715 254.465 68.260 ;
        RECT 241.345 67.020 248.465 67.270 ;
        RECT 248.635 67.020 248.950 67.580 ;
        RECT 240.010 66.625 246.755 66.850 ;
        RECT 240.010 65.710 240.280 66.455 ;
        RECT 240.450 65.885 240.740 66.625 ;
        RECT 241.350 66.610 246.755 66.625 ;
        RECT 240.910 65.715 241.165 66.440 ;
        RECT 241.350 65.885 241.610 66.610 ;
        RECT 241.780 65.715 242.025 66.440 ;
        RECT 242.210 65.885 242.470 66.610 ;
        RECT 242.640 65.715 242.885 66.440 ;
        RECT 243.070 65.885 243.330 66.610 ;
        RECT 243.500 65.715 243.745 66.440 ;
        RECT 243.915 65.885 244.175 66.610 ;
        RECT 244.345 65.715 244.605 66.440 ;
        RECT 244.775 65.885 245.035 66.610 ;
        RECT 245.205 65.715 245.465 66.440 ;
        RECT 245.635 65.885 245.895 66.610 ;
        RECT 246.065 65.715 246.325 66.440 ;
        RECT 246.495 65.885 246.755 66.610 ;
        RECT 246.925 65.715 247.185 66.510 ;
        RECT 247.355 65.885 247.605 67.020 ;
        RECT 240.910 65.710 247.185 65.715 ;
        RECT 247.785 65.710 248.045 66.520 ;
        RECT 248.220 65.880 248.465 67.020 ;
        RECT 250.705 66.885 251.045 67.715 ;
        RECT 254.640 67.490 258.150 68.260 ;
        RECT 258.520 67.630 258.850 67.990 ;
        RECT 259.470 67.800 259.720 68.260 ;
        RECT 259.890 67.800 260.450 68.090 ;
        RECT 248.645 65.710 248.940 66.520 ;
        RECT 252.525 66.145 252.875 67.395 ;
        RECT 254.640 66.970 256.290 67.490 ;
        RECT 258.520 67.440 259.910 67.630 ;
        RECT 259.740 67.350 259.910 67.440 ;
        RECT 256.460 66.800 258.150 67.320 ;
        RECT 249.120 65.710 254.465 66.145 ;
        RECT 254.640 65.710 258.150 66.800 ;
        RECT 258.335 67.020 259.010 67.270 ;
        RECT 259.230 67.020 259.570 67.270 ;
        RECT 259.740 67.020 260.030 67.350 ;
        RECT 258.335 66.660 258.600 67.020 ;
        RECT 259.740 66.770 259.910 67.020 ;
        RECT 258.970 66.600 259.910 66.770 ;
        RECT 258.520 65.710 258.800 66.380 ;
        RECT 258.970 66.050 259.270 66.600 ;
        RECT 260.200 66.430 260.450 67.800 ;
        RECT 259.470 65.710 259.800 66.430 ;
        RECT 259.990 65.880 260.450 66.430 ;
        RECT 260.620 67.585 260.890 67.930 ;
        RECT 261.080 67.860 261.460 68.260 ;
        RECT 261.630 67.690 261.800 68.040 ;
        RECT 261.970 67.860 262.300 68.260 ;
        RECT 262.500 67.690 262.670 68.040 ;
        RECT 262.870 67.760 263.200 68.260 ;
        RECT 260.620 66.850 260.790 67.585 ;
        RECT 261.060 67.520 262.670 67.690 ;
        RECT 261.060 67.350 261.230 67.520 ;
        RECT 260.960 67.020 261.230 67.350 ;
        RECT 261.400 67.020 261.805 67.350 ;
        RECT 261.060 66.850 261.230 67.020 ;
        RECT 260.620 65.880 260.890 66.850 ;
        RECT 261.060 66.680 261.785 66.850 ;
        RECT 261.975 66.730 262.685 67.350 ;
        RECT 262.855 67.020 263.205 67.590 ;
        RECT 263.380 67.490 265.050 68.260 ;
        RECT 265.220 67.535 265.510 68.260 ;
        RECT 265.680 67.490 269.190 68.260 ;
        RECT 269.360 67.510 270.570 68.260 ;
        RECT 263.380 66.970 264.130 67.490 ;
        RECT 261.615 66.560 261.785 66.680 ;
        RECT 262.885 66.560 263.205 66.850 ;
        RECT 264.300 66.800 265.050 67.320 ;
        RECT 265.680 66.970 267.330 67.490 ;
        RECT 261.100 65.710 261.380 66.510 ;
        RECT 261.615 66.390 263.205 66.560 ;
        RECT 261.550 65.930 263.205 66.220 ;
        RECT 263.380 65.710 265.050 66.800 ;
        RECT 265.220 65.710 265.510 66.875 ;
        RECT 267.500 66.800 269.190 67.320 ;
        RECT 269.360 66.970 269.880 67.510 ;
        RECT 270.745 67.440 271.020 68.260 ;
        RECT 271.190 67.620 271.520 68.090 ;
        RECT 271.690 67.790 271.860 68.260 ;
        RECT 272.030 67.620 272.360 68.090 ;
        RECT 272.530 67.790 272.820 68.260 ;
        RECT 273.040 67.715 278.385 68.260 ;
        RECT 271.190 67.610 272.360 67.620 ;
        RECT 271.190 67.580 272.790 67.610 ;
        RECT 271.190 67.440 272.810 67.580 ;
        RECT 272.575 67.410 272.810 67.440 ;
        RECT 270.050 66.800 270.570 67.340 ;
        RECT 270.745 67.070 271.465 67.270 ;
        RECT 271.635 67.070 272.405 67.270 ;
        RECT 272.575 66.900 272.790 67.410 ;
        RECT 265.680 65.710 269.190 66.800 ;
        RECT 269.360 65.710 270.570 66.800 ;
        RECT 270.745 66.680 271.860 66.890 ;
        RECT 270.745 65.880 271.020 66.680 ;
        RECT 271.190 65.710 271.520 66.510 ;
        RECT 271.690 66.050 271.860 66.680 ;
        RECT 272.030 66.680 272.790 66.900 ;
        RECT 274.625 66.885 274.965 67.715 ;
        RECT 279.485 67.520 279.740 68.090 ;
        RECT 279.910 67.860 280.240 68.260 ;
        RECT 280.665 67.725 281.195 68.090 ;
        RECT 280.665 67.690 280.840 67.725 ;
        RECT 279.910 67.520 280.840 67.690 ;
        RECT 272.030 66.220 272.360 66.680 ;
        RECT 272.530 66.050 272.830 66.510 ;
        RECT 276.445 66.145 276.795 67.395 ;
        RECT 279.485 66.850 279.655 67.520 ;
        RECT 279.910 67.350 280.080 67.520 ;
        RECT 279.825 67.020 280.080 67.350 ;
        RECT 280.305 67.020 280.500 67.350 ;
        RECT 271.690 65.880 272.830 66.050 ;
        RECT 273.040 65.710 278.385 66.145 ;
        RECT 279.485 65.880 279.820 66.850 ;
        RECT 279.990 65.710 280.160 66.850 ;
        RECT 280.330 66.050 280.500 67.020 ;
        RECT 280.670 66.390 280.840 67.520 ;
        RECT 281.010 66.730 281.180 67.530 ;
        RECT 281.385 67.240 281.660 68.090 ;
        RECT 281.380 67.070 281.660 67.240 ;
        RECT 281.385 66.930 281.660 67.070 ;
        RECT 281.830 66.730 282.020 68.090 ;
        RECT 282.200 67.725 282.710 68.260 ;
        RECT 282.930 67.450 283.175 68.055 ;
        RECT 283.620 67.630 283.960 68.090 ;
        RECT 284.130 67.800 284.300 68.260 ;
        RECT 284.930 67.825 285.290 68.090 ;
        RECT 284.935 67.820 285.290 67.825 ;
        RECT 284.940 67.810 285.290 67.820 ;
        RECT 284.945 67.805 285.290 67.810 ;
        RECT 284.950 67.795 285.290 67.805 ;
        RECT 285.530 67.800 285.700 68.260 ;
        RECT 284.955 67.790 285.290 67.795 ;
        RECT 284.965 67.780 285.290 67.790 ;
        RECT 284.975 67.770 285.290 67.780 ;
        RECT 284.470 67.630 284.800 67.710 ;
        RECT 282.220 67.280 283.450 67.450 ;
        RECT 283.620 67.440 284.800 67.630 ;
        RECT 284.990 67.630 285.290 67.770 ;
        RECT 284.990 67.440 285.700 67.630 ;
        RECT 281.010 66.560 282.020 66.730 ;
        RECT 282.190 66.715 282.940 66.905 ;
        RECT 280.670 66.220 281.795 66.390 ;
        RECT 282.190 66.050 282.360 66.715 ;
        RECT 283.110 66.470 283.450 67.280 ;
        RECT 283.620 67.070 283.950 67.270 ;
        RECT 284.260 67.250 284.590 67.270 ;
        RECT 284.140 67.070 284.590 67.250 ;
        RECT 283.620 66.730 283.850 67.070 ;
        RECT 280.330 65.880 282.360 66.050 ;
        RECT 282.530 65.710 282.700 66.470 ;
        RECT 282.935 66.060 283.450 66.470 ;
        RECT 283.630 65.710 283.960 66.430 ;
        RECT 284.140 65.955 284.355 67.070 ;
        RECT 284.760 67.040 285.230 67.270 ;
        RECT 285.415 66.870 285.700 67.440 ;
        RECT 285.870 67.315 286.210 68.090 ;
        RECT 284.550 66.655 285.700 66.870 ;
        RECT 284.550 65.880 284.880 66.655 ;
        RECT 285.050 65.710 285.760 66.485 ;
        RECT 285.930 65.880 286.210 67.315 ;
        RECT 286.380 67.490 289.890 68.260 ;
        RECT 290.980 67.535 291.270 68.260 ;
        RECT 291.445 67.520 291.700 68.090 ;
        RECT 291.870 67.860 292.200 68.260 ;
        RECT 292.625 67.725 293.155 68.090 ;
        RECT 293.345 67.920 293.620 68.090 ;
        RECT 293.340 67.750 293.620 67.920 ;
        RECT 292.625 67.690 292.800 67.725 ;
        RECT 291.870 67.520 292.800 67.690 ;
        RECT 286.380 66.970 288.030 67.490 ;
        RECT 288.200 66.800 289.890 67.320 ;
        RECT 286.380 65.710 289.890 66.800 ;
        RECT 290.980 65.710 291.270 66.875 ;
        RECT 291.445 66.850 291.615 67.520 ;
        RECT 291.870 67.350 292.040 67.520 ;
        RECT 291.785 67.020 292.040 67.350 ;
        RECT 292.265 67.020 292.460 67.350 ;
        RECT 291.445 65.880 291.780 66.850 ;
        RECT 291.950 65.710 292.120 66.850 ;
        RECT 292.290 66.050 292.460 67.020 ;
        RECT 292.630 66.390 292.800 67.520 ;
        RECT 292.970 66.730 293.140 67.530 ;
        RECT 293.345 66.930 293.620 67.750 ;
        RECT 293.790 66.730 293.980 68.090 ;
        RECT 294.160 67.725 294.670 68.260 ;
        RECT 294.890 67.450 295.135 68.055 ;
        RECT 295.580 67.490 298.170 68.260 ;
        RECT 298.805 67.710 299.060 68.000 ;
        RECT 299.230 67.880 299.560 68.260 ;
        RECT 298.805 67.540 299.555 67.710 ;
        RECT 294.180 67.280 295.410 67.450 ;
        RECT 292.970 66.560 293.980 66.730 ;
        RECT 294.150 66.715 294.900 66.905 ;
        RECT 292.630 66.220 293.755 66.390 ;
        RECT 294.150 66.050 294.320 66.715 ;
        RECT 295.070 66.470 295.410 67.280 ;
        RECT 295.580 66.970 296.790 67.490 ;
        RECT 296.960 66.800 298.170 67.320 ;
        RECT 292.290 65.880 294.320 66.050 ;
        RECT 294.490 65.710 294.660 66.470 ;
        RECT 294.895 66.060 295.410 66.470 ;
        RECT 295.580 65.710 298.170 66.800 ;
        RECT 298.805 66.720 299.155 67.370 ;
        RECT 299.325 66.550 299.555 67.540 ;
        RECT 298.805 66.380 299.555 66.550 ;
        RECT 298.805 65.880 299.060 66.380 ;
        RECT 299.230 65.710 299.560 66.210 ;
        RECT 299.730 65.880 299.900 68.000 ;
        RECT 300.260 67.900 300.590 68.260 ;
        RECT 300.760 67.870 301.255 68.040 ;
        RECT 301.460 67.870 302.315 68.040 ;
        RECT 300.130 66.680 300.590 67.730 ;
        RECT 300.070 65.895 300.395 66.680 ;
        RECT 300.760 66.510 300.930 67.870 ;
        RECT 301.100 66.960 301.450 67.580 ;
        RECT 301.620 67.360 301.975 67.580 ;
        RECT 301.620 66.770 301.790 67.360 ;
        RECT 302.145 67.160 302.315 67.870 ;
        RECT 303.190 67.800 303.520 68.260 ;
        RECT 303.730 67.900 304.080 68.070 ;
        RECT 302.520 67.330 303.310 67.580 ;
        RECT 303.730 67.510 303.990 67.900 ;
        RECT 304.300 67.810 305.250 68.090 ;
        RECT 305.420 67.820 305.610 68.260 ;
        RECT 305.780 67.880 306.850 68.050 ;
        RECT 303.480 67.160 303.650 67.340 ;
        RECT 300.760 66.340 301.155 66.510 ;
        RECT 301.325 66.380 301.790 66.770 ;
        RECT 301.960 66.990 303.650 67.160 ;
        RECT 300.985 66.210 301.155 66.340 ;
        RECT 301.960 66.210 302.130 66.990 ;
        RECT 303.820 66.820 303.990 67.510 ;
        RECT 302.490 66.650 303.990 66.820 ;
        RECT 304.180 66.850 304.390 67.640 ;
        RECT 304.560 67.020 304.910 67.640 ;
        RECT 305.080 67.030 305.250 67.810 ;
        RECT 305.780 67.650 305.950 67.880 ;
        RECT 305.420 67.480 305.950 67.650 ;
        RECT 305.420 67.200 305.640 67.480 ;
        RECT 306.120 67.310 306.360 67.710 ;
        RECT 305.080 66.860 305.485 67.030 ;
        RECT 305.820 66.940 306.360 67.310 ;
        RECT 306.530 67.525 306.850 67.880 ;
        RECT 307.095 67.800 307.400 68.260 ;
        RECT 307.570 67.550 307.820 68.080 ;
        RECT 306.530 67.350 306.855 67.525 ;
        RECT 306.530 67.050 307.445 67.350 ;
        RECT 306.705 67.020 307.445 67.050 ;
        RECT 304.180 66.690 304.855 66.850 ;
        RECT 305.315 66.770 305.485 66.860 ;
        RECT 304.180 66.680 305.145 66.690 ;
        RECT 303.820 66.510 303.990 66.650 ;
        RECT 300.565 65.710 300.815 66.170 ;
        RECT 300.985 65.880 301.235 66.210 ;
        RECT 301.450 65.880 302.130 66.210 ;
        RECT 302.300 66.310 303.375 66.480 ;
        RECT 303.820 66.340 304.380 66.510 ;
        RECT 304.685 66.390 305.145 66.680 ;
        RECT 305.315 66.600 306.535 66.770 ;
        RECT 302.300 65.970 302.470 66.310 ;
        RECT 302.705 65.710 303.035 66.140 ;
        RECT 303.205 65.970 303.375 66.310 ;
        RECT 303.670 65.710 304.040 66.170 ;
        RECT 304.210 65.880 304.380 66.340 ;
        RECT 305.315 66.220 305.485 66.600 ;
        RECT 306.705 66.430 306.875 67.020 ;
        RECT 307.615 66.900 307.820 67.550 ;
        RECT 307.990 67.505 308.240 68.260 ;
        RECT 308.460 67.585 308.720 68.090 ;
        RECT 308.900 67.880 309.230 68.260 ;
        RECT 309.410 67.710 309.580 68.090 ;
        RECT 304.615 65.880 305.485 66.220 ;
        RECT 306.075 66.260 306.875 66.430 ;
        RECT 305.655 65.710 305.905 66.170 ;
        RECT 306.075 65.970 306.245 66.260 ;
        RECT 306.425 65.710 306.755 66.090 ;
        RECT 307.095 65.710 307.400 66.850 ;
        RECT 307.570 66.020 307.820 66.900 ;
        RECT 307.990 65.710 308.240 66.850 ;
        RECT 308.460 66.785 308.630 67.585 ;
        RECT 308.915 67.540 309.580 67.710 ;
        RECT 308.915 67.285 309.085 67.540 ;
        RECT 309.840 67.510 311.050 68.260 ;
        RECT 308.800 66.955 309.085 67.285 ;
        RECT 309.320 66.990 309.650 67.360 ;
        RECT 308.915 66.810 309.085 66.955 ;
        RECT 308.460 65.880 308.730 66.785 ;
        RECT 308.915 66.640 309.580 66.810 ;
        RECT 308.900 65.710 309.230 66.470 ;
        RECT 309.410 65.880 309.580 66.640 ;
        RECT 309.840 66.800 310.360 67.340 ;
        RECT 310.530 66.970 311.050 67.510 ;
        RECT 309.840 65.710 311.050 66.800 ;
        RECT 162.095 65.540 311.135 65.710 ;
        RECT 162.180 64.450 163.390 65.540 ;
        RECT 163.560 64.450 165.230 65.540 ;
        RECT 162.180 63.740 162.700 64.280 ;
        RECT 162.870 63.910 163.390 64.450 ;
        RECT 163.560 63.760 164.310 64.280 ;
        RECT 164.480 63.930 165.230 64.450 ;
        RECT 165.450 64.400 165.700 65.540 ;
        RECT 165.870 64.350 166.120 65.230 ;
        RECT 166.290 64.400 166.595 65.540 ;
        RECT 166.935 65.160 167.265 65.540 ;
        RECT 167.445 64.990 167.615 65.280 ;
        RECT 167.785 65.080 168.035 65.540 ;
        RECT 166.815 64.820 167.615 64.990 ;
        RECT 168.205 65.030 169.075 65.370 ;
        RECT 162.180 62.990 163.390 63.740 ;
        RECT 163.560 62.990 165.230 63.760 ;
        RECT 165.450 62.990 165.700 63.745 ;
        RECT 165.870 63.700 166.075 64.350 ;
        RECT 166.815 64.230 166.985 64.820 ;
        RECT 168.205 64.650 168.375 65.030 ;
        RECT 169.310 64.910 169.480 65.370 ;
        RECT 169.650 65.080 170.020 65.540 ;
        RECT 170.315 64.940 170.485 65.280 ;
        RECT 170.655 65.110 170.985 65.540 ;
        RECT 171.220 64.940 171.390 65.280 ;
        RECT 167.155 64.480 168.375 64.650 ;
        RECT 168.545 64.570 169.005 64.860 ;
        RECT 169.310 64.740 169.870 64.910 ;
        RECT 170.315 64.770 171.390 64.940 ;
        RECT 171.560 65.040 172.240 65.370 ;
        RECT 172.455 65.040 172.705 65.370 ;
        RECT 172.875 65.080 173.125 65.540 ;
        RECT 169.700 64.600 169.870 64.740 ;
        RECT 168.545 64.560 169.510 64.570 ;
        RECT 168.205 64.390 168.375 64.480 ;
        RECT 168.835 64.400 169.510 64.560 ;
        RECT 166.245 64.200 166.985 64.230 ;
        RECT 166.245 63.900 167.160 64.200 ;
        RECT 166.835 63.725 167.160 63.900 ;
        RECT 165.870 63.170 166.120 63.700 ;
        RECT 166.290 62.990 166.595 63.450 ;
        RECT 166.840 63.370 167.160 63.725 ;
        RECT 167.330 63.940 167.870 64.310 ;
        RECT 168.205 64.220 168.610 64.390 ;
        RECT 167.330 63.540 167.570 63.940 ;
        RECT 168.050 63.770 168.270 64.050 ;
        RECT 167.740 63.600 168.270 63.770 ;
        RECT 167.740 63.370 167.910 63.600 ;
        RECT 168.440 63.440 168.610 64.220 ;
        RECT 168.780 63.610 169.130 64.230 ;
        RECT 169.300 63.610 169.510 64.400 ;
        RECT 169.700 64.430 171.200 64.600 ;
        RECT 169.700 63.740 169.870 64.430 ;
        RECT 171.560 64.260 171.730 65.040 ;
        RECT 172.535 64.910 172.705 65.040 ;
        RECT 170.040 64.090 171.730 64.260 ;
        RECT 171.900 64.480 172.365 64.870 ;
        RECT 172.535 64.740 172.930 64.910 ;
        RECT 170.040 63.910 170.210 64.090 ;
        RECT 166.840 63.200 167.910 63.370 ;
        RECT 168.080 62.990 168.270 63.430 ;
        RECT 168.440 63.160 169.390 63.440 ;
        RECT 169.700 63.350 169.960 63.740 ;
        RECT 170.380 63.670 171.170 63.920 ;
        RECT 169.610 63.180 169.960 63.350 ;
        RECT 170.170 62.990 170.500 63.450 ;
        RECT 171.375 63.380 171.545 64.090 ;
        RECT 171.900 63.890 172.070 64.480 ;
        RECT 171.715 63.670 172.070 63.890 ;
        RECT 172.240 63.670 172.590 64.290 ;
        RECT 172.760 63.380 172.930 64.740 ;
        RECT 173.295 64.570 173.620 65.355 ;
        RECT 173.100 63.520 173.560 64.570 ;
        RECT 171.375 63.210 172.230 63.380 ;
        RECT 172.435 63.210 172.930 63.380 ;
        RECT 173.100 62.990 173.430 63.350 ;
        RECT 173.790 63.250 173.960 65.370 ;
        RECT 174.130 65.040 174.460 65.540 ;
        RECT 174.630 64.870 174.885 65.370 ;
        RECT 174.135 64.700 174.885 64.870 ;
        RECT 174.135 63.710 174.365 64.700 ;
        RECT 174.535 63.880 174.885 64.530 ;
        RECT 175.060 64.375 175.350 65.540 ;
        RECT 175.525 64.400 175.860 65.370 ;
        RECT 176.030 64.400 176.200 65.540 ;
        RECT 176.370 65.200 178.400 65.370 ;
        RECT 175.525 63.730 175.695 64.400 ;
        RECT 176.370 64.230 176.540 65.200 ;
        RECT 175.865 63.900 176.120 64.230 ;
        RECT 176.345 63.900 176.540 64.230 ;
        RECT 176.710 64.860 177.835 65.030 ;
        RECT 175.950 63.730 176.120 63.900 ;
        RECT 176.710 63.730 176.880 64.860 ;
        RECT 174.135 63.540 174.885 63.710 ;
        RECT 174.130 62.990 174.460 63.370 ;
        RECT 174.630 63.250 174.885 63.540 ;
        RECT 175.060 62.990 175.350 63.715 ;
        RECT 175.525 63.160 175.780 63.730 ;
        RECT 175.950 63.560 176.880 63.730 ;
        RECT 177.050 64.520 178.060 64.690 ;
        RECT 177.050 63.720 177.220 64.520 ;
        RECT 177.425 64.180 177.700 64.320 ;
        RECT 177.420 64.010 177.700 64.180 ;
        RECT 176.705 63.525 176.880 63.560 ;
        RECT 175.950 62.990 176.280 63.390 ;
        RECT 176.705 63.160 177.235 63.525 ;
        RECT 177.425 63.160 177.700 64.010 ;
        RECT 177.870 63.160 178.060 64.520 ;
        RECT 178.230 64.535 178.400 65.200 ;
        RECT 178.570 64.780 178.740 65.540 ;
        RECT 178.975 64.780 179.490 65.190 ;
        RECT 178.230 64.345 178.980 64.535 ;
        RECT 179.150 63.970 179.490 64.780 ;
        RECT 178.260 63.800 179.490 63.970 ;
        RECT 180.585 64.400 180.920 65.370 ;
        RECT 181.090 64.400 181.260 65.540 ;
        RECT 181.430 65.200 183.460 65.370 ;
        RECT 178.240 62.990 178.750 63.525 ;
        RECT 178.970 63.195 179.215 63.800 ;
        RECT 180.585 63.730 180.755 64.400 ;
        RECT 181.430 64.230 181.600 65.200 ;
        RECT 180.925 63.900 181.180 64.230 ;
        RECT 181.405 63.900 181.600 64.230 ;
        RECT 181.770 64.860 182.895 65.030 ;
        RECT 181.010 63.730 181.180 63.900 ;
        RECT 181.770 63.730 181.940 64.860 ;
        RECT 180.585 63.160 180.840 63.730 ;
        RECT 181.010 63.560 181.940 63.730 ;
        RECT 182.110 64.520 183.120 64.690 ;
        RECT 182.110 63.720 182.280 64.520 ;
        RECT 182.485 63.840 182.760 64.320 ;
        RECT 182.480 63.670 182.760 63.840 ;
        RECT 181.765 63.525 181.940 63.560 ;
        RECT 181.010 62.990 181.340 63.390 ;
        RECT 181.765 63.160 182.295 63.525 ;
        RECT 182.485 63.160 182.760 63.670 ;
        RECT 182.930 63.160 183.120 64.520 ;
        RECT 183.290 64.535 183.460 65.200 ;
        RECT 183.630 64.780 183.800 65.540 ;
        RECT 184.035 64.780 184.550 65.190 ;
        RECT 183.290 64.345 184.040 64.535 ;
        RECT 184.210 63.970 184.550 64.780 ;
        RECT 185.645 64.740 185.960 65.540 ;
        RECT 186.225 65.200 187.305 65.355 ;
        RECT 186.160 65.185 187.305 65.200 ;
        RECT 186.160 65.030 186.395 65.185 ;
        RECT 186.225 64.570 186.395 65.030 ;
        RECT 183.320 63.800 184.550 63.970 ;
        RECT 183.300 62.990 183.810 63.525 ;
        RECT 184.030 63.195 184.275 63.800 ;
        RECT 185.640 63.560 185.910 64.570 ;
        RECT 186.080 64.400 186.395 64.570 ;
        RECT 186.080 63.730 186.250 64.400 ;
        RECT 186.565 64.230 186.800 64.910 ;
        RECT 186.970 64.400 187.305 65.185 ;
        RECT 187.480 64.450 190.990 65.540 ;
        RECT 191.160 64.450 192.370 65.540 ;
        RECT 192.540 65.030 193.730 65.320 ;
        RECT 186.420 63.900 186.800 64.230 ;
        RECT 186.970 63.900 187.305 64.230 ;
        RECT 187.480 63.760 189.130 64.280 ;
        RECT 189.300 63.930 190.990 64.450 ;
        RECT 186.080 63.560 187.305 63.730 ;
        RECT 185.710 62.990 186.040 63.390 ;
        RECT 186.210 63.290 186.380 63.560 ;
        RECT 186.550 62.990 186.880 63.390 ;
        RECT 187.050 63.290 187.305 63.560 ;
        RECT 187.480 62.990 190.990 63.760 ;
        RECT 191.160 63.740 191.680 64.280 ;
        RECT 191.850 63.910 192.370 64.450 ;
        RECT 192.560 64.690 193.730 64.860 ;
        RECT 193.900 64.740 194.180 65.540 ;
        RECT 192.560 64.400 192.885 64.690 ;
        RECT 193.560 64.570 193.730 64.690 ;
        RECT 193.055 64.230 193.250 64.520 ;
        RECT 193.560 64.400 194.220 64.570 ;
        RECT 194.390 64.400 194.665 65.370 ;
        RECT 194.050 64.230 194.220 64.400 ;
        RECT 192.540 63.900 192.885 64.230 ;
        RECT 193.055 63.900 193.880 64.230 ;
        RECT 194.050 63.900 194.325 64.230 ;
        RECT 191.160 62.990 192.370 63.740 ;
        RECT 194.050 63.730 194.220 63.900 ;
        RECT 192.555 63.560 194.220 63.730 ;
        RECT 194.495 63.665 194.665 64.400 ;
        RECT 194.915 64.570 195.190 65.370 ;
        RECT 195.360 64.740 195.690 65.540 ;
        RECT 195.860 65.200 196.940 65.370 ;
        RECT 195.860 64.570 196.030 65.200 ;
        RECT 194.915 64.360 196.030 64.570 ;
        RECT 196.245 64.520 196.490 65.030 ;
        RECT 196.660 64.700 196.940 65.200 ;
        RECT 197.175 64.700 197.425 65.540 ;
        RECT 197.640 64.520 197.810 65.370 ;
        RECT 197.980 64.780 198.310 65.540 ;
        RECT 198.545 64.570 198.715 64.820 ;
        RECT 196.245 64.350 197.810 64.520 ;
        RECT 198.030 64.400 198.715 64.570 ;
        RECT 198.980 64.450 200.650 65.540 ;
        RECT 194.840 63.980 195.635 64.180 ;
        RECT 195.805 63.980 196.945 64.180 ;
        RECT 197.115 63.810 197.370 64.350 ;
        RECT 198.030 64.150 198.200 64.400 ;
        RECT 197.560 63.980 198.200 64.150 ;
        RECT 192.555 63.210 192.810 63.560 ;
        RECT 192.980 62.990 193.310 63.390 ;
        RECT 193.480 63.210 193.650 63.560 ;
        RECT 193.820 62.990 194.200 63.390 ;
        RECT 194.390 63.320 194.665 63.665 ;
        RECT 194.915 63.630 196.870 63.810 ;
        RECT 194.915 63.170 195.270 63.630 ;
        RECT 195.440 62.990 195.610 63.460 ;
        RECT 195.780 63.160 196.110 63.630 ;
        RECT 196.280 62.990 196.450 63.460 ;
        RECT 196.620 63.380 196.870 63.630 ;
        RECT 197.040 63.550 197.370 63.810 ;
        RECT 197.540 63.380 197.820 63.810 ;
        RECT 196.620 63.160 197.820 63.380 ;
        RECT 198.030 63.730 198.200 63.980 ;
        RECT 198.370 63.900 198.810 64.230 ;
        RECT 198.980 63.760 199.730 64.280 ;
        RECT 199.900 63.930 200.650 64.450 ;
        RECT 200.820 64.375 201.110 65.540 ;
        RECT 201.280 64.400 201.620 65.370 ;
        RECT 201.790 64.400 201.960 65.540 ;
        RECT 202.230 64.740 202.480 65.540 ;
        RECT 203.125 64.570 203.455 65.370 ;
        RECT 203.755 64.740 204.085 65.540 ;
        RECT 204.255 64.570 204.585 65.370 ;
        RECT 202.150 64.400 204.585 64.570 ;
        RECT 204.960 64.450 208.470 65.540 ;
        RECT 201.280 63.790 201.455 64.400 ;
        RECT 202.150 64.150 202.320 64.400 ;
        RECT 201.625 63.980 202.320 64.150 ;
        RECT 202.495 63.980 202.915 64.180 ;
        RECT 203.085 63.980 203.415 64.180 ;
        RECT 203.585 63.980 203.915 64.180 ;
        RECT 198.030 63.350 198.295 63.730 ;
        RECT 198.545 62.990 198.715 63.730 ;
        RECT 198.980 62.990 200.650 63.760 ;
        RECT 200.820 62.990 201.110 63.715 ;
        RECT 201.280 63.160 201.620 63.790 ;
        RECT 201.790 62.990 202.040 63.790 ;
        RECT 202.230 63.640 203.455 63.810 ;
        RECT 202.230 63.160 202.560 63.640 ;
        RECT 202.730 62.990 202.955 63.450 ;
        RECT 203.125 63.160 203.455 63.640 ;
        RECT 204.085 63.770 204.255 64.400 ;
        RECT 204.440 63.980 204.790 64.230 ;
        RECT 204.085 63.160 204.585 63.770 ;
        RECT 204.960 63.760 206.610 64.280 ;
        RECT 206.780 63.930 208.470 64.450 ;
        RECT 208.845 64.570 209.175 65.370 ;
        RECT 209.345 64.740 209.675 65.540 ;
        RECT 209.975 64.570 210.305 65.370 ;
        RECT 210.950 64.740 211.200 65.540 ;
        RECT 208.845 64.400 211.280 64.570 ;
        RECT 211.470 64.400 211.640 65.540 ;
        RECT 211.810 64.400 212.150 65.370 ;
        RECT 212.525 64.570 212.855 65.370 ;
        RECT 213.025 64.740 213.355 65.540 ;
        RECT 213.655 64.570 213.985 65.370 ;
        RECT 214.630 64.740 214.880 65.540 ;
        RECT 212.525 64.400 214.960 64.570 ;
        RECT 215.150 64.400 215.320 65.540 ;
        RECT 215.490 64.400 215.830 65.370 ;
        RECT 216.205 64.570 216.535 65.370 ;
        RECT 216.705 64.740 217.035 65.540 ;
        RECT 217.335 64.570 217.665 65.370 ;
        RECT 218.310 64.740 218.560 65.540 ;
        RECT 216.205 64.400 218.640 64.570 ;
        RECT 218.830 64.400 219.000 65.540 ;
        RECT 219.170 64.400 219.510 65.370 ;
        RECT 208.640 63.980 208.990 64.230 ;
        RECT 209.175 63.770 209.345 64.400 ;
        RECT 209.515 63.980 209.845 64.180 ;
        RECT 210.015 63.980 210.345 64.180 ;
        RECT 210.515 63.980 210.935 64.180 ;
        RECT 211.110 64.150 211.280 64.400 ;
        RECT 211.110 63.980 211.805 64.150 ;
        RECT 204.960 62.990 208.470 63.760 ;
        RECT 208.845 63.160 209.345 63.770 ;
        RECT 209.975 63.640 211.200 63.810 ;
        RECT 211.975 63.790 212.150 64.400 ;
        RECT 212.320 63.980 212.670 64.230 ;
        RECT 209.975 63.160 210.305 63.640 ;
        RECT 210.475 62.990 210.700 63.450 ;
        RECT 210.870 63.160 211.200 63.640 ;
        RECT 211.390 62.990 211.640 63.790 ;
        RECT 211.810 63.160 212.150 63.790 ;
        RECT 212.855 63.770 213.025 64.400 ;
        RECT 213.195 63.980 213.525 64.180 ;
        RECT 213.695 63.980 214.025 64.180 ;
        RECT 214.195 63.980 214.615 64.180 ;
        RECT 214.790 64.150 214.960 64.400 ;
        RECT 214.790 63.980 215.485 64.150 ;
        RECT 212.525 63.160 213.025 63.770 ;
        RECT 213.655 63.640 214.880 63.810 ;
        RECT 215.655 63.790 215.830 64.400 ;
        RECT 216.000 63.980 216.350 64.230 ;
        RECT 213.655 63.160 213.985 63.640 ;
        RECT 214.155 62.990 214.380 63.450 ;
        RECT 214.550 63.160 214.880 63.640 ;
        RECT 215.070 62.990 215.320 63.790 ;
        RECT 215.490 63.160 215.830 63.790 ;
        RECT 216.535 63.770 216.705 64.400 ;
        RECT 216.875 63.980 217.205 64.180 ;
        RECT 217.375 63.980 217.705 64.180 ;
        RECT 217.875 63.980 218.295 64.180 ;
        RECT 218.470 64.150 218.640 64.400 ;
        RECT 218.470 63.980 219.165 64.150 ;
        RECT 216.205 63.160 216.705 63.770 ;
        RECT 217.335 63.640 218.560 63.810 ;
        RECT 219.335 63.790 219.510 64.400 ;
        RECT 217.335 63.160 217.665 63.640 ;
        RECT 217.835 62.990 218.060 63.450 ;
        RECT 218.230 63.160 218.560 63.640 ;
        RECT 218.750 62.990 219.000 63.790 ;
        RECT 219.170 63.160 219.510 63.790 ;
        RECT 219.680 64.820 220.140 65.370 ;
        RECT 220.330 64.820 220.660 65.540 ;
        RECT 219.680 63.450 219.930 64.820 ;
        RECT 220.860 64.650 221.160 65.200 ;
        RECT 221.330 64.870 221.610 65.540 ;
        RECT 220.220 64.480 221.160 64.650 ;
        RECT 220.220 64.230 220.390 64.480 ;
        RECT 221.530 64.230 221.795 64.590 ;
        RECT 221.980 64.450 225.490 65.540 ;
        RECT 220.100 63.900 220.390 64.230 ;
        RECT 220.560 63.980 220.900 64.230 ;
        RECT 221.120 63.980 221.795 64.230 ;
        RECT 220.220 63.810 220.390 63.900 ;
        RECT 220.220 63.620 221.610 63.810 ;
        RECT 219.680 63.160 220.240 63.450 ;
        RECT 220.410 62.990 220.660 63.450 ;
        RECT 221.280 63.260 221.610 63.620 ;
        RECT 221.980 63.760 223.630 64.280 ;
        RECT 223.800 63.930 225.490 64.450 ;
        RECT 226.580 64.375 226.870 65.540 ;
        RECT 227.040 65.105 232.385 65.540 ;
        RECT 232.560 65.105 237.905 65.540 ;
        RECT 221.980 62.990 225.490 63.760 ;
        RECT 226.580 62.990 226.870 63.715 ;
        RECT 228.625 63.535 228.965 64.365 ;
        RECT 230.445 63.855 230.795 65.105 ;
        RECT 234.145 63.535 234.485 64.365 ;
        RECT 235.965 63.855 236.315 65.105 ;
        RECT 238.080 64.450 240.670 65.540 ;
        RECT 238.080 63.760 239.290 64.280 ;
        RECT 239.460 63.930 240.670 64.450 ;
        RECT 240.890 64.525 241.145 65.365 ;
        RECT 241.320 64.720 241.650 65.540 ;
        RECT 241.890 64.550 242.100 65.365 ;
        RECT 227.040 62.990 232.385 63.535 ;
        RECT 232.560 62.990 237.905 63.535 ;
        RECT 238.080 62.990 240.670 63.760 ;
        RECT 240.890 63.160 241.220 64.525 ;
        RECT 241.450 64.370 242.100 64.550 ;
        RECT 241.450 63.730 241.670 64.370 ;
        RECT 242.270 64.195 242.475 65.370 ;
        RECT 242.045 63.955 242.475 64.195 ;
        RECT 242.645 63.955 242.975 65.370 ;
        RECT 243.155 63.900 243.435 65.370 ;
        RECT 243.615 64.570 243.900 65.365 ;
        RECT 244.080 64.740 244.295 65.540 ;
        RECT 244.475 64.570 244.745 65.365 ;
        RECT 243.615 64.400 244.745 64.570 ;
        RECT 244.980 64.570 245.250 65.340 ;
        RECT 245.420 64.760 245.750 65.540 ;
        RECT 245.955 64.935 246.140 65.340 ;
        RECT 246.310 65.115 246.645 65.540 ;
        RECT 246.820 65.105 252.165 65.540 ;
        RECT 245.955 64.760 246.620 64.935 ;
        RECT 244.980 64.400 246.110 64.570 ;
        RECT 243.660 63.900 244.045 64.230 ;
        RECT 244.265 63.930 244.765 64.195 ;
        RECT 243.740 63.750 244.045 63.900 ;
        RECT 241.450 63.560 243.560 63.730 ;
        RECT 241.450 63.555 242.670 63.560 ;
        RECT 241.390 62.990 242.065 63.375 ;
        RECT 242.340 63.165 242.670 63.555 ;
        RECT 242.840 62.990 243.185 63.390 ;
        RECT 243.355 63.165 243.560 63.560 ;
        RECT 243.740 63.190 244.295 63.750 ;
        RECT 244.470 62.990 244.710 63.665 ;
        RECT 244.980 63.490 245.150 64.400 ;
        RECT 245.320 63.650 245.680 64.230 ;
        RECT 245.860 63.900 246.110 64.400 ;
        RECT 246.280 63.730 246.620 64.760 ;
        RECT 245.935 63.560 246.620 63.730 ;
        RECT 244.980 63.160 245.240 63.490 ;
        RECT 245.450 62.990 245.725 63.470 ;
        RECT 245.935 63.160 246.140 63.560 ;
        RECT 248.405 63.535 248.745 64.365 ;
        RECT 250.225 63.855 250.575 65.105 ;
        RECT 252.340 64.375 252.630 65.540 ;
        RECT 252.800 65.105 258.145 65.540 ;
        RECT 258.320 65.105 263.665 65.540 ;
        RECT 263.840 65.105 269.185 65.540 ;
        RECT 246.310 62.990 246.645 63.390 ;
        RECT 246.820 62.990 252.165 63.535 ;
        RECT 252.340 62.990 252.630 63.715 ;
        RECT 254.385 63.535 254.725 64.365 ;
        RECT 256.205 63.855 256.555 65.105 ;
        RECT 259.905 63.535 260.245 64.365 ;
        RECT 261.725 63.855 262.075 65.105 ;
        RECT 265.425 63.535 265.765 64.365 ;
        RECT 267.245 63.855 267.595 65.105 ;
        RECT 270.280 65.035 270.910 65.540 ;
        RECT 270.295 64.500 270.550 64.865 ;
        RECT 270.720 64.860 270.910 65.035 ;
        RECT 271.090 65.030 271.565 65.370 ;
        RECT 270.720 64.670 271.050 64.860 ;
        RECT 271.275 64.500 271.525 64.795 ;
        RECT 271.750 64.695 271.965 65.540 ;
        RECT 272.165 64.700 272.440 65.370 ;
        RECT 270.295 64.330 272.085 64.500 ;
        RECT 272.270 64.350 272.440 64.700 ;
        RECT 272.610 64.530 272.870 65.540 ;
        RECT 273.040 64.450 276.550 65.540 ;
        RECT 276.720 64.450 277.930 65.540 ;
        RECT 270.280 63.670 270.665 64.150 ;
        RECT 252.800 62.990 258.145 63.535 ;
        RECT 258.320 62.990 263.665 63.535 ;
        RECT 263.840 62.990 269.185 63.535 ;
        RECT 270.835 63.475 271.090 64.330 ;
        RECT 270.300 63.210 271.090 63.475 ;
        RECT 271.260 63.655 271.670 64.150 ;
        RECT 271.855 63.900 272.085 64.330 ;
        RECT 272.255 63.830 272.870 64.350 ;
        RECT 271.260 63.210 271.490 63.655 ;
        RECT 272.255 63.620 272.425 63.830 ;
        RECT 273.040 63.760 274.690 64.280 ;
        RECT 274.860 63.930 276.550 64.450 ;
        RECT 271.670 62.990 272.000 63.485 ;
        RECT 272.175 63.160 272.425 63.620 ;
        RECT 272.595 62.990 272.870 63.650 ;
        RECT 273.040 62.990 276.550 63.760 ;
        RECT 276.720 63.740 277.240 64.280 ;
        RECT 277.410 63.910 277.930 64.450 ;
        RECT 278.100 64.375 278.390 65.540 ;
        RECT 278.560 64.450 281.150 65.540 ;
        RECT 278.560 63.760 279.770 64.280 ;
        RECT 279.940 63.930 281.150 64.450 ;
        RECT 281.785 64.400 282.120 65.370 ;
        RECT 282.290 64.400 282.460 65.540 ;
        RECT 282.630 65.200 284.660 65.370 ;
        RECT 276.720 62.990 277.930 63.740 ;
        RECT 278.100 62.990 278.390 63.715 ;
        RECT 278.560 62.990 281.150 63.760 ;
        RECT 281.785 63.730 281.955 64.400 ;
        RECT 282.630 64.230 282.800 65.200 ;
        RECT 282.125 63.900 282.380 64.230 ;
        RECT 282.605 63.900 282.800 64.230 ;
        RECT 282.970 64.860 284.095 65.030 ;
        RECT 282.210 63.730 282.380 63.900 ;
        RECT 282.970 63.730 283.140 64.860 ;
        RECT 281.785 63.160 282.040 63.730 ;
        RECT 282.210 63.560 283.140 63.730 ;
        RECT 283.310 64.520 284.320 64.690 ;
        RECT 283.310 63.720 283.480 64.520 ;
        RECT 283.685 64.180 283.960 64.320 ;
        RECT 283.680 64.010 283.960 64.180 ;
        RECT 282.965 63.525 283.140 63.560 ;
        RECT 282.210 62.990 282.540 63.390 ;
        RECT 282.965 63.160 283.495 63.525 ;
        RECT 283.685 63.160 283.960 64.010 ;
        RECT 284.130 63.160 284.320 64.520 ;
        RECT 284.490 64.535 284.660 65.200 ;
        RECT 284.830 64.780 285.000 65.540 ;
        RECT 285.235 64.780 285.750 65.190 ;
        RECT 284.490 64.345 285.240 64.535 ;
        RECT 285.410 63.970 285.750 64.780 ;
        RECT 284.520 63.800 285.750 63.970 ;
        RECT 285.925 64.400 286.260 65.370 ;
        RECT 286.430 64.400 286.600 65.540 ;
        RECT 286.770 65.200 288.800 65.370 ;
        RECT 284.500 62.990 285.010 63.525 ;
        RECT 285.230 63.195 285.475 63.800 ;
        RECT 285.925 63.730 286.095 64.400 ;
        RECT 286.770 64.230 286.940 65.200 ;
        RECT 286.265 63.900 286.520 64.230 ;
        RECT 286.745 63.900 286.940 64.230 ;
        RECT 287.110 64.860 288.235 65.030 ;
        RECT 286.350 63.730 286.520 63.900 ;
        RECT 287.110 63.730 287.280 64.860 ;
        RECT 285.925 63.160 286.180 63.730 ;
        RECT 286.350 63.560 287.280 63.730 ;
        RECT 287.450 64.520 288.460 64.690 ;
        RECT 287.450 63.720 287.620 64.520 ;
        RECT 287.105 63.525 287.280 63.560 ;
        RECT 286.350 62.990 286.680 63.390 ;
        RECT 287.105 63.160 287.635 63.525 ;
        RECT 287.825 63.500 288.100 64.320 ;
        RECT 287.820 63.330 288.100 63.500 ;
        RECT 287.825 63.160 288.100 63.330 ;
        RECT 288.270 63.160 288.460 64.520 ;
        RECT 288.630 64.535 288.800 65.200 ;
        RECT 288.970 64.780 289.140 65.540 ;
        RECT 289.375 64.780 289.890 65.190 ;
        RECT 288.630 64.345 289.380 64.535 ;
        RECT 289.550 63.970 289.890 64.780 ;
        RECT 290.060 64.450 293.570 65.540 ;
        RECT 294.205 64.870 294.460 65.370 ;
        RECT 294.630 65.040 294.960 65.540 ;
        RECT 294.205 64.700 294.955 64.870 ;
        RECT 288.660 63.800 289.890 63.970 ;
        RECT 288.640 62.990 289.150 63.525 ;
        RECT 289.370 63.195 289.615 63.800 ;
        RECT 290.060 63.760 291.710 64.280 ;
        RECT 291.880 63.930 293.570 64.450 ;
        RECT 294.205 63.880 294.555 64.530 ;
        RECT 290.060 62.990 293.570 63.760 ;
        RECT 294.725 63.710 294.955 64.700 ;
        RECT 294.205 63.540 294.955 63.710 ;
        RECT 294.205 63.250 294.460 63.540 ;
        RECT 294.630 62.990 294.960 63.370 ;
        RECT 295.130 63.250 295.300 65.370 ;
        RECT 295.470 64.570 295.795 65.355 ;
        RECT 295.965 65.080 296.215 65.540 ;
        RECT 296.385 65.040 296.635 65.370 ;
        RECT 296.850 65.040 297.530 65.370 ;
        RECT 296.385 64.910 296.555 65.040 ;
        RECT 296.160 64.740 296.555 64.910 ;
        RECT 295.530 63.520 295.990 64.570 ;
        RECT 296.160 63.380 296.330 64.740 ;
        RECT 296.725 64.480 297.190 64.870 ;
        RECT 296.500 63.670 296.850 64.290 ;
        RECT 297.020 63.890 297.190 64.480 ;
        RECT 297.360 64.260 297.530 65.040 ;
        RECT 297.700 64.940 297.870 65.280 ;
        RECT 298.105 65.110 298.435 65.540 ;
        RECT 298.605 64.940 298.775 65.280 ;
        RECT 299.070 65.080 299.440 65.540 ;
        RECT 297.700 64.770 298.775 64.940 ;
        RECT 299.610 64.910 299.780 65.370 ;
        RECT 300.015 65.030 300.885 65.370 ;
        RECT 301.055 65.080 301.305 65.540 ;
        RECT 299.220 64.740 299.780 64.910 ;
        RECT 299.220 64.600 299.390 64.740 ;
        RECT 297.890 64.430 299.390 64.600 ;
        RECT 300.085 64.570 300.545 64.860 ;
        RECT 297.360 64.090 299.050 64.260 ;
        RECT 297.020 63.670 297.375 63.890 ;
        RECT 297.545 63.380 297.715 64.090 ;
        RECT 297.920 63.670 298.710 63.920 ;
        RECT 298.880 63.910 299.050 64.090 ;
        RECT 299.220 63.740 299.390 64.430 ;
        RECT 295.660 62.990 295.990 63.350 ;
        RECT 296.160 63.210 296.655 63.380 ;
        RECT 296.860 63.210 297.715 63.380 ;
        RECT 298.590 62.990 298.920 63.450 ;
        RECT 299.130 63.350 299.390 63.740 ;
        RECT 299.580 64.560 300.545 64.570 ;
        RECT 300.715 64.650 300.885 65.030 ;
        RECT 301.475 64.990 301.645 65.280 ;
        RECT 301.825 65.160 302.155 65.540 ;
        RECT 301.475 64.820 302.275 64.990 ;
        RECT 299.580 64.400 300.255 64.560 ;
        RECT 300.715 64.480 301.935 64.650 ;
        RECT 299.580 63.610 299.790 64.400 ;
        RECT 300.715 64.390 300.885 64.480 ;
        RECT 299.960 63.610 300.310 64.230 ;
        RECT 300.480 64.220 300.885 64.390 ;
        RECT 300.480 63.440 300.650 64.220 ;
        RECT 300.820 63.770 301.040 64.050 ;
        RECT 301.220 63.940 301.760 64.310 ;
        RECT 302.105 64.230 302.275 64.820 ;
        RECT 302.495 64.400 302.800 65.540 ;
        RECT 302.970 64.350 303.220 65.230 ;
        RECT 303.390 64.400 303.640 65.540 ;
        RECT 303.860 64.375 304.150 65.540 ;
        RECT 304.320 65.105 309.665 65.540 ;
        RECT 302.105 64.200 302.845 64.230 ;
        RECT 300.820 63.600 301.350 63.770 ;
        RECT 299.130 63.180 299.480 63.350 ;
        RECT 299.700 63.160 300.650 63.440 ;
        RECT 300.820 62.990 301.010 63.430 ;
        RECT 301.180 63.370 301.350 63.600 ;
        RECT 301.520 63.540 301.760 63.940 ;
        RECT 301.930 63.900 302.845 64.200 ;
        RECT 301.930 63.725 302.255 63.900 ;
        RECT 301.930 63.370 302.250 63.725 ;
        RECT 303.015 63.700 303.220 64.350 ;
        RECT 301.180 63.200 302.250 63.370 ;
        RECT 302.495 62.990 302.800 63.450 ;
        RECT 302.970 63.170 303.220 63.700 ;
        RECT 303.390 62.990 303.640 63.745 ;
        RECT 303.860 62.990 304.150 63.715 ;
        RECT 305.905 63.535 306.245 64.365 ;
        RECT 307.725 63.855 308.075 65.105 ;
        RECT 309.840 64.450 311.050 65.540 ;
        RECT 309.840 63.910 310.360 64.450 ;
        RECT 310.530 63.740 311.050 64.280 ;
        RECT 304.320 62.990 309.665 63.535 ;
        RECT 309.840 62.990 311.050 63.740 ;
        RECT 162.095 62.820 311.135 62.990 ;
        RECT 162.180 62.070 163.390 62.820 ;
        RECT 162.180 61.530 162.700 62.070 ;
        RECT 163.565 61.980 163.825 62.820 ;
        RECT 164.000 62.075 164.255 62.650 ;
        RECT 164.425 62.440 164.755 62.820 ;
        RECT 164.970 62.270 165.140 62.650 ;
        RECT 164.425 62.100 165.140 62.270 ;
        RECT 162.870 61.360 163.390 61.900 ;
        RECT 162.180 60.270 163.390 61.360 ;
        RECT 163.565 60.270 163.825 61.420 ;
        RECT 164.000 61.345 164.170 62.075 ;
        RECT 164.425 61.910 164.595 62.100 ;
        RECT 165.400 62.050 168.910 62.820 ;
        RECT 169.130 62.065 169.380 62.820 ;
        RECT 169.550 62.110 169.800 62.640 ;
        RECT 169.970 62.360 170.275 62.820 ;
        RECT 170.520 62.440 171.590 62.610 ;
        RECT 164.340 61.580 164.595 61.910 ;
        RECT 164.425 61.370 164.595 61.580 ;
        RECT 164.875 61.550 165.230 61.920 ;
        RECT 165.400 61.530 167.050 62.050 ;
        RECT 164.000 60.440 164.255 61.345 ;
        RECT 164.425 61.200 165.140 61.370 ;
        RECT 167.220 61.360 168.910 61.880 ;
        RECT 169.550 61.460 169.755 62.110 ;
        RECT 170.520 62.085 170.840 62.440 ;
        RECT 170.515 61.910 170.840 62.085 ;
        RECT 169.925 61.610 170.840 61.910 ;
        RECT 171.010 61.870 171.250 62.270 ;
        RECT 171.420 62.210 171.590 62.440 ;
        RECT 171.760 62.380 171.950 62.820 ;
        RECT 172.120 62.370 173.070 62.650 ;
        RECT 173.290 62.460 173.640 62.630 ;
        RECT 171.420 62.040 171.950 62.210 ;
        RECT 169.925 61.580 170.665 61.610 ;
        RECT 164.425 60.270 164.755 61.030 ;
        RECT 164.970 60.440 165.140 61.200 ;
        RECT 165.400 60.270 168.910 61.360 ;
        RECT 169.130 60.270 169.380 61.410 ;
        RECT 169.550 60.580 169.800 61.460 ;
        RECT 169.970 60.270 170.275 61.410 ;
        RECT 170.495 60.990 170.665 61.580 ;
        RECT 171.010 61.500 171.550 61.870 ;
        RECT 171.730 61.760 171.950 62.040 ;
        RECT 172.120 61.590 172.290 62.370 ;
        RECT 171.885 61.420 172.290 61.590 ;
        RECT 172.460 61.580 172.810 62.200 ;
        RECT 171.885 61.330 172.055 61.420 ;
        RECT 172.980 61.410 173.190 62.200 ;
        RECT 170.835 61.160 172.055 61.330 ;
        RECT 172.515 61.250 173.190 61.410 ;
        RECT 170.495 60.820 171.295 60.990 ;
        RECT 170.615 60.270 170.945 60.650 ;
        RECT 171.125 60.530 171.295 60.820 ;
        RECT 171.885 60.780 172.055 61.160 ;
        RECT 172.225 61.240 173.190 61.250 ;
        RECT 173.380 62.070 173.640 62.460 ;
        RECT 173.850 62.360 174.180 62.820 ;
        RECT 175.055 62.430 175.910 62.600 ;
        RECT 176.115 62.430 176.610 62.600 ;
        RECT 176.780 62.460 177.110 62.820 ;
        RECT 173.380 61.380 173.550 62.070 ;
        RECT 173.720 61.720 173.890 61.900 ;
        RECT 174.060 61.890 174.850 62.140 ;
        RECT 175.055 61.720 175.225 62.430 ;
        RECT 175.395 61.920 175.750 62.140 ;
        RECT 173.720 61.550 175.410 61.720 ;
        RECT 172.225 60.950 172.685 61.240 ;
        RECT 173.380 61.210 174.880 61.380 ;
        RECT 173.380 61.070 173.550 61.210 ;
        RECT 172.990 60.900 173.550 61.070 ;
        RECT 171.465 60.270 171.715 60.730 ;
        RECT 171.885 60.440 172.755 60.780 ;
        RECT 172.990 60.440 173.160 60.900 ;
        RECT 173.995 60.870 175.070 61.040 ;
        RECT 173.330 60.270 173.700 60.730 ;
        RECT 173.995 60.530 174.165 60.870 ;
        RECT 174.335 60.270 174.665 60.700 ;
        RECT 174.900 60.530 175.070 60.870 ;
        RECT 175.240 60.770 175.410 61.550 ;
        RECT 175.580 61.330 175.750 61.920 ;
        RECT 175.920 61.520 176.270 62.140 ;
        RECT 175.580 60.940 176.045 61.330 ;
        RECT 176.440 61.070 176.610 62.430 ;
        RECT 176.780 61.240 177.240 62.290 ;
        RECT 176.215 60.900 176.610 61.070 ;
        RECT 176.215 60.770 176.385 60.900 ;
        RECT 175.240 60.440 175.920 60.770 ;
        RECT 176.135 60.440 176.385 60.770 ;
        RECT 176.555 60.270 176.805 60.730 ;
        RECT 176.975 60.455 177.300 61.240 ;
        RECT 177.470 60.440 177.640 62.560 ;
        RECT 177.810 62.440 178.140 62.820 ;
        RECT 178.310 62.270 178.565 62.560 ;
        RECT 177.815 62.100 178.565 62.270 ;
        RECT 177.815 61.110 178.045 62.100 ;
        RECT 178.740 62.020 179.030 62.820 ;
        RECT 179.200 62.360 179.750 62.650 ;
        RECT 179.920 62.360 180.170 62.820 ;
        RECT 178.215 61.280 178.565 61.930 ;
        RECT 177.815 60.940 178.565 61.110 ;
        RECT 177.810 60.270 178.140 60.770 ;
        RECT 178.310 60.440 178.565 60.940 ;
        RECT 178.740 60.270 179.030 61.410 ;
        RECT 179.200 60.990 179.450 62.360 ;
        RECT 180.800 62.190 181.130 62.550 ;
        RECT 179.740 62.000 181.130 62.190 ;
        RECT 181.500 62.050 185.010 62.820 ;
        RECT 179.740 61.910 179.910 62.000 ;
        RECT 179.620 61.580 179.910 61.910 ;
        RECT 180.080 61.580 180.410 61.830 ;
        RECT 180.640 61.580 181.330 61.830 ;
        RECT 179.740 61.330 179.910 61.580 ;
        RECT 179.740 61.160 180.680 61.330 ;
        RECT 179.200 60.440 179.650 60.990 ;
        RECT 179.840 60.270 180.170 60.990 ;
        RECT 180.380 60.610 180.680 61.160 ;
        RECT 181.015 61.140 181.330 61.580 ;
        RECT 181.500 61.530 183.150 62.050 ;
        RECT 185.180 62.020 185.470 62.820 ;
        RECT 185.640 62.360 186.190 62.650 ;
        RECT 186.360 62.360 186.610 62.820 ;
        RECT 183.320 61.360 185.010 61.880 ;
        RECT 180.850 60.270 181.130 60.940 ;
        RECT 181.500 60.270 185.010 61.360 ;
        RECT 185.180 60.270 185.470 61.410 ;
        RECT 185.640 60.990 185.890 62.360 ;
        RECT 187.240 62.190 187.570 62.550 ;
        RECT 186.180 62.000 187.570 62.190 ;
        RECT 187.940 62.095 188.230 62.820 ;
        RECT 188.860 62.440 189.190 62.820 ;
        RECT 188.415 62.270 188.690 62.410 ;
        RECT 189.360 62.270 189.570 62.440 ;
        RECT 188.415 62.080 189.570 62.270 ;
        RECT 189.740 62.270 190.070 62.650 ;
        RECT 190.260 62.440 190.590 62.820 ;
        RECT 189.740 62.065 190.590 62.270 ;
        RECT 186.180 61.910 186.350 62.000 ;
        RECT 186.060 61.580 186.350 61.910 ;
        RECT 186.520 61.580 186.850 61.830 ;
        RECT 187.080 61.580 187.770 61.830 ;
        RECT 186.180 61.330 186.350 61.580 ;
        RECT 186.180 61.160 187.120 61.330 ;
        RECT 185.640 60.440 186.090 60.990 ;
        RECT 186.280 60.270 186.610 60.990 ;
        RECT 186.820 60.610 187.120 61.160 ;
        RECT 187.455 61.140 187.770 61.580 ;
        RECT 188.410 61.455 188.670 61.910 ;
        RECT 188.925 61.505 189.510 61.880 ;
        RECT 187.290 60.270 187.570 60.940 ;
        RECT 187.940 60.270 188.230 61.435 ;
        RECT 188.415 60.270 188.740 61.255 ;
        RECT 188.925 61.120 189.130 61.505 ;
        RECT 189.680 61.290 190.090 61.895 ;
        RECT 190.260 61.575 190.590 62.065 ;
        RECT 190.260 61.120 190.430 61.575 ;
        RECT 188.920 60.950 189.130 61.120 ;
        RECT 188.925 60.920 189.130 60.950 ;
        RECT 189.310 60.900 190.430 61.120 ;
        RECT 189.310 60.440 189.570 60.900 ;
        RECT 189.740 60.270 190.590 60.720 ;
        RECT 190.760 60.440 191.005 62.650 ;
        RECT 191.190 62.020 191.430 62.820 ;
        RECT 191.620 62.145 191.880 62.650 ;
        RECT 192.060 62.440 192.390 62.820 ;
        RECT 192.570 62.270 192.740 62.650 ;
        RECT 193.010 62.315 193.340 62.820 ;
        RECT 191.620 61.345 191.800 62.145 ;
        RECT 192.075 62.100 192.740 62.270 ;
        RECT 193.510 62.250 193.750 62.625 ;
        RECT 194.030 62.490 194.200 62.635 ;
        RECT 194.030 62.295 194.430 62.490 ;
        RECT 194.790 62.325 195.190 62.820 ;
        RECT 192.075 61.845 192.245 62.100 ;
        RECT 191.970 61.515 192.245 61.845 ;
        RECT 192.470 61.550 192.810 61.920 ;
        RECT 192.075 61.370 192.245 61.515 ;
        RECT 193.065 61.460 193.365 62.140 ;
        RECT 191.190 60.270 191.445 61.270 ;
        RECT 191.620 60.440 191.890 61.345 ;
        RECT 192.075 61.200 192.750 61.370 ;
        RECT 193.060 61.290 193.365 61.460 ;
        RECT 193.535 62.100 193.750 62.250 ;
        RECT 193.535 61.770 194.090 62.100 ;
        RECT 194.260 61.960 194.430 62.295 ;
        RECT 195.360 62.130 195.595 62.650 ;
        RECT 195.780 62.185 196.050 62.820 ;
        RECT 192.060 60.270 192.390 61.030 ;
        RECT 192.570 60.440 192.750 61.200 ;
        RECT 193.535 61.120 193.770 61.770 ;
        RECT 194.260 61.600 195.250 61.960 ;
        RECT 193.090 60.890 193.770 61.120 ;
        RECT 193.960 61.580 195.250 61.600 ;
        RECT 193.960 61.430 194.820 61.580 ;
        RECT 193.090 60.460 193.260 60.890 ;
        RECT 193.430 60.270 193.760 60.720 ;
        RECT 193.960 60.485 194.245 61.430 ;
        RECT 195.420 61.325 195.595 62.130 ;
        RECT 194.420 60.950 195.115 61.260 ;
        RECT 194.425 60.270 195.110 60.740 ;
        RECT 195.290 60.540 195.595 61.325 ;
        RECT 196.680 62.020 197.020 62.650 ;
        RECT 197.310 62.360 197.480 62.820 ;
        RECT 197.750 62.190 198.080 62.635 ;
        RECT 196.680 61.450 196.950 62.020 ;
        RECT 197.330 62.000 198.080 62.190 ;
        RECT 198.250 62.170 198.420 62.490 ;
        RECT 198.645 62.360 198.975 62.820 ;
        RECT 199.175 62.170 199.505 62.650 ;
        RECT 199.720 62.360 200.050 62.820 ;
        RECT 200.220 62.170 200.550 62.650 ;
        RECT 200.820 62.275 206.165 62.820 ;
        RECT 198.250 62.000 200.550 62.170 ;
        RECT 197.330 61.830 197.700 62.000 ;
        RECT 197.120 61.620 197.700 61.830 ;
        RECT 197.870 61.620 198.290 61.830 ;
        RECT 197.440 61.450 197.700 61.620 ;
        RECT 195.780 60.270 196.050 61.225 ;
        RECT 196.680 60.440 197.205 61.450 ;
        RECT 197.440 61.160 198.190 61.450 ;
        RECT 197.440 60.270 197.770 60.990 ;
        RECT 197.940 60.440 198.190 61.160 ;
        RECT 198.460 60.515 198.790 61.830 ;
        RECT 199.000 60.515 199.330 61.830 ;
        RECT 199.500 60.515 199.870 61.830 ;
        RECT 200.080 61.580 200.590 61.830 ;
        RECT 202.405 61.445 202.745 62.275 ;
        RECT 206.340 62.050 208.010 62.820 ;
        RECT 200.200 60.270 200.530 61.390 ;
        RECT 204.225 60.705 204.575 61.955 ;
        RECT 206.340 61.530 207.090 62.050 ;
        RECT 208.640 62.020 208.980 62.650 ;
        RECT 209.270 62.360 209.440 62.820 ;
        RECT 209.710 62.190 210.040 62.635 ;
        RECT 207.260 61.360 208.010 61.880 ;
        RECT 200.820 60.270 206.165 60.705 ;
        RECT 206.340 60.270 208.010 61.360 ;
        RECT 208.640 61.450 208.910 62.020 ;
        RECT 209.290 62.000 210.040 62.190 ;
        RECT 210.210 62.170 210.380 62.490 ;
        RECT 210.605 62.360 210.935 62.820 ;
        RECT 211.135 62.170 211.465 62.650 ;
        RECT 211.680 62.360 212.010 62.820 ;
        RECT 212.180 62.170 212.510 62.650 ;
        RECT 210.210 62.000 212.510 62.170 ;
        RECT 213.700 62.095 213.990 62.820 ;
        RECT 214.160 62.020 214.500 62.650 ;
        RECT 214.790 62.360 214.960 62.820 ;
        RECT 215.230 62.190 215.560 62.635 ;
        RECT 209.290 61.830 209.660 62.000 ;
        RECT 209.080 61.620 209.660 61.830 ;
        RECT 209.830 61.620 210.250 61.830 ;
        RECT 209.400 61.450 209.660 61.620 ;
        RECT 208.640 60.440 209.165 61.450 ;
        RECT 209.400 61.160 210.150 61.450 ;
        RECT 209.400 60.270 209.730 60.990 ;
        RECT 209.900 60.440 210.150 61.160 ;
        RECT 210.420 60.515 210.750 61.830 ;
        RECT 210.960 60.515 211.290 61.830 ;
        RECT 211.460 60.515 211.830 61.830 ;
        RECT 212.040 61.580 212.550 61.830 ;
        RECT 214.160 61.450 214.430 62.020 ;
        RECT 214.810 62.000 215.560 62.190 ;
        RECT 215.730 62.170 215.900 62.490 ;
        RECT 216.125 62.360 216.455 62.820 ;
        RECT 216.655 62.170 216.985 62.650 ;
        RECT 217.200 62.360 217.530 62.820 ;
        RECT 217.700 62.170 218.030 62.650 ;
        RECT 215.730 62.000 218.030 62.170 ;
        RECT 218.300 62.050 219.970 62.820 ;
        RECT 220.140 62.080 220.580 62.640 ;
        RECT 220.750 62.080 221.200 62.820 ;
        RECT 221.370 62.250 221.540 62.650 ;
        RECT 221.710 62.420 222.130 62.820 ;
        RECT 222.300 62.250 222.530 62.650 ;
        RECT 221.370 62.080 222.530 62.250 ;
        RECT 222.700 62.080 223.190 62.650 ;
        RECT 214.810 61.830 215.180 62.000 ;
        RECT 214.600 61.620 215.180 61.830 ;
        RECT 215.350 61.620 215.770 61.830 ;
        RECT 214.920 61.450 215.180 61.620 ;
        RECT 212.160 60.270 212.490 61.390 ;
        RECT 213.700 60.270 213.990 61.435 ;
        RECT 214.160 60.440 214.685 61.450 ;
        RECT 214.920 61.160 215.670 61.450 ;
        RECT 214.920 60.270 215.250 60.990 ;
        RECT 215.420 60.440 215.670 61.160 ;
        RECT 215.940 60.515 216.270 61.830 ;
        RECT 216.480 60.515 216.810 61.830 ;
        RECT 216.980 60.515 217.350 61.830 ;
        RECT 217.560 61.580 218.070 61.830 ;
        RECT 218.300 61.530 219.050 62.050 ;
        RECT 217.680 60.270 218.010 61.390 ;
        RECT 219.220 61.360 219.970 61.880 ;
        RECT 218.300 60.270 219.970 61.360 ;
        RECT 220.140 61.070 220.450 62.080 ;
        RECT 220.620 61.460 220.790 61.910 ;
        RECT 220.960 61.630 221.350 61.910 ;
        RECT 221.535 61.580 221.780 61.910 ;
        RECT 220.620 61.290 221.410 61.460 ;
        RECT 220.140 60.440 220.580 61.070 ;
        RECT 220.755 60.270 221.070 61.120 ;
        RECT 221.240 60.610 221.410 61.290 ;
        RECT 221.580 60.780 221.780 61.580 ;
        RECT 221.980 60.780 222.230 61.910 ;
        RECT 222.445 61.580 222.850 61.910 ;
        RECT 223.020 61.410 223.190 62.080 ;
        RECT 222.420 61.240 223.190 61.410 ;
        RECT 223.820 62.080 224.205 62.650 ;
        RECT 224.375 62.360 224.700 62.820 ;
        RECT 225.220 62.190 225.500 62.650 ;
        RECT 223.820 61.410 224.100 62.080 ;
        RECT 224.375 62.020 225.500 62.190 ;
        RECT 224.375 61.910 224.825 62.020 ;
        RECT 224.270 61.580 224.825 61.910 ;
        RECT 225.690 61.850 226.090 62.650 ;
        RECT 226.490 62.360 226.760 62.820 ;
        RECT 226.930 62.190 227.215 62.650 ;
        RECT 222.420 60.610 222.670 61.240 ;
        RECT 221.240 60.440 222.670 60.610 ;
        RECT 222.850 60.270 223.180 61.070 ;
        RECT 223.820 60.440 224.205 61.410 ;
        RECT 224.375 61.120 224.825 61.580 ;
        RECT 224.995 61.290 226.090 61.850 ;
        RECT 224.375 60.900 225.500 61.120 ;
        RECT 224.375 60.270 224.700 60.730 ;
        RECT 225.220 60.440 225.500 60.900 ;
        RECT 225.690 60.440 226.090 61.290 ;
        RECT 226.260 62.020 227.215 62.190 ;
        RECT 227.500 62.050 230.090 62.820 ;
        RECT 230.265 62.080 230.520 62.650 ;
        RECT 230.690 62.420 231.020 62.820 ;
        RECT 231.445 62.285 231.975 62.650 ;
        RECT 231.445 62.250 231.620 62.285 ;
        RECT 230.690 62.080 231.620 62.250 ;
        RECT 226.260 61.120 226.470 62.020 ;
        RECT 226.640 61.290 227.330 61.850 ;
        RECT 227.500 61.530 228.710 62.050 ;
        RECT 228.880 61.360 230.090 61.880 ;
        RECT 226.260 60.900 227.215 61.120 ;
        RECT 226.490 60.270 226.760 60.730 ;
        RECT 226.930 60.440 227.215 60.900 ;
        RECT 227.500 60.270 230.090 61.360 ;
        RECT 230.265 61.410 230.435 62.080 ;
        RECT 230.690 61.910 230.860 62.080 ;
        RECT 230.605 61.580 230.860 61.910 ;
        RECT 231.085 61.580 231.280 61.910 ;
        RECT 230.265 60.440 230.600 61.410 ;
        RECT 230.770 60.270 230.940 61.410 ;
        RECT 231.110 60.610 231.280 61.580 ;
        RECT 231.450 60.950 231.620 62.080 ;
        RECT 231.790 61.290 231.960 62.090 ;
        RECT 232.165 61.800 232.440 62.650 ;
        RECT 232.160 61.630 232.440 61.800 ;
        RECT 232.165 61.490 232.440 61.630 ;
        RECT 232.610 61.290 232.800 62.650 ;
        RECT 232.980 62.285 233.490 62.820 ;
        RECT 233.710 62.010 233.955 62.615 ;
        RECT 234.405 62.080 234.660 62.650 ;
        RECT 234.830 62.420 235.160 62.820 ;
        RECT 235.585 62.285 236.115 62.650 ;
        RECT 235.585 62.250 235.760 62.285 ;
        RECT 234.830 62.080 235.760 62.250 ;
        RECT 233.000 61.840 234.230 62.010 ;
        RECT 231.790 61.120 232.800 61.290 ;
        RECT 232.970 61.275 233.720 61.465 ;
        RECT 231.450 60.780 232.575 60.950 ;
        RECT 232.970 60.610 233.140 61.275 ;
        RECT 233.890 61.030 234.230 61.840 ;
        RECT 231.110 60.440 233.140 60.610 ;
        RECT 233.310 60.270 233.480 61.030 ;
        RECT 233.715 60.620 234.230 61.030 ;
        RECT 234.405 61.410 234.575 62.080 ;
        RECT 234.830 61.910 235.000 62.080 ;
        RECT 234.745 61.580 235.000 61.910 ;
        RECT 235.225 61.580 235.420 61.910 ;
        RECT 234.405 60.440 234.740 61.410 ;
        RECT 234.910 60.270 235.080 61.410 ;
        RECT 235.250 60.610 235.420 61.580 ;
        RECT 235.590 60.950 235.760 62.080 ;
        RECT 235.930 61.290 236.100 62.090 ;
        RECT 236.305 61.800 236.580 62.650 ;
        RECT 236.300 61.630 236.580 61.800 ;
        RECT 236.305 61.490 236.580 61.630 ;
        RECT 236.750 61.290 236.940 62.650 ;
        RECT 237.120 62.285 237.630 62.820 ;
        RECT 237.850 62.010 238.095 62.615 ;
        RECT 239.460 62.095 239.750 62.820 ;
        RECT 239.920 62.080 240.305 62.650 ;
        RECT 240.475 62.360 240.800 62.820 ;
        RECT 241.320 62.190 241.600 62.650 ;
        RECT 237.140 61.840 238.370 62.010 ;
        RECT 235.930 61.120 236.940 61.290 ;
        RECT 237.110 61.275 237.860 61.465 ;
        RECT 235.590 60.780 236.715 60.950 ;
        RECT 237.110 60.610 237.280 61.275 ;
        RECT 238.030 61.030 238.370 61.840 ;
        RECT 235.250 60.440 237.280 60.610 ;
        RECT 237.450 60.270 237.620 61.030 ;
        RECT 237.855 60.620 238.370 61.030 ;
        RECT 239.460 60.270 239.750 61.435 ;
        RECT 239.920 61.410 240.200 62.080 ;
        RECT 240.475 62.020 241.600 62.190 ;
        RECT 240.475 61.910 240.925 62.020 ;
        RECT 240.370 61.580 240.925 61.910 ;
        RECT 241.790 61.850 242.190 62.650 ;
        RECT 242.590 62.360 242.860 62.820 ;
        RECT 243.030 62.190 243.315 62.650 ;
        RECT 243.605 62.565 243.940 62.610 ;
        RECT 239.920 60.440 240.305 61.410 ;
        RECT 240.475 61.120 240.925 61.580 ;
        RECT 241.095 61.290 242.190 61.850 ;
        RECT 240.475 60.900 241.600 61.120 ;
        RECT 240.475 60.270 240.800 60.730 ;
        RECT 241.320 60.440 241.600 60.900 ;
        RECT 241.790 60.440 242.190 61.290 ;
        RECT 242.360 62.020 243.315 62.190 ;
        RECT 243.600 62.100 243.940 62.565 ;
        RECT 244.110 62.440 244.440 62.820 ;
        RECT 242.360 61.120 242.570 62.020 ;
        RECT 242.740 61.290 243.430 61.850 ;
        RECT 243.600 61.410 243.770 62.100 ;
        RECT 243.940 61.580 244.200 61.910 ;
        RECT 242.360 60.900 243.315 61.120 ;
        RECT 242.590 60.270 242.860 60.730 ;
        RECT 243.030 60.440 243.315 60.900 ;
        RECT 243.600 60.440 243.860 61.410 ;
        RECT 244.030 61.030 244.200 61.580 ;
        RECT 244.370 61.210 244.710 62.240 ;
        RECT 244.900 61.460 245.170 62.485 ;
        RECT 244.900 61.290 245.210 61.460 ;
        RECT 244.900 61.210 245.170 61.290 ;
        RECT 245.395 61.210 245.675 62.485 ;
        RECT 245.875 62.320 246.105 62.650 ;
        RECT 246.350 62.440 246.680 62.820 ;
        RECT 245.875 61.030 246.045 62.320 ;
        RECT 246.850 62.250 247.025 62.650 ;
        RECT 246.395 62.080 247.025 62.250 ;
        RECT 247.370 62.270 247.540 62.650 ;
        RECT 247.720 62.440 248.050 62.820 ;
        RECT 247.370 62.100 248.035 62.270 ;
        RECT 248.230 62.145 248.490 62.650 ;
        RECT 246.395 61.910 246.565 62.080 ;
        RECT 246.215 61.580 246.565 61.910 ;
        RECT 244.030 60.860 246.045 61.030 ;
        RECT 246.395 61.060 246.565 61.580 ;
        RECT 246.745 61.230 247.110 61.910 ;
        RECT 247.300 61.550 247.640 61.920 ;
        RECT 247.865 61.845 248.035 62.100 ;
        RECT 247.865 61.515 248.140 61.845 ;
        RECT 247.865 61.370 248.035 61.515 ;
        RECT 247.360 61.200 248.035 61.370 ;
        RECT 248.310 61.345 248.490 62.145 ;
        RECT 248.660 62.190 249.000 62.650 ;
        RECT 249.170 62.360 249.340 62.820 ;
        RECT 249.970 62.385 250.330 62.650 ;
        RECT 249.975 62.380 250.330 62.385 ;
        RECT 249.980 62.370 250.330 62.380 ;
        RECT 249.985 62.365 250.330 62.370 ;
        RECT 249.990 62.355 250.330 62.365 ;
        RECT 250.570 62.360 250.740 62.820 ;
        RECT 249.995 62.350 250.330 62.355 ;
        RECT 250.005 62.340 250.330 62.350 ;
        RECT 250.015 62.330 250.330 62.340 ;
        RECT 249.510 62.190 249.840 62.270 ;
        RECT 248.660 62.000 249.840 62.190 ;
        RECT 250.030 62.190 250.330 62.330 ;
        RECT 250.030 62.000 250.740 62.190 ;
        RECT 246.395 60.890 247.025 61.060 ;
        RECT 244.055 60.270 244.385 60.680 ;
        RECT 244.585 60.440 244.755 60.860 ;
        RECT 244.970 60.270 245.640 60.680 ;
        RECT 245.875 60.440 246.045 60.860 ;
        RECT 246.350 60.270 246.680 60.710 ;
        RECT 246.850 60.440 247.025 60.890 ;
        RECT 247.360 60.440 247.540 61.200 ;
        RECT 247.720 60.270 248.050 61.030 ;
        RECT 248.220 60.440 248.490 61.345 ;
        RECT 248.660 61.630 248.990 61.830 ;
        RECT 249.300 61.810 249.630 61.830 ;
        RECT 249.180 61.630 249.630 61.810 ;
        RECT 248.660 61.290 248.890 61.630 ;
        RECT 248.670 60.270 249.000 60.990 ;
        RECT 249.180 60.515 249.395 61.630 ;
        RECT 249.800 61.600 250.270 61.830 ;
        RECT 250.455 61.430 250.740 62.000 ;
        RECT 250.910 61.875 251.250 62.650 ;
        RECT 249.590 61.215 250.740 61.430 ;
        RECT 249.590 60.440 249.920 61.215 ;
        RECT 250.090 60.270 250.800 61.045 ;
        RECT 250.970 60.440 251.250 61.875 ;
        RECT 251.425 62.080 251.680 62.650 ;
        RECT 251.850 62.420 252.180 62.820 ;
        RECT 252.605 62.285 253.135 62.650 ;
        RECT 253.325 62.480 253.600 62.650 ;
        RECT 253.320 62.310 253.600 62.480 ;
        RECT 252.605 62.250 252.780 62.285 ;
        RECT 251.850 62.080 252.780 62.250 ;
        RECT 251.425 61.410 251.595 62.080 ;
        RECT 251.850 61.910 252.020 62.080 ;
        RECT 251.765 61.580 252.020 61.910 ;
        RECT 252.245 61.580 252.440 61.910 ;
        RECT 251.425 60.440 251.760 61.410 ;
        RECT 251.930 60.270 252.100 61.410 ;
        RECT 252.270 60.610 252.440 61.580 ;
        RECT 252.610 60.950 252.780 62.080 ;
        RECT 252.950 61.290 253.120 62.090 ;
        RECT 253.325 61.490 253.600 62.310 ;
        RECT 253.770 61.290 253.960 62.650 ;
        RECT 254.140 62.285 254.650 62.820 ;
        RECT 254.870 62.010 255.115 62.615 ;
        RECT 255.560 62.050 257.230 62.820 ;
        RECT 257.400 62.330 257.670 62.820 ;
        RECT 254.160 61.840 255.390 62.010 ;
        RECT 252.950 61.120 253.960 61.290 ;
        RECT 254.130 61.275 254.880 61.465 ;
        RECT 252.610 60.780 253.735 60.950 ;
        RECT 254.130 60.610 254.300 61.275 ;
        RECT 255.050 61.030 255.390 61.840 ;
        RECT 255.560 61.530 256.310 62.050 ;
        RECT 256.480 61.360 257.230 61.880 ;
        RECT 257.460 61.580 257.725 62.160 ;
        RECT 257.895 61.890 258.170 62.600 ;
        RECT 258.370 62.335 259.155 62.600 ;
        RECT 257.895 61.660 258.730 61.890 ;
        RECT 252.270 60.440 254.300 60.610 ;
        RECT 254.470 60.270 254.640 61.030 ;
        RECT 254.875 60.620 255.390 61.030 ;
        RECT 255.560 60.270 257.230 61.360 ;
        RECT 257.400 60.270 257.715 61.330 ;
        RECT 257.895 61.000 258.170 61.660 ;
        RECT 258.900 61.480 259.155 62.335 ;
        RECT 259.325 62.140 259.535 62.600 ;
        RECT 259.725 62.325 260.055 62.820 ;
        RECT 260.230 62.190 260.475 62.650 ;
        RECT 259.325 61.660 259.735 62.140 ;
        RECT 260.305 61.980 260.475 62.190 ;
        RECT 260.645 62.160 260.910 62.820 ;
        RECT 261.080 62.100 261.420 62.610 ;
        RECT 259.905 61.480 260.135 61.910 ;
        RECT 258.365 61.310 260.135 61.480 ;
        RECT 260.305 61.460 260.910 61.980 ;
        RECT 258.365 60.945 258.600 61.310 ;
        RECT 258.770 60.950 259.100 61.140 ;
        RECT 259.325 61.015 259.515 61.310 ;
        RECT 260.305 61.120 260.475 61.460 ;
        RECT 258.770 60.775 258.960 60.950 ;
        RECT 258.345 60.270 258.960 60.775 ;
        RECT 259.130 60.440 259.605 60.780 ;
        RECT 259.775 60.270 259.990 61.115 ;
        RECT 260.220 61.110 260.475 61.120 ;
        RECT 260.190 60.440 260.475 61.110 ;
        RECT 260.645 60.270 260.910 61.280 ;
        RECT 261.080 60.700 261.340 62.100 ;
        RECT 261.590 62.020 261.860 62.820 ;
        RECT 261.515 61.580 261.845 61.830 ;
        RECT 262.040 61.580 262.320 62.550 ;
        RECT 262.500 61.580 262.800 62.550 ;
        RECT 262.980 61.580 263.330 62.545 ;
        RECT 263.550 62.320 264.045 62.650 ;
        RECT 261.530 61.410 261.845 61.580 ;
        RECT 263.550 61.410 263.720 62.320 ;
        RECT 261.530 61.240 263.720 61.410 ;
        RECT 261.080 60.440 261.420 60.700 ;
        RECT 261.590 60.270 261.920 61.070 ;
        RECT 262.385 60.440 262.635 61.240 ;
        RECT 262.820 60.270 263.150 60.990 ;
        RECT 263.370 60.440 263.620 61.240 ;
        RECT 263.890 60.830 264.130 62.140 ;
        RECT 265.220 62.095 265.510 62.820 ;
        RECT 265.680 62.275 271.025 62.820 ;
        RECT 271.200 62.275 276.545 62.820 ;
        RECT 267.265 61.445 267.605 62.275 ;
        RECT 263.790 60.270 264.125 60.650 ;
        RECT 265.220 60.270 265.510 61.435 ;
        RECT 269.085 60.705 269.435 61.955 ;
        RECT 272.785 61.445 273.125 62.275 ;
        RECT 277.640 62.190 277.980 62.650 ;
        RECT 278.150 62.360 278.320 62.820 ;
        RECT 278.950 62.385 279.310 62.650 ;
        RECT 278.955 62.380 279.310 62.385 ;
        RECT 278.960 62.370 279.310 62.380 ;
        RECT 278.965 62.365 279.310 62.370 ;
        RECT 278.970 62.355 279.310 62.365 ;
        RECT 279.550 62.360 279.720 62.820 ;
        RECT 278.975 62.350 279.310 62.355 ;
        RECT 278.985 62.340 279.310 62.350 ;
        RECT 278.995 62.330 279.310 62.340 ;
        RECT 278.490 62.190 278.820 62.270 ;
        RECT 277.640 62.000 278.820 62.190 ;
        RECT 279.010 62.190 279.310 62.330 ;
        RECT 279.010 62.000 279.720 62.190 ;
        RECT 274.605 60.705 274.955 61.955 ;
        RECT 277.640 61.630 277.970 61.830 ;
        RECT 278.280 61.810 278.610 61.830 ;
        RECT 278.160 61.630 278.610 61.810 ;
        RECT 277.640 61.290 277.870 61.630 ;
        RECT 265.680 60.270 271.025 60.705 ;
        RECT 271.200 60.270 276.545 60.705 ;
        RECT 277.650 60.270 277.980 60.990 ;
        RECT 278.160 60.515 278.375 61.630 ;
        RECT 278.780 61.600 279.250 61.830 ;
        RECT 279.435 61.430 279.720 62.000 ;
        RECT 279.890 61.875 280.230 62.650 ;
        RECT 280.405 62.270 280.660 62.560 ;
        RECT 280.830 62.440 281.160 62.820 ;
        RECT 280.405 62.100 281.155 62.270 ;
        RECT 278.570 61.215 279.720 61.430 ;
        RECT 278.570 60.440 278.900 61.215 ;
        RECT 279.070 60.270 279.780 61.045 ;
        RECT 279.950 60.440 280.230 61.875 ;
        RECT 280.405 61.280 280.755 61.930 ;
        RECT 280.925 61.110 281.155 62.100 ;
        RECT 280.405 60.940 281.155 61.110 ;
        RECT 280.405 60.440 280.660 60.940 ;
        RECT 280.830 60.270 281.160 60.770 ;
        RECT 281.330 60.440 281.500 62.560 ;
        RECT 281.860 62.460 282.190 62.820 ;
        RECT 282.360 62.430 282.855 62.600 ;
        RECT 283.060 62.430 283.915 62.600 ;
        RECT 281.730 61.240 282.190 62.290 ;
        RECT 281.670 60.455 281.995 61.240 ;
        RECT 282.360 61.070 282.530 62.430 ;
        RECT 282.700 61.520 283.050 62.140 ;
        RECT 283.220 61.920 283.575 62.140 ;
        RECT 283.220 61.330 283.390 61.920 ;
        RECT 283.745 61.720 283.915 62.430 ;
        RECT 284.790 62.360 285.120 62.820 ;
        RECT 285.330 62.460 285.680 62.630 ;
        RECT 284.120 61.890 284.910 62.140 ;
        RECT 285.330 62.070 285.590 62.460 ;
        RECT 285.900 62.370 286.850 62.650 ;
        RECT 287.020 62.380 287.210 62.820 ;
        RECT 287.380 62.440 288.450 62.610 ;
        RECT 285.080 61.720 285.250 61.900 ;
        RECT 282.360 60.900 282.755 61.070 ;
        RECT 282.925 60.940 283.390 61.330 ;
        RECT 283.560 61.550 285.250 61.720 ;
        RECT 282.585 60.770 282.755 60.900 ;
        RECT 283.560 60.770 283.730 61.550 ;
        RECT 285.420 61.380 285.590 62.070 ;
        RECT 284.090 61.210 285.590 61.380 ;
        RECT 285.780 61.410 285.990 62.200 ;
        RECT 286.160 61.580 286.510 62.200 ;
        RECT 286.680 61.590 286.850 62.370 ;
        RECT 287.380 62.210 287.550 62.440 ;
        RECT 287.020 62.040 287.550 62.210 ;
        RECT 287.020 61.760 287.240 62.040 ;
        RECT 287.720 61.870 287.960 62.270 ;
        RECT 286.680 61.420 287.085 61.590 ;
        RECT 287.420 61.500 287.960 61.870 ;
        RECT 288.130 62.085 288.450 62.440 ;
        RECT 288.695 62.360 289.000 62.820 ;
        RECT 289.170 62.110 289.425 62.640 ;
        RECT 288.130 61.910 288.455 62.085 ;
        RECT 288.130 61.610 289.045 61.910 ;
        RECT 288.305 61.580 289.045 61.610 ;
        RECT 285.780 61.250 286.455 61.410 ;
        RECT 286.915 61.330 287.085 61.420 ;
        RECT 285.780 61.240 286.745 61.250 ;
        RECT 285.420 61.070 285.590 61.210 ;
        RECT 282.165 60.270 282.415 60.730 ;
        RECT 282.585 60.440 282.835 60.770 ;
        RECT 283.050 60.440 283.730 60.770 ;
        RECT 283.900 60.870 284.975 61.040 ;
        RECT 285.420 60.900 285.980 61.070 ;
        RECT 286.285 60.950 286.745 61.240 ;
        RECT 286.915 61.160 288.135 61.330 ;
        RECT 283.900 60.530 284.070 60.870 ;
        RECT 284.305 60.270 284.635 60.700 ;
        RECT 284.805 60.530 284.975 60.870 ;
        RECT 285.270 60.270 285.640 60.730 ;
        RECT 285.810 60.440 285.980 60.900 ;
        RECT 286.915 60.780 287.085 61.160 ;
        RECT 288.305 60.990 288.475 61.580 ;
        RECT 289.215 61.460 289.425 62.110 ;
        RECT 289.600 62.070 290.810 62.820 ;
        RECT 290.980 62.095 291.270 62.820 ;
        RECT 289.600 61.530 290.120 62.070 ;
        RECT 291.440 62.050 294.030 62.820 ;
        RECT 286.215 60.440 287.085 60.780 ;
        RECT 287.675 60.820 288.475 60.990 ;
        RECT 287.255 60.270 287.505 60.730 ;
        RECT 287.675 60.530 287.845 60.820 ;
        RECT 288.025 60.270 288.355 60.650 ;
        RECT 288.695 60.270 289.000 61.410 ;
        RECT 289.170 60.580 289.425 61.460 ;
        RECT 290.290 61.360 290.810 61.900 ;
        RECT 291.440 61.530 292.650 62.050 ;
        RECT 294.935 62.010 295.180 62.615 ;
        RECT 295.400 62.285 295.910 62.820 ;
        RECT 289.600 60.270 290.810 61.360 ;
        RECT 290.980 60.270 291.270 61.435 ;
        RECT 292.820 61.360 294.030 61.880 ;
        RECT 291.440 60.270 294.030 61.360 ;
        RECT 294.660 61.840 295.890 62.010 ;
        RECT 294.660 61.030 295.000 61.840 ;
        RECT 295.170 61.275 295.920 61.465 ;
        RECT 294.660 60.620 295.175 61.030 ;
        RECT 295.410 60.270 295.580 61.030 ;
        RECT 295.750 60.610 295.920 61.275 ;
        RECT 296.090 61.290 296.280 62.650 ;
        RECT 296.450 62.480 296.725 62.650 ;
        RECT 296.450 62.310 296.730 62.480 ;
        RECT 296.450 61.490 296.725 62.310 ;
        RECT 296.915 62.285 297.445 62.650 ;
        RECT 297.870 62.420 298.200 62.820 ;
        RECT 297.270 62.250 297.445 62.285 ;
        RECT 296.930 61.290 297.100 62.090 ;
        RECT 296.090 61.120 297.100 61.290 ;
        RECT 297.270 62.080 298.200 62.250 ;
        RECT 298.370 62.080 298.625 62.650 ;
        RECT 297.270 60.950 297.440 62.080 ;
        RECT 298.030 61.910 298.200 62.080 ;
        RECT 296.315 60.780 297.440 60.950 ;
        RECT 297.610 61.580 297.805 61.910 ;
        RECT 298.030 61.580 298.285 61.910 ;
        RECT 297.610 60.610 297.780 61.580 ;
        RECT 298.455 61.410 298.625 62.080 ;
        RECT 295.750 60.440 297.780 60.610 ;
        RECT 297.950 60.270 298.120 61.410 ;
        RECT 298.290 60.440 298.625 61.410 ;
        RECT 298.805 62.080 299.060 62.650 ;
        RECT 299.230 62.420 299.560 62.820 ;
        RECT 299.985 62.285 300.515 62.650 ;
        RECT 299.985 62.250 300.160 62.285 ;
        RECT 299.230 62.080 300.160 62.250 ;
        RECT 300.705 62.140 300.980 62.650 ;
        RECT 298.805 61.410 298.975 62.080 ;
        RECT 299.230 61.910 299.400 62.080 ;
        RECT 299.145 61.580 299.400 61.910 ;
        RECT 299.625 61.580 299.820 61.910 ;
        RECT 298.805 60.440 299.140 61.410 ;
        RECT 299.310 60.270 299.480 61.410 ;
        RECT 299.650 60.610 299.820 61.580 ;
        RECT 299.990 60.950 300.160 62.080 ;
        RECT 300.330 61.290 300.500 62.090 ;
        RECT 300.700 61.970 300.980 62.140 ;
        RECT 300.705 61.490 300.980 61.970 ;
        RECT 301.150 61.290 301.340 62.650 ;
        RECT 301.520 62.285 302.030 62.820 ;
        RECT 302.250 62.010 302.495 62.615 ;
        RECT 302.945 62.080 303.200 62.650 ;
        RECT 303.370 62.420 303.700 62.820 ;
        RECT 304.125 62.285 304.655 62.650 ;
        RECT 304.125 62.250 304.300 62.285 ;
        RECT 303.370 62.080 304.300 62.250 ;
        RECT 301.540 61.840 302.770 62.010 ;
        RECT 300.330 61.120 301.340 61.290 ;
        RECT 301.510 61.275 302.260 61.465 ;
        RECT 299.990 60.780 301.115 60.950 ;
        RECT 301.510 60.610 301.680 61.275 ;
        RECT 302.430 61.030 302.770 61.840 ;
        RECT 299.650 60.440 301.680 60.610 ;
        RECT 301.850 60.270 302.020 61.030 ;
        RECT 302.255 60.620 302.770 61.030 ;
        RECT 302.945 61.410 303.115 62.080 ;
        RECT 303.370 61.910 303.540 62.080 ;
        RECT 303.285 61.580 303.540 61.910 ;
        RECT 303.765 61.580 303.960 61.910 ;
        RECT 302.945 60.440 303.280 61.410 ;
        RECT 303.450 60.270 303.620 61.410 ;
        RECT 303.790 60.610 303.960 61.580 ;
        RECT 304.130 60.950 304.300 62.080 ;
        RECT 304.470 61.290 304.640 62.090 ;
        RECT 304.845 61.800 305.120 62.650 ;
        RECT 304.840 61.630 305.120 61.800 ;
        RECT 304.845 61.490 305.120 61.630 ;
        RECT 305.290 61.290 305.480 62.650 ;
        RECT 305.660 62.285 306.170 62.820 ;
        RECT 306.390 62.010 306.635 62.615 ;
        RECT 307.080 62.050 309.670 62.820 ;
        RECT 309.840 62.070 311.050 62.820 ;
        RECT 305.680 61.840 306.910 62.010 ;
        RECT 304.470 61.120 305.480 61.290 ;
        RECT 305.650 61.275 306.400 61.465 ;
        RECT 304.130 60.780 305.255 60.950 ;
        RECT 305.650 60.610 305.820 61.275 ;
        RECT 306.570 61.030 306.910 61.840 ;
        RECT 307.080 61.530 308.290 62.050 ;
        RECT 308.460 61.360 309.670 61.880 ;
        RECT 303.790 60.440 305.820 60.610 ;
        RECT 305.990 60.270 306.160 61.030 ;
        RECT 306.395 60.620 306.910 61.030 ;
        RECT 307.080 60.270 309.670 61.360 ;
        RECT 309.840 61.360 310.360 61.900 ;
        RECT 310.530 61.530 311.050 62.070 ;
        RECT 309.840 60.270 311.050 61.360 ;
        RECT 162.095 60.100 311.135 60.270 ;
        RECT 162.180 59.010 163.390 60.100 ;
        RECT 163.560 59.665 168.905 60.100 ;
        RECT 162.180 58.300 162.700 58.840 ;
        RECT 162.870 58.470 163.390 59.010 ;
        RECT 162.180 57.550 163.390 58.300 ;
        RECT 165.145 58.095 165.485 58.925 ;
        RECT 166.965 58.415 167.315 59.665 ;
        RECT 169.080 59.010 170.750 60.100 ;
        RECT 169.080 58.320 169.830 58.840 ;
        RECT 170.000 58.490 170.750 59.010 ;
        RECT 170.925 58.960 171.260 59.930 ;
        RECT 171.430 58.960 171.600 60.100 ;
        RECT 171.770 59.760 173.800 59.930 ;
        RECT 163.560 57.550 168.905 58.095 ;
        RECT 169.080 57.550 170.750 58.320 ;
        RECT 170.925 58.290 171.095 58.960 ;
        RECT 171.770 58.790 171.940 59.760 ;
        RECT 171.265 58.460 171.520 58.790 ;
        RECT 171.745 58.460 171.940 58.790 ;
        RECT 172.110 59.420 173.235 59.590 ;
        RECT 171.350 58.290 171.520 58.460 ;
        RECT 172.110 58.290 172.280 59.420 ;
        RECT 170.925 57.720 171.180 58.290 ;
        RECT 171.350 58.120 172.280 58.290 ;
        RECT 172.450 59.080 173.460 59.250 ;
        RECT 172.450 58.280 172.620 59.080 ;
        RECT 172.825 58.740 173.100 58.880 ;
        RECT 172.820 58.570 173.100 58.740 ;
        RECT 172.105 58.085 172.280 58.120 ;
        RECT 171.350 57.550 171.680 57.950 ;
        RECT 172.105 57.720 172.635 58.085 ;
        RECT 172.825 57.720 173.100 58.570 ;
        RECT 173.270 57.720 173.460 59.080 ;
        RECT 173.630 59.095 173.800 59.760 ;
        RECT 173.970 59.340 174.140 60.100 ;
        RECT 174.375 59.340 174.890 59.750 ;
        RECT 173.630 58.905 174.380 59.095 ;
        RECT 174.550 58.530 174.890 59.340 ;
        RECT 175.060 58.935 175.350 60.100 ;
        RECT 175.525 58.950 175.785 60.100 ;
        RECT 175.960 59.025 176.215 59.930 ;
        RECT 176.385 59.340 176.715 60.100 ;
        RECT 176.930 59.170 177.100 59.930 ;
        RECT 173.660 58.360 174.890 58.530 ;
        RECT 173.640 57.550 174.150 58.085 ;
        RECT 174.370 57.755 174.615 58.360 ;
        RECT 175.060 57.550 175.350 58.275 ;
        RECT 175.525 57.550 175.785 58.390 ;
        RECT 175.960 58.295 176.130 59.025 ;
        RECT 176.385 59.000 177.100 59.170 ;
        RECT 176.385 58.790 176.555 59.000 ;
        RECT 177.820 58.960 178.110 60.100 ;
        RECT 178.280 59.380 178.730 59.930 ;
        RECT 178.920 59.380 179.250 60.100 ;
        RECT 176.300 58.460 176.555 58.790 ;
        RECT 175.960 57.720 176.215 58.295 ;
        RECT 176.385 58.270 176.555 58.460 ;
        RECT 176.835 58.450 177.190 58.820 ;
        RECT 176.385 58.100 177.100 58.270 ;
        RECT 176.385 57.550 176.715 57.930 ;
        RECT 176.930 57.720 177.100 58.100 ;
        RECT 177.820 57.550 178.110 58.350 ;
        RECT 178.280 58.010 178.530 59.380 ;
        RECT 179.460 59.210 179.760 59.760 ;
        RECT 179.930 59.430 180.210 60.100 ;
        RECT 178.820 59.040 179.760 59.210 ;
        RECT 178.820 58.790 178.990 59.040 ;
        RECT 180.095 58.790 180.410 59.230 ;
        RECT 180.580 59.010 181.790 60.100 ;
        RECT 178.700 58.460 178.990 58.790 ;
        RECT 179.160 58.540 179.490 58.790 ;
        RECT 179.720 58.540 180.410 58.790 ;
        RECT 178.820 58.370 178.990 58.460 ;
        RECT 178.820 58.180 180.210 58.370 ;
        RECT 178.280 57.720 178.830 58.010 ;
        RECT 179.000 57.550 179.250 58.010 ;
        RECT 179.880 57.820 180.210 58.180 ;
        RECT 180.580 58.300 181.100 58.840 ;
        RECT 181.270 58.470 181.790 59.010 ;
        RECT 181.960 59.675 182.495 59.890 ;
        RECT 183.420 59.675 183.760 60.100 ;
        RECT 184.265 59.675 184.595 60.100 ;
        RECT 185.105 59.675 185.465 60.100 ;
        RECT 180.580 57.550 181.790 58.300 ;
        RECT 181.960 58.290 182.165 59.675 ;
        RECT 185.670 59.505 185.930 59.685 ;
        RECT 182.395 59.335 185.930 59.505 ;
        RECT 186.100 59.400 186.460 60.100 ;
        RECT 186.990 59.570 187.320 59.910 ;
        RECT 187.850 59.740 188.520 60.100 ;
        RECT 188.690 59.570 188.880 59.930 ;
        RECT 189.050 59.720 189.400 60.100 ;
        RECT 186.990 59.550 188.880 59.570 ;
        RECT 186.990 59.340 189.410 59.550 ;
        RECT 182.395 58.790 182.625 59.335 ;
        RECT 185.250 59.275 185.930 59.335 ;
        RECT 188.690 59.295 189.410 59.340 ;
        RECT 182.335 58.460 182.625 58.790 ;
        RECT 182.815 58.460 183.125 59.165 ;
        RECT 183.295 58.880 183.615 59.165 ;
        RECT 183.795 58.880 185.080 59.165 ;
        RECT 183.295 58.460 183.480 58.880 ;
        RECT 183.650 58.540 184.740 58.710 ;
        RECT 183.650 58.355 183.820 58.540 ;
        RECT 184.910 58.370 185.080 58.880 ;
        RECT 183.615 58.290 183.820 58.355 ;
        RECT 181.960 58.185 183.820 58.290 ;
        RECT 183.990 58.200 185.080 58.370 ;
        RECT 185.250 58.370 185.420 59.275 ;
        RECT 185.590 58.540 185.930 59.105 ;
        RECT 186.135 58.960 188.055 59.170 ;
        RECT 186.135 58.460 186.505 58.960 ;
        RECT 186.845 58.460 187.395 58.790 ;
        RECT 187.750 58.455 188.055 58.960 ;
        RECT 188.380 58.540 189.050 59.080 ;
        RECT 189.220 58.800 189.410 59.295 ;
        RECT 189.580 59.165 189.760 59.930 ;
        RECT 189.930 59.335 190.260 60.100 ;
        RECT 190.430 59.165 190.620 59.930 ;
        RECT 190.790 59.335 191.120 60.100 ;
        RECT 191.620 59.760 192.800 59.930 ;
        RECT 189.580 58.995 191.445 59.165 ;
        RECT 189.220 58.460 191.045 58.800 ;
        RECT 185.250 58.200 185.930 58.370 ;
        RECT 189.220 58.335 189.420 58.460 ;
        RECT 181.960 58.120 183.765 58.185 ;
        RECT 181.960 58.070 182.355 58.120 ;
        RECT 182.100 57.770 182.355 58.070 ;
        RECT 182.525 57.550 182.915 57.950 ;
        RECT 183.085 57.770 183.255 58.120 ;
        RECT 183.990 58.050 184.160 58.200 ;
        RECT 183.425 57.550 183.755 57.950 ;
        RECT 183.925 57.720 184.160 58.050 ;
        RECT 184.345 57.550 184.515 58.030 ;
        RECT 184.685 57.750 185.015 58.200 ;
        RECT 185.225 57.550 185.395 58.030 ;
        RECT 185.670 57.755 185.930 58.200 ;
        RECT 186.130 58.080 188.260 58.250 ;
        RECT 188.440 58.120 189.420 58.335 ;
        RECT 191.215 58.270 191.445 58.995 ;
        RECT 191.620 58.960 191.960 59.760 ;
        RECT 192.130 58.790 192.365 59.515 ;
        RECT 192.535 59.130 192.800 59.760 ;
        RECT 192.970 59.300 193.670 60.100 ;
        RECT 192.535 58.960 193.625 59.130 ;
        RECT 191.620 58.540 191.960 58.790 ;
        RECT 192.130 58.540 192.590 58.790 ;
        RECT 192.760 58.540 193.235 58.790 ;
        RECT 193.405 58.710 193.625 58.960 ;
        RECT 193.880 59.090 194.130 59.930 ;
        RECT 194.300 59.260 194.550 60.100 ;
        RECT 194.720 59.090 194.970 59.930 ;
        RECT 195.140 59.260 195.390 60.100 ;
        RECT 195.960 59.430 196.240 60.100 ;
        RECT 196.410 59.210 196.710 59.760 ;
        RECT 196.910 59.380 197.240 60.100 ;
        RECT 197.430 59.380 197.890 59.930 ;
        RECT 193.880 58.920 195.590 59.090 ;
        RECT 193.980 58.910 194.150 58.920 ;
        RECT 193.405 58.540 195.130 58.710 ;
        RECT 193.405 58.370 193.625 58.540 ;
        RECT 195.300 58.370 195.590 58.920 ;
        RECT 195.775 58.790 196.040 59.150 ;
        RECT 196.410 59.040 197.350 59.210 ;
        RECT 197.180 58.790 197.350 59.040 ;
        RECT 195.775 58.540 196.450 58.790 ;
        RECT 196.670 58.540 197.010 58.790 ;
        RECT 197.180 58.460 197.470 58.790 ;
        RECT 197.180 58.370 197.350 58.460 ;
        RECT 189.820 58.100 191.445 58.270 ;
        RECT 191.620 58.190 193.625 58.370 ;
        RECT 193.840 58.200 195.590 58.370 ;
        RECT 189.820 58.080 190.940 58.100 ;
        RECT 187.930 57.950 188.260 58.080 ;
        RECT 186.560 57.550 186.890 57.910 ;
        RECT 187.420 57.550 187.760 57.910 ;
        RECT 187.930 57.720 189.200 57.950 ;
        RECT 189.390 57.550 189.720 57.930 ;
        RECT 190.250 57.550 190.580 57.910 ;
        RECT 191.110 57.550 191.440 57.930 ;
        RECT 191.620 57.720 191.960 58.190 ;
        RECT 192.130 57.550 192.300 58.020 ;
        RECT 192.470 57.720 192.800 58.190 ;
        RECT 192.970 57.550 193.670 58.020 ;
        RECT 193.840 57.730 194.170 58.200 ;
        RECT 194.340 57.550 194.510 58.020 ;
        RECT 194.680 57.730 195.010 58.200 ;
        RECT 195.960 58.180 197.350 58.370 ;
        RECT 195.180 57.550 195.350 58.020 ;
        RECT 195.960 57.820 196.290 58.180 ;
        RECT 197.640 58.010 197.890 59.380 ;
        RECT 198.060 59.010 200.650 60.100 ;
        RECT 196.910 57.550 197.160 58.010 ;
        RECT 197.330 57.720 197.890 58.010 ;
        RECT 198.060 58.320 199.270 58.840 ;
        RECT 199.440 58.490 200.650 59.010 ;
        RECT 200.820 58.935 201.110 60.100 ;
        RECT 201.280 59.300 201.720 59.930 ;
        RECT 198.060 57.550 200.650 58.320 ;
        RECT 201.280 58.290 201.590 59.300 ;
        RECT 201.895 59.250 202.210 60.100 ;
        RECT 202.380 59.760 203.810 59.930 ;
        RECT 202.380 59.080 202.550 59.760 ;
        RECT 201.760 58.910 202.550 59.080 ;
        RECT 201.760 58.460 201.930 58.910 ;
        RECT 202.720 58.790 202.920 59.590 ;
        RECT 202.100 58.460 202.490 58.740 ;
        RECT 202.675 58.460 202.920 58.790 ;
        RECT 203.120 58.460 203.370 59.590 ;
        RECT 203.560 59.130 203.810 59.760 ;
        RECT 203.990 59.300 204.320 60.100 ;
        RECT 204.500 59.665 209.845 60.100 ;
        RECT 203.560 58.960 204.330 59.130 ;
        RECT 203.585 58.460 203.990 58.790 ;
        RECT 204.160 58.290 204.330 58.960 ;
        RECT 200.820 57.550 201.110 58.275 ;
        RECT 201.280 57.730 201.720 58.290 ;
        RECT 201.890 57.550 202.340 58.290 ;
        RECT 202.510 58.120 203.670 58.290 ;
        RECT 202.510 57.720 202.680 58.120 ;
        RECT 202.850 57.550 203.270 57.950 ;
        RECT 203.440 57.720 203.670 58.120 ;
        RECT 203.840 57.720 204.330 58.290 ;
        RECT 206.085 58.095 206.425 58.925 ;
        RECT 207.905 58.415 208.255 59.665 ;
        RECT 210.020 59.010 212.610 60.100 ;
        RECT 210.020 58.320 211.230 58.840 ;
        RECT 211.400 58.490 212.610 59.010 ;
        RECT 213.240 58.960 213.625 59.920 ;
        RECT 213.840 59.300 214.130 60.100 ;
        RECT 214.300 59.760 215.665 59.930 ;
        RECT 214.300 59.130 214.470 59.760 ;
        RECT 213.795 58.960 214.470 59.130 ;
        RECT 204.500 57.550 209.845 58.095 ;
        RECT 210.020 57.550 212.610 58.320 ;
        RECT 213.240 58.290 213.415 58.960 ;
        RECT 213.795 58.790 213.965 58.960 ;
        RECT 214.640 58.790 214.965 59.590 ;
        RECT 215.335 59.550 215.665 59.760 ;
        RECT 215.335 59.300 216.290 59.550 ;
        RECT 213.600 58.540 213.965 58.790 ;
        RECT 214.160 58.540 214.410 58.790 ;
        RECT 213.600 58.460 213.790 58.540 ;
        RECT 214.160 58.460 214.330 58.540 ;
        RECT 214.620 58.460 214.965 58.790 ;
        RECT 215.135 58.460 215.410 59.125 ;
        RECT 215.595 58.460 215.950 59.125 ;
        RECT 216.120 58.290 216.290 59.300 ;
        RECT 216.460 58.960 216.750 60.100 ;
        RECT 216.920 59.300 217.360 59.930 ;
        RECT 216.475 58.460 216.750 58.790 ;
        RECT 213.240 57.720 213.750 58.290 ;
        RECT 214.295 58.120 215.695 58.290 ;
        RECT 213.920 57.550 214.090 58.110 ;
        RECT 214.295 57.720 214.625 58.120 ;
        RECT 214.800 57.550 215.130 57.950 ;
        RECT 215.365 57.930 215.695 58.120 ;
        RECT 215.865 58.100 216.290 58.290 ;
        RECT 216.920 58.290 217.230 59.300 ;
        RECT 217.535 59.250 217.850 60.100 ;
        RECT 218.020 59.760 219.450 59.930 ;
        RECT 218.020 59.080 218.190 59.760 ;
        RECT 217.400 58.910 218.190 59.080 ;
        RECT 217.400 58.460 217.570 58.910 ;
        RECT 218.360 58.790 218.560 59.590 ;
        RECT 217.740 58.460 218.130 58.740 ;
        RECT 218.315 58.460 218.560 58.790 ;
        RECT 218.760 58.460 219.010 59.590 ;
        RECT 219.200 59.130 219.450 59.760 ;
        RECT 219.630 59.300 219.960 60.100 ;
        RECT 219.200 58.960 219.970 59.130 ;
        RECT 219.225 58.460 219.630 58.790 ;
        RECT 219.800 58.290 219.970 58.960 ;
        RECT 216.460 57.930 216.750 58.200 ;
        RECT 215.365 57.720 216.750 57.930 ;
        RECT 216.920 57.730 217.360 58.290 ;
        RECT 217.530 57.550 217.980 58.290 ;
        RECT 218.150 58.120 219.310 58.290 ;
        RECT 218.150 57.720 218.320 58.120 ;
        RECT 218.490 57.550 218.910 57.950 ;
        RECT 219.080 57.720 219.310 58.120 ;
        RECT 219.480 57.720 219.970 58.290 ;
        RECT 220.145 58.960 220.480 59.930 ;
        RECT 220.650 58.960 220.820 60.100 ;
        RECT 220.990 59.760 223.020 59.930 ;
        RECT 220.145 58.290 220.315 58.960 ;
        RECT 220.990 58.790 221.160 59.760 ;
        RECT 220.485 58.460 220.740 58.790 ;
        RECT 220.965 58.460 221.160 58.790 ;
        RECT 221.330 59.420 222.455 59.590 ;
        RECT 220.570 58.290 220.740 58.460 ;
        RECT 221.330 58.290 221.500 59.420 ;
        RECT 220.145 57.720 220.400 58.290 ;
        RECT 220.570 58.120 221.500 58.290 ;
        RECT 221.670 59.080 222.680 59.250 ;
        RECT 221.670 58.280 221.840 59.080 ;
        RECT 222.045 58.740 222.320 58.880 ;
        RECT 222.040 58.570 222.320 58.740 ;
        RECT 221.325 58.085 221.500 58.120 ;
        RECT 220.570 57.550 220.900 57.950 ;
        RECT 221.325 57.720 221.855 58.085 ;
        RECT 222.045 57.720 222.320 58.570 ;
        RECT 222.490 57.720 222.680 59.080 ;
        RECT 222.850 59.095 223.020 59.760 ;
        RECT 223.190 59.340 223.360 60.100 ;
        RECT 223.595 59.340 224.110 59.750 ;
        RECT 222.850 58.905 223.600 59.095 ;
        RECT 223.770 58.530 224.110 59.340 ;
        RECT 222.880 58.360 224.110 58.530 ;
        RECT 224.315 59.310 224.850 59.930 ;
        RECT 222.860 57.550 223.370 58.085 ;
        RECT 223.590 57.755 223.835 58.360 ;
        RECT 224.315 58.290 224.630 59.310 ;
        RECT 225.020 59.300 225.350 60.100 ;
        RECT 225.835 59.130 226.225 59.305 ;
        RECT 224.800 58.960 226.225 59.130 ;
        RECT 224.800 58.460 224.970 58.960 ;
        RECT 224.315 57.720 224.930 58.290 ;
        RECT 225.220 58.230 225.485 58.790 ;
        RECT 225.655 58.060 225.825 58.960 ;
        RECT 226.580 58.935 226.870 60.100 ;
        RECT 227.155 59.470 227.440 59.930 ;
        RECT 227.610 59.640 227.880 60.100 ;
        RECT 227.155 59.250 228.110 59.470 ;
        RECT 225.995 58.230 226.350 58.790 ;
        RECT 227.040 58.520 227.730 59.080 ;
        RECT 227.900 58.350 228.110 59.250 ;
        RECT 225.100 57.550 225.315 58.060 ;
        RECT 225.545 57.730 225.825 58.060 ;
        RECT 226.005 57.550 226.245 58.060 ;
        RECT 226.580 57.550 226.870 58.275 ;
        RECT 227.155 58.180 228.110 58.350 ;
        RECT 228.280 59.080 228.680 59.930 ;
        RECT 228.870 59.470 229.150 59.930 ;
        RECT 229.670 59.640 229.995 60.100 ;
        RECT 228.870 59.250 229.995 59.470 ;
        RECT 228.280 58.520 229.375 59.080 ;
        RECT 229.545 58.790 229.995 59.250 ;
        RECT 230.165 58.960 230.550 59.930 ;
        RECT 230.720 59.010 232.390 60.100 ;
        RECT 232.565 59.430 232.820 59.930 ;
        RECT 232.990 59.600 233.320 60.100 ;
        RECT 232.565 59.260 233.315 59.430 ;
        RECT 227.155 57.720 227.440 58.180 ;
        RECT 227.610 57.550 227.880 58.010 ;
        RECT 228.280 57.720 228.680 58.520 ;
        RECT 229.545 58.460 230.100 58.790 ;
        RECT 229.545 58.350 229.995 58.460 ;
        RECT 228.870 58.180 229.995 58.350 ;
        RECT 230.270 58.290 230.550 58.960 ;
        RECT 228.870 57.720 229.150 58.180 ;
        RECT 229.670 57.550 229.995 58.010 ;
        RECT 230.165 57.720 230.550 58.290 ;
        RECT 230.720 58.320 231.470 58.840 ;
        RECT 231.640 58.490 232.390 59.010 ;
        RECT 232.565 58.440 232.915 59.090 ;
        RECT 230.720 57.550 232.390 58.320 ;
        RECT 233.085 58.270 233.315 59.260 ;
        RECT 232.565 58.100 233.315 58.270 ;
        RECT 232.565 57.810 232.820 58.100 ;
        RECT 232.990 57.550 233.320 57.930 ;
        RECT 233.490 57.810 233.660 59.930 ;
        RECT 233.830 59.130 234.155 59.915 ;
        RECT 234.325 59.640 234.575 60.100 ;
        RECT 234.745 59.600 234.995 59.930 ;
        RECT 235.210 59.600 235.890 59.930 ;
        RECT 234.745 59.470 234.915 59.600 ;
        RECT 234.520 59.300 234.915 59.470 ;
        RECT 233.890 58.080 234.350 59.130 ;
        RECT 234.520 57.940 234.690 59.300 ;
        RECT 235.085 59.040 235.550 59.430 ;
        RECT 234.860 58.230 235.210 58.850 ;
        RECT 235.380 58.450 235.550 59.040 ;
        RECT 235.720 58.820 235.890 59.600 ;
        RECT 236.060 59.500 236.230 59.840 ;
        RECT 236.465 59.670 236.795 60.100 ;
        RECT 236.965 59.500 237.135 59.840 ;
        RECT 237.430 59.640 237.800 60.100 ;
        RECT 236.060 59.330 237.135 59.500 ;
        RECT 237.970 59.470 238.140 59.930 ;
        RECT 238.375 59.590 239.245 59.930 ;
        RECT 239.415 59.640 239.665 60.100 ;
        RECT 237.580 59.300 238.140 59.470 ;
        RECT 237.580 59.160 237.750 59.300 ;
        RECT 236.250 58.990 237.750 59.160 ;
        RECT 238.445 59.130 238.905 59.420 ;
        RECT 235.720 58.650 237.410 58.820 ;
        RECT 235.380 58.230 235.735 58.450 ;
        RECT 235.905 57.940 236.075 58.650 ;
        RECT 236.280 58.230 237.070 58.480 ;
        RECT 237.240 58.470 237.410 58.650 ;
        RECT 237.580 58.300 237.750 58.990 ;
        RECT 234.020 57.550 234.350 57.910 ;
        RECT 234.520 57.770 235.015 57.940 ;
        RECT 235.220 57.770 236.075 57.940 ;
        RECT 236.950 57.550 237.280 58.010 ;
        RECT 237.490 57.910 237.750 58.300 ;
        RECT 237.940 59.120 238.905 59.130 ;
        RECT 239.075 59.210 239.245 59.590 ;
        RECT 239.835 59.550 240.005 59.840 ;
        RECT 240.185 59.720 240.515 60.100 ;
        RECT 239.835 59.380 240.635 59.550 ;
        RECT 237.940 58.960 238.615 59.120 ;
        RECT 239.075 59.040 240.295 59.210 ;
        RECT 237.940 58.170 238.150 58.960 ;
        RECT 239.075 58.950 239.245 59.040 ;
        RECT 238.320 58.170 238.670 58.790 ;
        RECT 238.840 58.780 239.245 58.950 ;
        RECT 238.840 58.000 239.010 58.780 ;
        RECT 239.180 58.330 239.400 58.610 ;
        RECT 239.580 58.500 240.120 58.870 ;
        RECT 240.465 58.790 240.635 59.380 ;
        RECT 240.855 58.960 241.160 60.100 ;
        RECT 241.330 58.910 241.585 59.790 ;
        RECT 241.845 59.480 242.020 59.930 ;
        RECT 242.190 59.660 242.520 60.100 ;
        RECT 242.825 59.510 242.995 59.930 ;
        RECT 243.230 59.690 243.900 60.100 ;
        RECT 244.115 59.510 244.285 59.930 ;
        RECT 244.485 59.690 244.815 60.100 ;
        RECT 241.845 59.310 242.475 59.480 ;
        RECT 240.465 58.760 241.205 58.790 ;
        RECT 239.180 58.160 239.710 58.330 ;
        RECT 237.490 57.740 237.840 57.910 ;
        RECT 238.060 57.720 239.010 58.000 ;
        RECT 239.180 57.550 239.370 57.990 ;
        RECT 239.540 57.930 239.710 58.160 ;
        RECT 239.880 58.100 240.120 58.500 ;
        RECT 240.290 58.460 241.205 58.760 ;
        RECT 240.290 58.285 240.615 58.460 ;
        RECT 240.290 57.930 240.610 58.285 ;
        RECT 241.375 58.260 241.585 58.910 ;
        RECT 241.760 58.460 242.125 59.140 ;
        RECT 242.305 58.790 242.475 59.310 ;
        RECT 242.825 59.340 244.840 59.510 ;
        RECT 242.305 58.460 242.655 58.790 ;
        RECT 242.305 58.290 242.475 58.460 ;
        RECT 239.540 57.760 240.610 57.930 ;
        RECT 240.855 57.550 241.160 58.010 ;
        RECT 241.330 57.730 241.585 58.260 ;
        RECT 241.845 58.120 242.475 58.290 ;
        RECT 241.845 57.720 242.020 58.120 ;
        RECT 242.825 58.050 242.995 59.340 ;
        RECT 242.190 57.550 242.520 57.930 ;
        RECT 242.765 57.720 242.995 58.050 ;
        RECT 243.195 57.885 243.475 59.160 ;
        RECT 243.700 58.060 243.970 59.160 ;
        RECT 244.160 58.130 244.500 59.160 ;
        RECT 244.670 58.790 244.840 59.340 ;
        RECT 245.010 58.960 245.270 59.930 ;
        RECT 245.440 59.010 246.650 60.100 ;
        RECT 244.670 58.460 244.930 58.790 ;
        RECT 245.100 58.270 245.270 58.960 ;
        RECT 243.660 57.890 243.970 58.060 ;
        RECT 243.700 57.885 243.970 57.890 ;
        RECT 244.430 57.550 244.760 57.930 ;
        RECT 244.930 57.805 245.270 58.270 ;
        RECT 245.440 58.300 245.960 58.840 ;
        RECT 246.130 58.470 246.650 59.010 ;
        RECT 246.900 59.170 247.080 59.930 ;
        RECT 247.260 59.340 247.590 60.100 ;
        RECT 246.900 59.000 247.575 59.170 ;
        RECT 247.760 59.025 248.030 59.930 ;
        RECT 247.405 58.855 247.575 59.000 ;
        RECT 246.840 58.450 247.180 58.820 ;
        RECT 247.405 58.525 247.680 58.855 ;
        RECT 244.930 57.760 245.265 57.805 ;
        RECT 245.440 57.550 246.650 58.300 ;
        RECT 247.405 58.270 247.575 58.525 ;
        RECT 246.910 58.100 247.575 58.270 ;
        RECT 247.850 58.225 248.030 59.025 ;
        RECT 248.200 59.340 248.715 59.750 ;
        RECT 248.950 59.340 249.120 60.100 ;
        RECT 249.290 59.760 251.320 59.930 ;
        RECT 248.200 58.530 248.540 59.340 ;
        RECT 249.290 59.095 249.460 59.760 ;
        RECT 249.855 59.420 250.980 59.590 ;
        RECT 248.710 58.905 249.460 59.095 ;
        RECT 249.630 59.080 250.640 59.250 ;
        RECT 248.200 58.360 249.430 58.530 ;
        RECT 246.910 57.720 247.080 58.100 ;
        RECT 247.260 57.550 247.590 57.930 ;
        RECT 247.770 57.720 248.030 58.225 ;
        RECT 248.475 57.755 248.720 58.360 ;
        RECT 248.940 57.550 249.450 58.085 ;
        RECT 249.630 57.720 249.820 59.080 ;
        RECT 249.990 58.740 250.265 58.880 ;
        RECT 249.990 58.570 250.270 58.740 ;
        RECT 249.990 57.720 250.265 58.570 ;
        RECT 250.470 58.280 250.640 59.080 ;
        RECT 250.810 58.290 250.980 59.420 ;
        RECT 251.150 58.790 251.320 59.760 ;
        RECT 251.490 58.960 251.660 60.100 ;
        RECT 251.830 58.960 252.165 59.930 ;
        RECT 251.150 58.460 251.345 58.790 ;
        RECT 251.570 58.460 251.825 58.790 ;
        RECT 251.570 58.290 251.740 58.460 ;
        RECT 251.995 58.290 252.165 58.960 ;
        RECT 252.340 58.935 252.630 60.100 ;
        RECT 252.805 59.430 253.060 59.930 ;
        RECT 253.230 59.600 253.560 60.100 ;
        RECT 252.805 59.260 253.555 59.430 ;
        RECT 252.805 58.440 253.155 59.090 ;
        RECT 250.810 58.120 251.740 58.290 ;
        RECT 250.810 58.085 250.985 58.120 ;
        RECT 250.455 57.720 250.985 58.085 ;
        RECT 251.410 57.550 251.740 57.950 ;
        RECT 251.910 57.720 252.165 58.290 ;
        RECT 252.340 57.550 252.630 58.275 ;
        RECT 253.325 58.270 253.555 59.260 ;
        RECT 252.805 58.100 253.555 58.270 ;
        RECT 252.805 57.810 253.060 58.100 ;
        RECT 253.230 57.550 253.560 57.930 ;
        RECT 253.730 57.810 253.900 59.930 ;
        RECT 254.070 59.130 254.395 59.915 ;
        RECT 254.565 59.640 254.815 60.100 ;
        RECT 254.985 59.600 255.235 59.930 ;
        RECT 255.450 59.600 256.130 59.930 ;
        RECT 254.985 59.470 255.155 59.600 ;
        RECT 254.760 59.300 255.155 59.470 ;
        RECT 254.130 58.080 254.590 59.130 ;
        RECT 254.760 57.940 254.930 59.300 ;
        RECT 255.325 59.040 255.790 59.430 ;
        RECT 255.100 58.230 255.450 58.850 ;
        RECT 255.620 58.450 255.790 59.040 ;
        RECT 255.960 58.820 256.130 59.600 ;
        RECT 256.300 59.500 256.470 59.840 ;
        RECT 256.705 59.670 257.035 60.100 ;
        RECT 257.205 59.500 257.375 59.840 ;
        RECT 257.670 59.640 258.040 60.100 ;
        RECT 256.300 59.330 257.375 59.500 ;
        RECT 258.210 59.470 258.380 59.930 ;
        RECT 258.615 59.590 259.485 59.930 ;
        RECT 259.655 59.640 259.905 60.100 ;
        RECT 257.820 59.300 258.380 59.470 ;
        RECT 257.820 59.160 257.990 59.300 ;
        RECT 256.490 58.990 257.990 59.160 ;
        RECT 258.685 59.130 259.145 59.420 ;
        RECT 255.960 58.650 257.650 58.820 ;
        RECT 255.620 58.230 255.975 58.450 ;
        RECT 256.145 57.940 256.315 58.650 ;
        RECT 256.520 58.230 257.310 58.480 ;
        RECT 257.480 58.470 257.650 58.650 ;
        RECT 257.820 58.300 257.990 58.990 ;
        RECT 254.260 57.550 254.590 57.910 ;
        RECT 254.760 57.770 255.255 57.940 ;
        RECT 255.460 57.770 256.315 57.940 ;
        RECT 257.190 57.550 257.520 58.010 ;
        RECT 257.730 57.910 257.990 58.300 ;
        RECT 258.180 59.120 259.145 59.130 ;
        RECT 259.315 59.210 259.485 59.590 ;
        RECT 260.075 59.550 260.245 59.840 ;
        RECT 260.425 59.720 260.755 60.100 ;
        RECT 260.075 59.380 260.875 59.550 ;
        RECT 258.180 58.960 258.855 59.120 ;
        RECT 259.315 59.040 260.535 59.210 ;
        RECT 258.180 58.170 258.390 58.960 ;
        RECT 259.315 58.950 259.485 59.040 ;
        RECT 258.560 58.170 258.910 58.790 ;
        RECT 259.080 58.780 259.485 58.950 ;
        RECT 259.080 58.000 259.250 58.780 ;
        RECT 259.420 58.330 259.640 58.610 ;
        RECT 259.820 58.500 260.360 58.870 ;
        RECT 260.705 58.790 260.875 59.380 ;
        RECT 261.095 58.960 261.400 60.100 ;
        RECT 261.570 58.910 261.825 59.790 ;
        RECT 262.000 59.665 267.345 60.100 ;
        RECT 269.120 59.740 269.450 60.100 ;
        RECT 269.975 59.740 270.310 60.100 ;
        RECT 270.880 59.740 271.210 60.100 ;
        RECT 271.775 59.740 272.225 60.100 ;
        RECT 260.705 58.760 261.445 58.790 ;
        RECT 259.420 58.160 259.950 58.330 ;
        RECT 257.730 57.740 258.080 57.910 ;
        RECT 258.300 57.720 259.250 58.000 ;
        RECT 259.420 57.550 259.610 57.990 ;
        RECT 259.780 57.930 259.950 58.160 ;
        RECT 260.120 58.100 260.360 58.500 ;
        RECT 260.530 58.460 261.445 58.760 ;
        RECT 260.530 58.285 260.855 58.460 ;
        RECT 260.530 57.930 260.850 58.285 ;
        RECT 261.615 58.260 261.825 58.910 ;
        RECT 259.780 57.760 260.850 57.930 ;
        RECT 261.095 57.550 261.400 58.010 ;
        RECT 261.570 57.730 261.825 58.260 ;
        RECT 263.585 58.095 263.925 58.925 ;
        RECT 265.405 58.415 265.755 59.665 ;
        RECT 268.510 59.340 272.275 59.570 ;
        RECT 262.000 57.550 267.345 58.095 ;
        RECT 268.510 57.890 268.790 59.340 ;
        RECT 268.960 58.080 269.240 59.170 ;
        RECT 269.420 59.000 270.730 59.170 ;
        RECT 269.420 58.310 269.685 59.000 ;
        RECT 270.900 58.990 271.675 59.160 ;
        RECT 270.900 58.820 271.070 58.990 ;
        RECT 269.855 58.485 271.070 58.820 ;
        RECT 269.420 58.080 270.670 58.310 ;
        RECT 270.840 58.270 271.070 58.485 ;
        RECT 271.240 58.460 271.430 58.805 ;
        RECT 270.840 58.080 271.535 58.270 ;
        RECT 271.720 58.190 271.935 58.805 ;
        RECT 272.105 58.790 272.275 59.340 ;
        RECT 272.445 58.960 272.805 59.630 ;
        RECT 273.040 59.010 276.550 60.100 ;
        RECT 276.720 59.010 277.930 60.100 ;
        RECT 272.105 58.460 272.415 58.790 ;
        RECT 272.585 58.270 272.805 58.960 ;
        RECT 269.120 57.550 269.450 57.910 ;
        RECT 269.620 57.720 269.810 58.080 ;
        RECT 270.480 57.980 270.670 58.080 ;
        RECT 271.355 58.010 271.535 58.080 ;
        RECT 272.320 58.010 272.805 58.270 ;
        RECT 269.980 57.550 270.310 57.910 ;
        RECT 270.845 57.550 271.175 57.910 ;
        RECT 271.355 57.820 272.805 58.010 ;
        RECT 272.320 57.720 272.805 57.820 ;
        RECT 273.040 58.320 274.690 58.840 ;
        RECT 274.860 58.490 276.550 59.010 ;
        RECT 273.040 57.550 276.550 58.320 ;
        RECT 276.720 58.300 277.240 58.840 ;
        RECT 277.410 58.470 277.930 59.010 ;
        RECT 278.100 58.935 278.390 60.100 ;
        RECT 278.560 59.340 279.075 59.750 ;
        RECT 279.310 59.340 279.480 60.100 ;
        RECT 279.650 59.760 281.680 59.930 ;
        RECT 278.560 58.530 278.900 59.340 ;
        RECT 279.650 59.095 279.820 59.760 ;
        RECT 280.215 59.420 281.340 59.590 ;
        RECT 279.070 58.905 279.820 59.095 ;
        RECT 279.990 59.080 281.000 59.250 ;
        RECT 278.560 58.360 279.790 58.530 ;
        RECT 276.720 57.550 277.930 58.300 ;
        RECT 278.100 57.550 278.390 58.275 ;
        RECT 278.835 57.755 279.080 58.360 ;
        RECT 279.300 57.550 279.810 58.085 ;
        RECT 279.990 57.720 280.180 59.080 ;
        RECT 280.350 58.400 280.625 58.880 ;
        RECT 280.350 58.230 280.630 58.400 ;
        RECT 280.830 58.280 281.000 59.080 ;
        RECT 281.170 58.290 281.340 59.420 ;
        RECT 281.510 58.790 281.680 59.760 ;
        RECT 281.850 58.960 282.020 60.100 ;
        RECT 282.190 58.960 282.525 59.930 ;
        RECT 283.625 59.430 283.880 59.930 ;
        RECT 284.050 59.600 284.380 60.100 ;
        RECT 283.625 59.260 284.375 59.430 ;
        RECT 281.510 58.460 281.705 58.790 ;
        RECT 281.930 58.460 282.185 58.790 ;
        RECT 281.930 58.290 282.100 58.460 ;
        RECT 282.355 58.290 282.525 58.960 ;
        RECT 283.625 58.440 283.975 59.090 ;
        RECT 280.350 57.720 280.625 58.230 ;
        RECT 281.170 58.120 282.100 58.290 ;
        RECT 281.170 58.085 281.345 58.120 ;
        RECT 280.815 57.720 281.345 58.085 ;
        RECT 281.770 57.550 282.100 57.950 ;
        RECT 282.270 57.720 282.525 58.290 ;
        RECT 284.145 58.270 284.375 59.260 ;
        RECT 283.625 58.100 284.375 58.270 ;
        RECT 283.625 57.810 283.880 58.100 ;
        RECT 284.050 57.550 284.380 57.930 ;
        RECT 284.550 57.810 284.720 59.930 ;
        RECT 284.890 59.130 285.215 59.915 ;
        RECT 285.385 59.640 285.635 60.100 ;
        RECT 285.805 59.600 286.055 59.930 ;
        RECT 286.270 59.600 286.950 59.930 ;
        RECT 285.805 59.470 285.975 59.600 ;
        RECT 285.580 59.300 285.975 59.470 ;
        RECT 284.950 58.080 285.410 59.130 ;
        RECT 285.580 57.940 285.750 59.300 ;
        RECT 286.145 59.040 286.610 59.430 ;
        RECT 285.920 58.230 286.270 58.850 ;
        RECT 286.440 58.450 286.610 59.040 ;
        RECT 286.780 58.820 286.950 59.600 ;
        RECT 287.120 59.500 287.290 59.840 ;
        RECT 287.525 59.670 287.855 60.100 ;
        RECT 288.025 59.500 288.195 59.840 ;
        RECT 288.490 59.640 288.860 60.100 ;
        RECT 287.120 59.330 288.195 59.500 ;
        RECT 289.030 59.470 289.200 59.930 ;
        RECT 289.435 59.590 290.305 59.930 ;
        RECT 290.475 59.640 290.725 60.100 ;
        RECT 288.640 59.300 289.200 59.470 ;
        RECT 288.640 59.160 288.810 59.300 ;
        RECT 287.310 58.990 288.810 59.160 ;
        RECT 289.505 59.130 289.965 59.420 ;
        RECT 286.780 58.650 288.470 58.820 ;
        RECT 286.440 58.230 286.795 58.450 ;
        RECT 286.965 57.940 287.135 58.650 ;
        RECT 287.340 58.230 288.130 58.480 ;
        RECT 288.300 58.470 288.470 58.650 ;
        RECT 288.640 58.300 288.810 58.990 ;
        RECT 285.080 57.550 285.410 57.910 ;
        RECT 285.580 57.770 286.075 57.940 ;
        RECT 286.280 57.770 287.135 57.940 ;
        RECT 288.010 57.550 288.340 58.010 ;
        RECT 288.550 57.910 288.810 58.300 ;
        RECT 289.000 59.120 289.965 59.130 ;
        RECT 290.135 59.210 290.305 59.590 ;
        RECT 290.895 59.550 291.065 59.840 ;
        RECT 291.245 59.720 291.575 60.100 ;
        RECT 290.895 59.380 291.695 59.550 ;
        RECT 289.000 58.960 289.675 59.120 ;
        RECT 290.135 59.040 291.355 59.210 ;
        RECT 289.000 58.170 289.210 58.960 ;
        RECT 290.135 58.950 290.305 59.040 ;
        RECT 289.380 58.170 289.730 58.790 ;
        RECT 289.900 58.780 290.305 58.950 ;
        RECT 289.900 58.000 290.070 58.780 ;
        RECT 290.240 58.330 290.460 58.610 ;
        RECT 290.640 58.500 291.180 58.870 ;
        RECT 291.525 58.790 291.695 59.380 ;
        RECT 291.915 58.960 292.220 60.100 ;
        RECT 292.390 58.910 292.640 59.790 ;
        RECT 292.810 58.960 293.060 60.100 ;
        RECT 293.280 59.010 294.490 60.100 ;
        RECT 291.525 58.760 292.265 58.790 ;
        RECT 290.240 58.160 290.770 58.330 ;
        RECT 288.550 57.740 288.900 57.910 ;
        RECT 289.120 57.720 290.070 58.000 ;
        RECT 290.240 57.550 290.430 57.990 ;
        RECT 290.600 57.930 290.770 58.160 ;
        RECT 290.940 58.100 291.180 58.500 ;
        RECT 291.350 58.460 292.265 58.760 ;
        RECT 291.350 58.285 291.675 58.460 ;
        RECT 291.350 57.930 291.670 58.285 ;
        RECT 292.435 58.260 292.640 58.910 ;
        RECT 290.600 57.760 291.670 57.930 ;
        RECT 291.915 57.550 292.220 58.010 ;
        RECT 292.390 57.730 292.640 58.260 ;
        RECT 292.810 57.550 293.060 58.305 ;
        RECT 293.280 58.300 293.800 58.840 ;
        RECT 293.970 58.470 294.490 59.010 ;
        RECT 294.665 58.910 294.920 59.790 ;
        RECT 295.090 58.960 295.395 60.100 ;
        RECT 295.735 59.720 296.065 60.100 ;
        RECT 296.245 59.550 296.415 59.840 ;
        RECT 296.585 59.640 296.835 60.100 ;
        RECT 295.615 59.380 296.415 59.550 ;
        RECT 297.005 59.590 297.875 59.930 ;
        RECT 293.280 57.550 294.490 58.300 ;
        RECT 294.665 58.260 294.875 58.910 ;
        RECT 295.615 58.790 295.785 59.380 ;
        RECT 297.005 59.210 297.175 59.590 ;
        RECT 298.110 59.470 298.280 59.930 ;
        RECT 298.450 59.640 298.820 60.100 ;
        RECT 299.115 59.500 299.285 59.840 ;
        RECT 299.455 59.670 299.785 60.100 ;
        RECT 300.020 59.500 300.190 59.840 ;
        RECT 295.955 59.040 297.175 59.210 ;
        RECT 297.345 59.130 297.805 59.420 ;
        RECT 298.110 59.300 298.670 59.470 ;
        RECT 299.115 59.330 300.190 59.500 ;
        RECT 300.360 59.600 301.040 59.930 ;
        RECT 301.255 59.600 301.505 59.930 ;
        RECT 301.675 59.640 301.925 60.100 ;
        RECT 298.500 59.160 298.670 59.300 ;
        RECT 297.345 59.120 298.310 59.130 ;
        RECT 297.005 58.950 297.175 59.040 ;
        RECT 297.635 58.960 298.310 59.120 ;
        RECT 295.045 58.760 295.785 58.790 ;
        RECT 295.045 58.460 295.960 58.760 ;
        RECT 295.635 58.285 295.960 58.460 ;
        RECT 294.665 57.730 294.920 58.260 ;
        RECT 295.090 57.550 295.395 58.010 ;
        RECT 295.640 57.930 295.960 58.285 ;
        RECT 296.130 58.500 296.670 58.870 ;
        RECT 297.005 58.780 297.410 58.950 ;
        RECT 296.130 58.100 296.370 58.500 ;
        RECT 296.850 58.330 297.070 58.610 ;
        RECT 296.540 58.160 297.070 58.330 ;
        RECT 296.540 57.930 296.710 58.160 ;
        RECT 297.240 58.000 297.410 58.780 ;
        RECT 297.580 58.170 297.930 58.790 ;
        RECT 298.100 58.170 298.310 58.960 ;
        RECT 298.500 58.990 300.000 59.160 ;
        RECT 298.500 58.300 298.670 58.990 ;
        RECT 300.360 58.820 300.530 59.600 ;
        RECT 301.335 59.470 301.505 59.600 ;
        RECT 298.840 58.650 300.530 58.820 ;
        RECT 300.700 59.040 301.165 59.430 ;
        RECT 301.335 59.300 301.730 59.470 ;
        RECT 298.840 58.470 299.010 58.650 ;
        RECT 295.640 57.760 296.710 57.930 ;
        RECT 296.880 57.550 297.070 57.990 ;
        RECT 297.240 57.720 298.190 58.000 ;
        RECT 298.500 57.910 298.760 58.300 ;
        RECT 299.180 58.230 299.970 58.480 ;
        RECT 298.410 57.740 298.760 57.910 ;
        RECT 298.970 57.550 299.300 58.010 ;
        RECT 300.175 57.940 300.345 58.650 ;
        RECT 300.700 58.450 300.870 59.040 ;
        RECT 300.515 58.230 300.870 58.450 ;
        RECT 301.040 58.230 301.390 58.850 ;
        RECT 301.560 57.940 301.730 59.300 ;
        RECT 302.095 59.130 302.420 59.915 ;
        RECT 301.900 58.080 302.360 59.130 ;
        RECT 300.175 57.770 301.030 57.940 ;
        RECT 301.235 57.770 301.730 57.940 ;
        RECT 301.900 57.550 302.230 57.910 ;
        RECT 302.590 57.810 302.760 59.930 ;
        RECT 302.930 59.600 303.260 60.100 ;
        RECT 303.430 59.430 303.685 59.930 ;
        RECT 302.935 59.260 303.685 59.430 ;
        RECT 302.935 58.270 303.165 59.260 ;
        RECT 303.335 58.440 303.685 59.090 ;
        RECT 303.860 58.935 304.150 60.100 ;
        RECT 304.320 59.665 309.665 60.100 ;
        RECT 302.935 58.100 303.685 58.270 ;
        RECT 302.930 57.550 303.260 57.930 ;
        RECT 303.430 57.810 303.685 58.100 ;
        RECT 303.860 57.550 304.150 58.275 ;
        RECT 305.905 58.095 306.245 58.925 ;
        RECT 307.725 58.415 308.075 59.665 ;
        RECT 309.840 59.010 311.050 60.100 ;
        RECT 309.840 58.470 310.360 59.010 ;
        RECT 310.530 58.300 311.050 58.840 ;
        RECT 304.320 57.550 309.665 58.095 ;
        RECT 309.840 57.550 311.050 58.300 ;
        RECT 162.095 57.380 311.135 57.550 ;
        RECT 162.180 56.630 163.390 57.380 ;
        RECT 162.180 56.090 162.700 56.630 ;
        RECT 163.560 56.610 166.150 57.380 ;
        RECT 166.325 56.830 166.580 57.120 ;
        RECT 166.750 57.000 167.080 57.380 ;
        RECT 166.325 56.660 167.075 56.830 ;
        RECT 162.870 55.920 163.390 56.460 ;
        RECT 163.560 56.090 164.770 56.610 ;
        RECT 164.940 55.920 166.150 56.440 ;
        RECT 162.180 54.830 163.390 55.920 ;
        RECT 163.560 54.830 166.150 55.920 ;
        RECT 166.325 55.840 166.675 56.490 ;
        RECT 166.845 55.670 167.075 56.660 ;
        RECT 166.325 55.500 167.075 55.670 ;
        RECT 166.325 55.000 166.580 55.500 ;
        RECT 166.750 54.830 167.080 55.330 ;
        RECT 167.250 55.000 167.420 57.120 ;
        RECT 167.780 57.020 168.110 57.380 ;
        RECT 168.280 56.990 168.775 57.160 ;
        RECT 168.980 56.990 169.835 57.160 ;
        RECT 167.650 55.800 168.110 56.850 ;
        RECT 167.590 55.015 167.915 55.800 ;
        RECT 168.280 55.630 168.450 56.990 ;
        RECT 168.620 56.080 168.970 56.700 ;
        RECT 169.140 56.480 169.495 56.700 ;
        RECT 169.140 55.890 169.310 56.480 ;
        RECT 169.665 56.280 169.835 56.990 ;
        RECT 170.710 56.920 171.040 57.380 ;
        RECT 171.250 57.020 171.600 57.190 ;
        RECT 170.040 56.450 170.830 56.700 ;
        RECT 171.250 56.630 171.510 57.020 ;
        RECT 171.820 56.930 172.770 57.210 ;
        RECT 172.940 56.940 173.130 57.380 ;
        RECT 173.300 57.000 174.370 57.170 ;
        RECT 171.000 56.280 171.170 56.460 ;
        RECT 168.280 55.460 168.675 55.630 ;
        RECT 168.845 55.500 169.310 55.890 ;
        RECT 169.480 56.110 171.170 56.280 ;
        RECT 168.505 55.330 168.675 55.460 ;
        RECT 169.480 55.330 169.650 56.110 ;
        RECT 171.340 55.940 171.510 56.630 ;
        RECT 170.010 55.770 171.510 55.940 ;
        RECT 171.700 55.970 171.910 56.760 ;
        RECT 172.080 56.140 172.430 56.760 ;
        RECT 172.600 56.150 172.770 56.930 ;
        RECT 173.300 56.770 173.470 57.000 ;
        RECT 172.940 56.600 173.470 56.770 ;
        RECT 172.940 56.320 173.160 56.600 ;
        RECT 173.640 56.430 173.880 56.830 ;
        RECT 172.600 55.980 173.005 56.150 ;
        RECT 173.340 56.060 173.880 56.430 ;
        RECT 174.050 56.645 174.370 57.000 ;
        RECT 174.615 56.920 174.920 57.380 ;
        RECT 175.090 56.670 175.345 57.200 ;
        RECT 174.050 56.470 174.375 56.645 ;
        RECT 174.050 56.170 174.965 56.470 ;
        RECT 174.225 56.140 174.965 56.170 ;
        RECT 171.700 55.810 172.375 55.970 ;
        RECT 172.835 55.890 173.005 55.980 ;
        RECT 171.700 55.800 172.665 55.810 ;
        RECT 171.340 55.630 171.510 55.770 ;
        RECT 168.085 54.830 168.335 55.290 ;
        RECT 168.505 55.000 168.755 55.330 ;
        RECT 168.970 55.000 169.650 55.330 ;
        RECT 169.820 55.430 170.895 55.600 ;
        RECT 171.340 55.460 171.900 55.630 ;
        RECT 172.205 55.510 172.665 55.800 ;
        RECT 172.835 55.720 174.055 55.890 ;
        RECT 169.820 55.090 169.990 55.430 ;
        RECT 170.225 54.830 170.555 55.260 ;
        RECT 170.725 55.090 170.895 55.430 ;
        RECT 171.190 54.830 171.560 55.290 ;
        RECT 171.730 55.000 171.900 55.460 ;
        RECT 172.835 55.340 173.005 55.720 ;
        RECT 174.225 55.550 174.395 56.140 ;
        RECT 175.135 56.020 175.345 56.670 ;
        RECT 172.135 55.000 173.005 55.340 ;
        RECT 173.595 55.380 174.395 55.550 ;
        RECT 173.175 54.830 173.425 55.290 ;
        RECT 173.595 55.090 173.765 55.380 ;
        RECT 173.945 54.830 174.275 55.210 ;
        RECT 174.615 54.830 174.920 55.970 ;
        RECT 175.090 55.140 175.345 56.020 ;
        RECT 175.525 56.640 175.780 57.210 ;
        RECT 175.950 56.980 176.280 57.380 ;
        RECT 176.705 56.845 177.235 57.210 ;
        RECT 177.425 57.040 177.700 57.210 ;
        RECT 177.420 56.870 177.700 57.040 ;
        RECT 176.705 56.810 176.880 56.845 ;
        RECT 175.950 56.640 176.880 56.810 ;
        RECT 175.525 55.970 175.695 56.640 ;
        RECT 175.950 56.470 176.120 56.640 ;
        RECT 175.865 56.140 176.120 56.470 ;
        RECT 176.345 56.140 176.540 56.470 ;
        RECT 175.525 55.000 175.860 55.970 ;
        RECT 176.030 54.830 176.200 55.970 ;
        RECT 176.370 55.170 176.540 56.140 ;
        RECT 176.710 55.510 176.880 56.640 ;
        RECT 177.050 55.850 177.220 56.650 ;
        RECT 177.425 56.050 177.700 56.870 ;
        RECT 177.870 55.850 178.060 57.210 ;
        RECT 178.240 56.845 178.750 57.380 ;
        RECT 178.970 56.570 179.215 57.175 ;
        RECT 179.660 56.580 179.950 57.380 ;
        RECT 180.120 56.920 180.670 57.210 ;
        RECT 180.840 56.920 181.090 57.380 ;
        RECT 178.260 56.400 179.490 56.570 ;
        RECT 177.050 55.680 178.060 55.850 ;
        RECT 178.230 55.835 178.980 56.025 ;
        RECT 176.710 55.340 177.835 55.510 ;
        RECT 178.230 55.170 178.400 55.835 ;
        RECT 179.150 55.590 179.490 56.400 ;
        RECT 176.370 55.000 178.400 55.170 ;
        RECT 178.570 54.830 178.740 55.590 ;
        RECT 178.975 55.180 179.490 55.590 ;
        RECT 179.660 54.830 179.950 55.970 ;
        RECT 180.120 55.550 180.370 56.920 ;
        RECT 181.720 56.750 182.050 57.110 ;
        RECT 180.660 56.560 182.050 56.750 ;
        RECT 183.345 56.810 183.600 57.080 ;
        RECT 183.770 56.980 184.100 57.380 ;
        RECT 184.270 56.810 184.440 57.080 ;
        RECT 184.610 56.980 184.940 57.380 ;
        RECT 185.225 56.920 185.975 57.210 ;
        RECT 186.485 56.920 186.815 57.380 ;
        RECT 183.345 56.640 184.570 56.810 ;
        RECT 180.660 56.470 180.830 56.560 ;
        RECT 180.540 56.140 180.830 56.470 ;
        RECT 181.000 56.140 181.330 56.390 ;
        RECT 181.560 56.140 182.250 56.390 ;
        RECT 183.345 56.140 183.680 56.470 ;
        RECT 183.850 56.140 184.230 56.470 ;
        RECT 180.660 55.890 180.830 56.140 ;
        RECT 180.660 55.720 181.600 55.890 ;
        RECT 180.120 55.000 180.570 55.550 ;
        RECT 180.760 54.830 181.090 55.550 ;
        RECT 181.300 55.170 181.600 55.720 ;
        RECT 181.935 55.700 182.250 56.140 ;
        RECT 181.770 54.830 182.050 55.500 ;
        RECT 183.345 55.185 183.680 55.970 ;
        RECT 183.850 55.460 184.085 56.140 ;
        RECT 184.400 55.970 184.570 56.640 ;
        RECT 184.255 55.800 184.570 55.970 ;
        RECT 184.740 55.800 185.010 56.810 ;
        RECT 184.255 55.340 184.425 55.800 ;
        RECT 185.225 55.630 185.595 56.920 ;
        RECT 187.035 56.730 187.305 56.940 ;
        RECT 185.970 56.560 187.305 56.730 ;
        RECT 187.940 56.655 188.230 57.380 ;
        RECT 188.405 57.125 188.740 57.170 ;
        RECT 188.400 56.660 188.740 57.125 ;
        RECT 188.910 57.000 189.240 57.380 ;
        RECT 185.970 56.390 186.140 56.560 ;
        RECT 185.765 56.140 186.140 56.390 ;
        RECT 186.310 56.150 186.785 56.390 ;
        RECT 186.955 56.150 187.305 56.390 ;
        RECT 185.970 55.970 186.140 56.140 ;
        RECT 185.970 55.800 187.305 55.970 ;
        RECT 187.025 55.640 187.305 55.800 ;
        RECT 184.255 55.185 184.490 55.340 ;
        RECT 183.345 55.170 184.490 55.185 ;
        RECT 183.345 55.015 184.425 55.170 ;
        RECT 184.690 54.830 185.005 55.630 ;
        RECT 185.225 55.460 186.395 55.630 ;
        RECT 185.680 54.830 185.895 55.290 ;
        RECT 186.065 55.000 186.395 55.460 ;
        RECT 186.565 54.830 186.815 55.630 ;
        RECT 187.940 54.830 188.230 55.995 ;
        RECT 188.400 55.970 188.570 56.660 ;
        RECT 188.740 56.140 189.000 56.470 ;
        RECT 188.400 55.000 188.660 55.970 ;
        RECT 188.830 55.590 189.000 56.140 ;
        RECT 189.170 55.770 189.510 56.800 ;
        RECT 189.700 56.700 189.970 57.045 ;
        RECT 189.700 56.530 190.010 56.700 ;
        RECT 189.700 55.770 189.970 56.530 ;
        RECT 190.195 55.770 190.475 57.045 ;
        RECT 190.675 56.880 190.905 57.210 ;
        RECT 191.150 57.000 191.480 57.380 ;
        RECT 190.675 55.590 190.845 56.880 ;
        RECT 191.650 56.810 191.825 57.210 ;
        RECT 192.165 56.880 192.660 57.210 ;
        RECT 191.195 56.640 191.825 56.810 ;
        RECT 191.195 56.470 191.365 56.640 ;
        RECT 191.015 56.140 191.365 56.470 ;
        RECT 188.830 55.420 190.845 55.590 ;
        RECT 191.195 55.620 191.365 56.140 ;
        RECT 191.545 55.790 191.910 56.470 ;
        RECT 191.195 55.450 191.825 55.620 ;
        RECT 188.855 54.830 189.185 55.240 ;
        RECT 189.385 55.000 189.555 55.420 ;
        RECT 189.770 54.830 190.440 55.240 ;
        RECT 190.675 55.000 190.845 55.420 ;
        RECT 191.150 54.830 191.480 55.270 ;
        RECT 191.650 55.000 191.825 55.450 ;
        RECT 192.080 55.390 192.320 56.700 ;
        RECT 192.490 55.970 192.660 56.880 ;
        RECT 192.880 56.140 193.230 57.105 ;
        RECT 193.410 56.140 193.710 57.110 ;
        RECT 193.890 56.140 194.170 57.110 ;
        RECT 194.350 56.580 194.620 57.380 ;
        RECT 194.790 56.660 195.130 57.170 ;
        RECT 195.305 56.830 195.560 57.120 ;
        RECT 195.730 57.000 196.060 57.380 ;
        RECT 195.305 56.660 196.055 56.830 ;
        RECT 194.365 56.140 194.695 56.390 ;
        RECT 194.365 55.970 194.680 56.140 ;
        RECT 192.490 55.800 194.680 55.970 ;
        RECT 192.085 54.830 192.420 55.210 ;
        RECT 192.590 55.000 192.840 55.800 ;
        RECT 193.060 54.830 193.390 55.550 ;
        RECT 193.575 55.000 193.825 55.800 ;
        RECT 194.290 54.830 194.620 55.630 ;
        RECT 194.870 55.260 195.130 56.660 ;
        RECT 195.305 55.840 195.655 56.490 ;
        RECT 195.825 55.670 196.055 56.660 ;
        RECT 194.790 55.000 195.130 55.260 ;
        RECT 195.305 55.500 196.055 55.670 ;
        RECT 195.305 55.000 195.560 55.500 ;
        RECT 195.730 54.830 196.060 55.330 ;
        RECT 196.230 55.000 196.400 57.120 ;
        RECT 196.760 57.020 197.090 57.380 ;
        RECT 197.260 56.990 197.755 57.160 ;
        RECT 197.960 56.990 198.815 57.160 ;
        RECT 196.630 55.800 197.090 56.850 ;
        RECT 196.570 55.015 196.895 55.800 ;
        RECT 197.260 55.630 197.430 56.990 ;
        RECT 197.600 56.080 197.950 56.700 ;
        RECT 198.120 56.480 198.475 56.700 ;
        RECT 198.120 55.890 198.290 56.480 ;
        RECT 198.645 56.280 198.815 56.990 ;
        RECT 199.690 56.920 200.020 57.380 ;
        RECT 200.230 57.020 200.580 57.190 ;
        RECT 199.020 56.450 199.810 56.700 ;
        RECT 200.230 56.630 200.490 57.020 ;
        RECT 200.800 56.930 201.750 57.210 ;
        RECT 201.920 56.940 202.110 57.380 ;
        RECT 202.280 57.000 203.350 57.170 ;
        RECT 199.980 56.280 200.150 56.460 ;
        RECT 197.260 55.460 197.655 55.630 ;
        RECT 197.825 55.500 198.290 55.890 ;
        RECT 198.460 56.110 200.150 56.280 ;
        RECT 197.485 55.330 197.655 55.460 ;
        RECT 198.460 55.330 198.630 56.110 ;
        RECT 200.320 55.940 200.490 56.630 ;
        RECT 198.990 55.770 200.490 55.940 ;
        RECT 200.680 55.970 200.890 56.760 ;
        RECT 201.060 56.140 201.410 56.760 ;
        RECT 201.580 56.150 201.750 56.930 ;
        RECT 202.280 56.770 202.450 57.000 ;
        RECT 201.920 56.600 202.450 56.770 ;
        RECT 201.920 56.320 202.140 56.600 ;
        RECT 202.620 56.430 202.860 56.830 ;
        RECT 201.580 55.980 201.985 56.150 ;
        RECT 202.320 56.060 202.860 56.430 ;
        RECT 203.030 56.645 203.350 57.000 ;
        RECT 203.595 56.920 203.900 57.380 ;
        RECT 204.070 56.670 204.325 57.200 ;
        RECT 203.030 56.470 203.355 56.645 ;
        RECT 203.030 56.170 203.945 56.470 ;
        RECT 203.205 56.140 203.945 56.170 ;
        RECT 200.680 55.810 201.355 55.970 ;
        RECT 201.815 55.890 201.985 55.980 ;
        RECT 200.680 55.800 201.645 55.810 ;
        RECT 200.320 55.630 200.490 55.770 ;
        RECT 197.065 54.830 197.315 55.290 ;
        RECT 197.485 55.000 197.735 55.330 ;
        RECT 197.950 55.000 198.630 55.330 ;
        RECT 198.800 55.430 199.875 55.600 ;
        RECT 200.320 55.460 200.880 55.630 ;
        RECT 201.185 55.510 201.645 55.800 ;
        RECT 201.815 55.720 203.035 55.890 ;
        RECT 198.800 55.090 198.970 55.430 ;
        RECT 199.205 54.830 199.535 55.260 ;
        RECT 199.705 55.090 199.875 55.430 ;
        RECT 200.170 54.830 200.540 55.290 ;
        RECT 200.710 55.000 200.880 55.460 ;
        RECT 201.815 55.340 201.985 55.720 ;
        RECT 203.205 55.550 203.375 56.140 ;
        RECT 204.115 56.020 204.325 56.670 ;
        RECT 201.115 55.000 201.985 55.340 ;
        RECT 202.575 55.380 203.375 55.550 ;
        RECT 202.155 54.830 202.405 55.290 ;
        RECT 202.575 55.090 202.745 55.380 ;
        RECT 202.925 54.830 203.255 55.210 ;
        RECT 203.595 54.830 203.900 55.970 ;
        RECT 204.070 55.140 204.325 56.020 ;
        RECT 204.535 56.640 205.150 57.210 ;
        RECT 205.320 56.870 205.535 57.380 ;
        RECT 205.765 56.870 206.045 57.200 ;
        RECT 206.225 56.870 206.465 57.380 ;
        RECT 204.535 55.620 204.850 56.640 ;
        RECT 205.020 55.970 205.190 56.470 ;
        RECT 205.440 56.140 205.705 56.700 ;
        RECT 205.875 55.970 206.045 56.870 ;
        RECT 206.215 56.140 206.570 56.700 ;
        RECT 206.800 56.610 210.310 57.380 ;
        RECT 211.565 56.870 211.805 57.380 ;
        RECT 211.985 56.870 212.265 57.200 ;
        RECT 212.495 56.870 212.710 57.380 ;
        RECT 206.800 56.090 208.450 56.610 ;
        RECT 205.020 55.800 206.445 55.970 ;
        RECT 208.620 55.920 210.310 56.440 ;
        RECT 211.460 56.140 211.815 56.700 ;
        RECT 211.985 55.970 212.155 56.870 ;
        RECT 212.325 56.140 212.590 56.700 ;
        RECT 212.880 56.640 213.495 57.210 ;
        RECT 213.700 56.655 213.990 57.380 ;
        RECT 212.840 55.970 213.010 56.470 ;
        RECT 204.535 55.000 205.070 55.620 ;
        RECT 205.240 54.830 205.570 55.630 ;
        RECT 206.055 55.625 206.445 55.800 ;
        RECT 206.800 54.830 210.310 55.920 ;
        RECT 211.585 55.800 213.010 55.970 ;
        RECT 211.585 55.625 211.975 55.800 ;
        RECT 212.460 54.830 212.790 55.630 ;
        RECT 213.180 55.620 213.495 56.640 ;
        RECT 214.160 56.630 215.370 57.380 ;
        RECT 215.540 56.640 215.925 57.210 ;
        RECT 216.095 56.920 216.420 57.380 ;
        RECT 216.940 56.750 217.220 57.210 ;
        RECT 214.160 56.090 214.680 56.630 ;
        RECT 212.960 55.000 213.495 55.620 ;
        RECT 213.700 54.830 213.990 55.995 ;
        RECT 214.850 55.920 215.370 56.460 ;
        RECT 214.160 54.830 215.370 55.920 ;
        RECT 215.540 55.970 215.820 56.640 ;
        RECT 216.095 56.580 217.220 56.750 ;
        RECT 216.095 56.470 216.545 56.580 ;
        RECT 215.990 56.140 216.545 56.470 ;
        RECT 217.410 56.410 217.810 57.210 ;
        RECT 218.210 56.920 218.480 57.380 ;
        RECT 218.650 56.750 218.935 57.210 ;
        RECT 215.540 55.000 215.925 55.970 ;
        RECT 216.095 55.680 216.545 56.140 ;
        RECT 216.715 55.850 217.810 56.410 ;
        RECT 216.095 55.460 217.220 55.680 ;
        RECT 216.095 54.830 216.420 55.290 ;
        RECT 216.940 55.000 217.220 55.460 ;
        RECT 217.410 55.000 217.810 55.850 ;
        RECT 217.980 56.580 218.935 56.750 ;
        RECT 219.225 56.830 219.480 57.120 ;
        RECT 219.650 57.000 219.980 57.380 ;
        RECT 219.225 56.660 219.975 56.830 ;
        RECT 217.980 55.680 218.190 56.580 ;
        RECT 218.360 55.850 219.050 56.410 ;
        RECT 219.225 55.840 219.575 56.490 ;
        RECT 217.980 55.460 218.935 55.680 ;
        RECT 219.745 55.670 219.975 56.660 ;
        RECT 218.210 54.830 218.480 55.290 ;
        RECT 218.650 55.000 218.935 55.460 ;
        RECT 219.225 55.500 219.975 55.670 ;
        RECT 219.225 55.000 219.480 55.500 ;
        RECT 219.650 54.830 219.980 55.330 ;
        RECT 220.150 55.000 220.320 57.120 ;
        RECT 220.680 57.020 221.010 57.380 ;
        RECT 221.180 56.990 221.675 57.160 ;
        RECT 221.880 56.990 222.735 57.160 ;
        RECT 220.550 55.800 221.010 56.850 ;
        RECT 220.490 55.015 220.815 55.800 ;
        RECT 221.180 55.630 221.350 56.990 ;
        RECT 221.520 56.080 221.870 56.700 ;
        RECT 222.040 56.480 222.395 56.700 ;
        RECT 222.040 55.890 222.210 56.480 ;
        RECT 222.565 56.280 222.735 56.990 ;
        RECT 223.610 56.920 223.940 57.380 ;
        RECT 224.150 57.020 224.500 57.190 ;
        RECT 222.940 56.450 223.730 56.700 ;
        RECT 224.150 56.630 224.410 57.020 ;
        RECT 224.720 56.930 225.670 57.210 ;
        RECT 225.840 56.940 226.030 57.380 ;
        RECT 226.200 57.000 227.270 57.170 ;
        RECT 223.900 56.280 224.070 56.460 ;
        RECT 221.180 55.460 221.575 55.630 ;
        RECT 221.745 55.500 222.210 55.890 ;
        RECT 222.380 56.110 224.070 56.280 ;
        RECT 221.405 55.330 221.575 55.460 ;
        RECT 222.380 55.330 222.550 56.110 ;
        RECT 224.240 55.940 224.410 56.630 ;
        RECT 222.910 55.770 224.410 55.940 ;
        RECT 224.600 55.970 224.810 56.760 ;
        RECT 224.980 56.140 225.330 56.760 ;
        RECT 225.500 56.150 225.670 56.930 ;
        RECT 226.200 56.770 226.370 57.000 ;
        RECT 225.840 56.600 226.370 56.770 ;
        RECT 225.840 56.320 226.060 56.600 ;
        RECT 226.540 56.430 226.780 56.830 ;
        RECT 225.500 55.980 225.905 56.150 ;
        RECT 226.240 56.060 226.780 56.430 ;
        RECT 226.950 56.645 227.270 57.000 ;
        RECT 227.515 56.920 227.820 57.380 ;
        RECT 227.990 56.670 228.245 57.200 ;
        RECT 226.950 56.470 227.275 56.645 ;
        RECT 226.950 56.170 227.865 56.470 ;
        RECT 227.125 56.140 227.865 56.170 ;
        RECT 224.600 55.810 225.275 55.970 ;
        RECT 225.735 55.890 225.905 55.980 ;
        RECT 224.600 55.800 225.565 55.810 ;
        RECT 224.240 55.630 224.410 55.770 ;
        RECT 220.985 54.830 221.235 55.290 ;
        RECT 221.405 55.000 221.655 55.330 ;
        RECT 221.870 55.000 222.550 55.330 ;
        RECT 222.720 55.430 223.795 55.600 ;
        RECT 224.240 55.460 224.800 55.630 ;
        RECT 225.105 55.510 225.565 55.800 ;
        RECT 225.735 55.720 226.955 55.890 ;
        RECT 222.720 55.090 222.890 55.430 ;
        RECT 223.125 54.830 223.455 55.260 ;
        RECT 223.625 55.090 223.795 55.430 ;
        RECT 224.090 54.830 224.460 55.290 ;
        RECT 224.630 55.000 224.800 55.460 ;
        RECT 225.735 55.340 225.905 55.720 ;
        RECT 227.125 55.550 227.295 56.140 ;
        RECT 228.035 56.020 228.245 56.670 ;
        RECT 228.425 56.830 228.680 57.120 ;
        RECT 228.850 57.000 229.180 57.380 ;
        RECT 228.425 56.660 229.175 56.830 ;
        RECT 225.035 55.000 225.905 55.340 ;
        RECT 226.495 55.380 227.295 55.550 ;
        RECT 226.075 54.830 226.325 55.290 ;
        RECT 226.495 55.090 226.665 55.380 ;
        RECT 226.845 54.830 227.175 55.210 ;
        RECT 227.515 54.830 227.820 55.970 ;
        RECT 227.990 55.140 228.245 56.020 ;
        RECT 228.425 55.840 228.775 56.490 ;
        RECT 228.945 55.670 229.175 56.660 ;
        RECT 228.425 55.500 229.175 55.670 ;
        RECT 228.425 55.000 228.680 55.500 ;
        RECT 228.850 54.830 229.180 55.330 ;
        RECT 229.350 55.000 229.520 57.120 ;
        RECT 229.880 57.020 230.210 57.380 ;
        RECT 230.380 56.990 230.875 57.160 ;
        RECT 231.080 56.990 231.935 57.160 ;
        RECT 229.750 55.800 230.210 56.850 ;
        RECT 229.690 55.015 230.015 55.800 ;
        RECT 230.380 55.630 230.550 56.990 ;
        RECT 230.720 56.080 231.070 56.700 ;
        RECT 231.240 56.480 231.595 56.700 ;
        RECT 231.240 55.890 231.410 56.480 ;
        RECT 231.765 56.280 231.935 56.990 ;
        RECT 232.810 56.920 233.140 57.380 ;
        RECT 233.350 57.020 233.700 57.190 ;
        RECT 232.140 56.450 232.930 56.700 ;
        RECT 233.350 56.630 233.610 57.020 ;
        RECT 233.920 56.930 234.870 57.210 ;
        RECT 235.040 56.940 235.230 57.380 ;
        RECT 235.400 57.000 236.470 57.170 ;
        RECT 233.100 56.280 233.270 56.460 ;
        RECT 230.380 55.460 230.775 55.630 ;
        RECT 230.945 55.500 231.410 55.890 ;
        RECT 231.580 56.110 233.270 56.280 ;
        RECT 230.605 55.330 230.775 55.460 ;
        RECT 231.580 55.330 231.750 56.110 ;
        RECT 233.440 55.940 233.610 56.630 ;
        RECT 232.110 55.770 233.610 55.940 ;
        RECT 233.800 55.970 234.010 56.760 ;
        RECT 234.180 56.140 234.530 56.760 ;
        RECT 234.700 56.150 234.870 56.930 ;
        RECT 235.400 56.770 235.570 57.000 ;
        RECT 235.040 56.600 235.570 56.770 ;
        RECT 235.040 56.320 235.260 56.600 ;
        RECT 235.740 56.430 235.980 56.830 ;
        RECT 234.700 55.980 235.105 56.150 ;
        RECT 235.440 56.060 235.980 56.430 ;
        RECT 236.150 56.645 236.470 57.000 ;
        RECT 236.715 56.920 237.020 57.380 ;
        RECT 237.190 56.670 237.445 57.200 ;
        RECT 236.150 56.470 236.475 56.645 ;
        RECT 236.150 56.170 237.065 56.470 ;
        RECT 236.325 56.140 237.065 56.170 ;
        RECT 233.800 55.810 234.475 55.970 ;
        RECT 234.935 55.890 235.105 55.980 ;
        RECT 233.800 55.800 234.765 55.810 ;
        RECT 233.440 55.630 233.610 55.770 ;
        RECT 230.185 54.830 230.435 55.290 ;
        RECT 230.605 55.000 230.855 55.330 ;
        RECT 231.070 55.000 231.750 55.330 ;
        RECT 231.920 55.430 232.995 55.600 ;
        RECT 233.440 55.460 234.000 55.630 ;
        RECT 234.305 55.510 234.765 55.800 ;
        RECT 234.935 55.720 236.155 55.890 ;
        RECT 231.920 55.090 232.090 55.430 ;
        RECT 232.325 54.830 232.655 55.260 ;
        RECT 232.825 55.090 232.995 55.430 ;
        RECT 233.290 54.830 233.660 55.290 ;
        RECT 233.830 55.000 234.000 55.460 ;
        RECT 234.935 55.340 235.105 55.720 ;
        RECT 236.325 55.550 236.495 56.140 ;
        RECT 237.235 56.020 237.445 56.670 ;
        RECT 237.620 56.610 239.290 57.380 ;
        RECT 239.460 56.655 239.750 57.380 ;
        RECT 239.955 56.640 240.570 57.210 ;
        RECT 240.740 56.870 240.955 57.380 ;
        RECT 241.185 56.870 241.465 57.200 ;
        RECT 241.645 56.870 241.885 57.380 ;
        RECT 237.620 56.090 238.370 56.610 ;
        RECT 234.235 55.000 235.105 55.340 ;
        RECT 235.695 55.380 236.495 55.550 ;
        RECT 235.275 54.830 235.525 55.290 ;
        RECT 235.695 55.090 235.865 55.380 ;
        RECT 236.045 54.830 236.375 55.210 ;
        RECT 236.715 54.830 237.020 55.970 ;
        RECT 237.190 55.140 237.445 56.020 ;
        RECT 238.540 55.920 239.290 56.440 ;
        RECT 237.620 54.830 239.290 55.920 ;
        RECT 239.460 54.830 239.750 55.995 ;
        RECT 239.955 55.620 240.270 56.640 ;
        RECT 240.440 55.970 240.610 56.470 ;
        RECT 240.860 56.140 241.125 56.700 ;
        RECT 241.295 55.970 241.465 56.870 ;
        RECT 241.635 56.140 241.990 56.700 ;
        RECT 242.255 56.640 242.870 57.210 ;
        RECT 243.040 56.870 243.255 57.380 ;
        RECT 243.485 56.870 243.765 57.200 ;
        RECT 243.945 56.870 244.185 57.380 ;
        RECT 240.440 55.800 241.865 55.970 ;
        RECT 239.955 55.000 240.490 55.620 ;
        RECT 240.660 54.830 240.990 55.630 ;
        RECT 241.475 55.625 241.865 55.800 ;
        RECT 242.255 55.620 242.570 56.640 ;
        RECT 242.740 55.970 242.910 56.470 ;
        RECT 243.160 56.140 243.425 56.700 ;
        RECT 243.595 55.970 243.765 56.870 ;
        RECT 243.935 56.140 244.290 56.700 ;
        RECT 244.555 56.640 245.170 57.210 ;
        RECT 245.340 56.870 245.555 57.380 ;
        RECT 245.785 56.870 246.065 57.200 ;
        RECT 246.245 56.870 246.485 57.380 ;
        RECT 242.740 55.800 244.165 55.970 ;
        RECT 242.255 55.000 242.790 55.620 ;
        RECT 242.960 54.830 243.290 55.630 ;
        RECT 243.775 55.625 244.165 55.800 ;
        RECT 244.555 55.620 244.870 56.640 ;
        RECT 245.040 55.970 245.210 56.470 ;
        RECT 245.460 56.140 245.725 56.700 ;
        RECT 245.895 55.970 246.065 56.870 ;
        RECT 246.235 56.140 246.590 56.700 ;
        RECT 246.820 56.610 250.330 57.380 ;
        RECT 251.425 56.830 251.680 57.120 ;
        RECT 251.850 57.000 252.180 57.380 ;
        RECT 251.425 56.660 252.175 56.830 ;
        RECT 246.820 56.090 248.470 56.610 ;
        RECT 245.040 55.800 246.465 55.970 ;
        RECT 248.640 55.920 250.330 56.440 ;
        RECT 244.555 55.000 245.090 55.620 ;
        RECT 245.260 54.830 245.590 55.630 ;
        RECT 246.075 55.625 246.465 55.800 ;
        RECT 246.820 54.830 250.330 55.920 ;
        RECT 251.425 55.840 251.775 56.490 ;
        RECT 251.945 55.670 252.175 56.660 ;
        RECT 251.425 55.500 252.175 55.670 ;
        RECT 251.425 55.000 251.680 55.500 ;
        RECT 251.850 54.830 252.180 55.330 ;
        RECT 252.350 55.000 252.520 57.120 ;
        RECT 252.880 57.020 253.210 57.380 ;
        RECT 253.380 56.990 253.875 57.160 ;
        RECT 254.080 56.990 254.935 57.160 ;
        RECT 252.750 55.800 253.210 56.850 ;
        RECT 252.690 55.015 253.015 55.800 ;
        RECT 253.380 55.630 253.550 56.990 ;
        RECT 253.720 56.080 254.070 56.700 ;
        RECT 254.240 56.480 254.595 56.700 ;
        RECT 254.240 55.890 254.410 56.480 ;
        RECT 254.765 56.280 254.935 56.990 ;
        RECT 255.810 56.920 256.140 57.380 ;
        RECT 256.350 57.020 256.700 57.190 ;
        RECT 255.140 56.450 255.930 56.700 ;
        RECT 256.350 56.630 256.610 57.020 ;
        RECT 256.920 56.930 257.870 57.210 ;
        RECT 258.040 56.940 258.230 57.380 ;
        RECT 258.400 57.000 259.470 57.170 ;
        RECT 256.100 56.280 256.270 56.460 ;
        RECT 253.380 55.460 253.775 55.630 ;
        RECT 253.945 55.500 254.410 55.890 ;
        RECT 254.580 56.110 256.270 56.280 ;
        RECT 253.605 55.330 253.775 55.460 ;
        RECT 254.580 55.330 254.750 56.110 ;
        RECT 256.440 55.940 256.610 56.630 ;
        RECT 255.110 55.770 256.610 55.940 ;
        RECT 256.800 55.970 257.010 56.760 ;
        RECT 257.180 56.140 257.530 56.760 ;
        RECT 257.700 56.150 257.870 56.930 ;
        RECT 258.400 56.770 258.570 57.000 ;
        RECT 258.040 56.600 258.570 56.770 ;
        RECT 258.040 56.320 258.260 56.600 ;
        RECT 258.740 56.430 258.980 56.830 ;
        RECT 257.700 55.980 258.105 56.150 ;
        RECT 258.440 56.060 258.980 56.430 ;
        RECT 259.150 56.645 259.470 57.000 ;
        RECT 259.715 56.920 260.020 57.380 ;
        RECT 260.190 56.670 260.445 57.200 ;
        RECT 261.290 56.690 261.620 57.380 ;
        RECT 262.080 56.785 262.700 57.210 ;
        RECT 262.870 56.890 263.200 57.380 ;
        RECT 259.150 56.470 259.475 56.645 ;
        RECT 259.150 56.170 260.065 56.470 ;
        RECT 259.325 56.140 260.065 56.170 ;
        RECT 256.800 55.810 257.475 55.970 ;
        RECT 257.935 55.890 258.105 55.980 ;
        RECT 256.800 55.800 257.765 55.810 ;
        RECT 256.440 55.630 256.610 55.770 ;
        RECT 253.185 54.830 253.435 55.290 ;
        RECT 253.605 55.000 253.855 55.330 ;
        RECT 254.070 55.000 254.750 55.330 ;
        RECT 254.920 55.430 255.995 55.600 ;
        RECT 256.440 55.460 257.000 55.630 ;
        RECT 257.305 55.510 257.765 55.800 ;
        RECT 257.935 55.720 259.155 55.890 ;
        RECT 254.920 55.090 255.090 55.430 ;
        RECT 255.325 54.830 255.655 55.260 ;
        RECT 255.825 55.090 255.995 55.430 ;
        RECT 256.290 54.830 256.660 55.290 ;
        RECT 256.830 55.000 257.000 55.460 ;
        RECT 257.935 55.340 258.105 55.720 ;
        RECT 259.325 55.550 259.495 56.140 ;
        RECT 260.235 56.020 260.445 56.670 ;
        RECT 262.340 56.450 262.700 56.785 ;
        RECT 257.235 55.000 258.105 55.340 ;
        RECT 258.695 55.380 259.495 55.550 ;
        RECT 258.275 54.830 258.525 55.290 ;
        RECT 258.695 55.090 258.865 55.380 ;
        RECT 259.045 54.830 259.375 55.210 ;
        RECT 259.715 54.830 260.020 55.970 ;
        RECT 260.190 55.140 260.445 56.020 ;
        RECT 261.280 56.170 262.700 56.450 ;
        RECT 260.750 54.830 261.080 56.000 ;
        RECT 261.280 55.000 261.610 56.170 ;
        RECT 261.810 54.830 262.140 56.000 ;
        RECT 262.340 55.000 262.700 56.170 ;
        RECT 262.870 56.140 263.210 56.720 ;
        RECT 263.380 56.610 265.050 57.380 ;
        RECT 265.220 56.655 265.510 57.380 ;
        RECT 265.680 56.640 266.065 57.210 ;
        RECT 266.235 56.920 266.560 57.380 ;
        RECT 267.080 56.750 267.360 57.210 ;
        RECT 263.380 56.090 264.130 56.610 ;
        RECT 262.870 54.830 263.200 55.970 ;
        RECT 264.300 55.920 265.050 56.440 ;
        RECT 263.380 54.830 265.050 55.920 ;
        RECT 265.220 54.830 265.510 55.995 ;
        RECT 265.680 55.970 265.960 56.640 ;
        RECT 266.235 56.580 267.360 56.750 ;
        RECT 266.235 56.470 266.685 56.580 ;
        RECT 266.130 56.140 266.685 56.470 ;
        RECT 267.550 56.410 267.950 57.210 ;
        RECT 268.350 56.920 268.620 57.380 ;
        RECT 268.790 56.750 269.075 57.210 ;
        RECT 269.360 56.835 274.705 57.380 ;
        RECT 265.680 55.000 266.065 55.970 ;
        RECT 266.235 55.680 266.685 56.140 ;
        RECT 266.855 55.850 267.950 56.410 ;
        RECT 266.235 55.460 267.360 55.680 ;
        RECT 266.235 54.830 266.560 55.290 ;
        RECT 267.080 55.000 267.360 55.460 ;
        RECT 267.550 55.000 267.950 55.850 ;
        RECT 268.120 56.580 269.075 56.750 ;
        RECT 268.120 55.680 268.330 56.580 ;
        RECT 268.500 55.850 269.190 56.410 ;
        RECT 270.945 56.005 271.285 56.835 ;
        RECT 274.885 56.670 275.140 57.200 ;
        RECT 275.310 56.920 275.615 57.380 ;
        RECT 275.860 57.000 276.930 57.170 ;
        RECT 268.120 55.460 269.075 55.680 ;
        RECT 268.350 54.830 268.620 55.290 ;
        RECT 268.790 55.000 269.075 55.460 ;
        RECT 272.765 55.265 273.115 56.515 ;
        RECT 274.885 56.020 275.095 56.670 ;
        RECT 275.860 56.645 276.180 57.000 ;
        RECT 275.855 56.470 276.180 56.645 ;
        RECT 275.265 56.170 276.180 56.470 ;
        RECT 276.350 56.430 276.590 56.830 ;
        RECT 276.760 56.770 276.930 57.000 ;
        RECT 277.100 56.940 277.290 57.380 ;
        RECT 277.460 56.930 278.410 57.210 ;
        RECT 278.630 57.020 278.980 57.190 ;
        RECT 276.760 56.600 277.290 56.770 ;
        RECT 275.265 56.140 276.005 56.170 ;
        RECT 269.360 54.830 274.705 55.265 ;
        RECT 274.885 55.140 275.140 56.020 ;
        RECT 275.310 54.830 275.615 55.970 ;
        RECT 275.835 55.550 276.005 56.140 ;
        RECT 276.350 56.060 276.890 56.430 ;
        RECT 277.070 56.320 277.290 56.600 ;
        RECT 277.460 56.150 277.630 56.930 ;
        RECT 277.225 55.980 277.630 56.150 ;
        RECT 277.800 56.140 278.150 56.760 ;
        RECT 277.225 55.890 277.395 55.980 ;
        RECT 278.320 55.970 278.530 56.760 ;
        RECT 276.175 55.720 277.395 55.890 ;
        RECT 277.855 55.810 278.530 55.970 ;
        RECT 275.835 55.380 276.635 55.550 ;
        RECT 275.955 54.830 276.285 55.210 ;
        RECT 276.465 55.090 276.635 55.380 ;
        RECT 277.225 55.340 277.395 55.720 ;
        RECT 277.565 55.800 278.530 55.810 ;
        RECT 278.720 56.630 278.980 57.020 ;
        RECT 279.190 56.920 279.520 57.380 ;
        RECT 280.395 56.990 281.250 57.160 ;
        RECT 281.455 56.990 281.950 57.160 ;
        RECT 282.120 57.020 282.450 57.380 ;
        RECT 278.720 55.940 278.890 56.630 ;
        RECT 279.060 56.280 279.230 56.460 ;
        RECT 279.400 56.450 280.190 56.700 ;
        RECT 280.395 56.280 280.565 56.990 ;
        RECT 280.735 56.480 281.090 56.700 ;
        RECT 279.060 56.110 280.750 56.280 ;
        RECT 277.565 55.510 278.025 55.800 ;
        RECT 278.720 55.770 280.220 55.940 ;
        RECT 278.720 55.630 278.890 55.770 ;
        RECT 278.330 55.460 278.890 55.630 ;
        RECT 276.805 54.830 277.055 55.290 ;
        RECT 277.225 55.000 278.095 55.340 ;
        RECT 278.330 55.000 278.500 55.460 ;
        RECT 279.335 55.430 280.410 55.600 ;
        RECT 278.670 54.830 279.040 55.290 ;
        RECT 279.335 55.090 279.505 55.430 ;
        RECT 279.675 54.830 280.005 55.260 ;
        RECT 280.240 55.090 280.410 55.430 ;
        RECT 280.580 55.330 280.750 56.110 ;
        RECT 280.920 55.890 281.090 56.480 ;
        RECT 281.260 56.080 281.610 56.700 ;
        RECT 280.920 55.500 281.385 55.890 ;
        RECT 281.780 55.630 281.950 56.990 ;
        RECT 282.120 55.800 282.580 56.850 ;
        RECT 281.555 55.460 281.950 55.630 ;
        RECT 281.555 55.330 281.725 55.460 ;
        RECT 280.580 55.000 281.260 55.330 ;
        RECT 281.475 55.000 281.725 55.330 ;
        RECT 281.895 54.830 282.145 55.290 ;
        RECT 282.315 55.015 282.640 55.800 ;
        RECT 282.810 55.000 282.980 57.120 ;
        RECT 283.150 57.000 283.480 57.380 ;
        RECT 283.650 56.830 283.905 57.120 ;
        RECT 283.155 56.660 283.905 56.830 ;
        RECT 283.155 55.670 283.385 56.660 ;
        RECT 284.080 56.630 285.290 57.380 ;
        RECT 285.705 56.900 286.005 57.380 ;
        RECT 286.175 56.730 286.435 57.185 ;
        RECT 286.605 56.900 286.865 57.380 ;
        RECT 287.035 56.730 287.295 57.185 ;
        RECT 287.465 56.900 287.725 57.380 ;
        RECT 287.895 56.730 288.155 57.185 ;
        RECT 288.325 56.900 288.585 57.380 ;
        RECT 288.755 56.730 289.015 57.185 ;
        RECT 289.185 56.855 289.445 57.380 ;
        RECT 283.555 55.840 283.905 56.490 ;
        RECT 284.080 56.090 284.600 56.630 ;
        RECT 285.705 56.560 289.015 56.730 ;
        RECT 284.770 55.920 285.290 56.460 ;
        RECT 283.155 55.500 283.905 55.670 ;
        RECT 283.150 54.830 283.480 55.330 ;
        RECT 283.650 55.000 283.905 55.500 ;
        RECT 284.080 54.830 285.290 55.920 ;
        RECT 285.705 55.970 286.675 56.560 ;
        RECT 289.615 56.390 289.865 57.200 ;
        RECT 290.045 56.920 290.290 57.380 ;
        RECT 286.845 56.140 289.865 56.390 ;
        RECT 290.035 56.140 290.350 56.750 ;
        RECT 290.980 56.655 291.270 57.380 ;
        RECT 291.500 56.920 291.745 57.380 ;
        RECT 291.440 56.140 291.755 56.750 ;
        RECT 291.925 56.390 292.175 57.200 ;
        RECT 292.345 56.855 292.605 57.380 ;
        RECT 292.775 56.730 293.035 57.185 ;
        RECT 293.205 56.900 293.465 57.380 ;
        RECT 293.635 56.730 293.895 57.185 ;
        RECT 294.065 56.900 294.325 57.380 ;
        RECT 294.495 56.730 294.755 57.185 ;
        RECT 294.925 56.900 295.185 57.380 ;
        RECT 295.355 56.730 295.615 57.185 ;
        RECT 295.785 56.900 296.085 57.380 ;
        RECT 292.775 56.560 296.085 56.730 ;
        RECT 291.925 56.140 294.945 56.390 ;
        RECT 285.705 55.730 289.015 55.970 ;
        RECT 285.710 54.830 286.005 55.560 ;
        RECT 286.175 55.005 286.435 55.730 ;
        RECT 286.605 54.830 286.865 55.560 ;
        RECT 287.035 55.005 287.295 55.730 ;
        RECT 287.465 54.830 287.725 55.560 ;
        RECT 287.895 55.005 288.155 55.730 ;
        RECT 288.325 54.830 288.585 55.560 ;
        RECT 288.755 55.005 289.015 55.730 ;
        RECT 289.185 54.830 289.445 55.940 ;
        RECT 289.615 55.005 289.865 56.140 ;
        RECT 290.045 54.830 290.340 55.940 ;
        RECT 290.980 54.830 291.270 55.995 ;
        RECT 291.450 54.830 291.745 55.940 ;
        RECT 291.925 55.005 292.175 56.140 ;
        RECT 295.115 55.970 296.085 56.560 ;
        RECT 296.500 56.610 299.090 57.380 ;
        RECT 299.810 56.830 299.980 57.120 ;
        RECT 300.150 57.000 300.480 57.380 ;
        RECT 299.810 56.660 300.475 56.830 ;
        RECT 296.500 56.090 297.710 56.610 ;
        RECT 292.345 54.830 292.605 55.940 ;
        RECT 292.775 55.730 296.085 55.970 ;
        RECT 297.880 55.920 299.090 56.440 ;
        RECT 292.775 55.005 293.035 55.730 ;
        RECT 293.205 54.830 293.465 55.560 ;
        RECT 293.635 55.005 293.895 55.730 ;
        RECT 294.065 54.830 294.325 55.560 ;
        RECT 294.495 55.005 294.755 55.730 ;
        RECT 294.925 54.830 295.185 55.560 ;
        RECT 295.355 55.005 295.615 55.730 ;
        RECT 295.785 54.830 296.080 55.560 ;
        RECT 296.500 54.830 299.090 55.920 ;
        RECT 299.725 55.840 300.075 56.490 ;
        RECT 300.245 55.670 300.475 56.660 ;
        RECT 299.810 55.500 300.475 55.670 ;
        RECT 299.810 55.000 299.980 55.500 ;
        RECT 300.150 54.830 300.480 55.330 ;
        RECT 300.650 55.000 300.875 57.120 ;
        RECT 301.090 57.000 301.420 57.380 ;
        RECT 301.590 56.830 301.760 57.160 ;
        RECT 302.060 57.000 303.075 57.200 ;
        RECT 301.065 56.640 301.760 56.830 ;
        RECT 301.065 55.670 301.235 56.640 ;
        RECT 301.405 55.840 301.815 56.460 ;
        RECT 301.985 55.890 302.205 56.760 ;
        RECT 302.385 56.450 302.735 56.820 ;
        RECT 302.905 56.270 303.075 57.000 ;
        RECT 303.245 56.940 303.655 57.380 ;
        RECT 303.945 56.740 304.195 57.170 ;
        RECT 304.395 56.920 304.715 57.380 ;
        RECT 305.275 56.990 306.125 57.160 ;
        RECT 303.245 56.400 303.655 56.730 ;
        RECT 303.945 56.400 304.365 56.740 ;
        RECT 302.655 56.230 303.075 56.270 ;
        RECT 302.655 56.060 304.005 56.230 ;
        RECT 301.065 55.500 301.760 55.670 ;
        RECT 301.985 55.510 302.485 55.890 ;
        RECT 301.090 54.830 301.420 55.330 ;
        RECT 301.590 55.000 301.760 55.500 ;
        RECT 302.655 55.215 302.825 56.060 ;
        RECT 303.755 55.900 304.005 56.060 ;
        RECT 302.995 55.630 303.245 55.890 ;
        RECT 304.175 55.630 304.365 56.400 ;
        RECT 302.995 55.380 304.365 55.630 ;
        RECT 304.535 56.570 305.785 56.740 ;
        RECT 304.535 55.810 304.705 56.570 ;
        RECT 305.455 56.450 305.785 56.570 ;
        RECT 304.875 55.990 305.055 56.400 ;
        RECT 305.955 56.230 306.125 56.990 ;
        RECT 306.325 56.900 306.985 57.380 ;
        RECT 307.165 56.785 307.485 57.115 ;
        RECT 306.315 56.460 306.975 56.730 ;
        RECT 306.315 56.400 306.645 56.460 ;
        RECT 306.795 56.230 307.125 56.290 ;
        RECT 305.225 56.060 307.125 56.230 ;
        RECT 304.535 55.500 305.055 55.810 ;
        RECT 305.225 55.550 305.395 56.060 ;
        RECT 307.295 55.890 307.485 56.785 ;
        RECT 305.565 55.720 307.485 55.890 ;
        RECT 307.165 55.700 307.485 55.720 ;
        RECT 307.685 56.470 307.935 57.120 ;
        RECT 308.115 56.920 308.400 57.380 ;
        RECT 308.580 56.670 308.835 57.200 ;
        RECT 307.685 56.140 308.485 56.470 ;
        RECT 305.225 55.380 306.435 55.550 ;
        RECT 301.995 55.045 302.825 55.215 ;
        RECT 303.065 54.830 303.445 55.210 ;
        RECT 303.625 55.090 303.795 55.380 ;
        RECT 305.225 55.300 305.395 55.380 ;
        RECT 303.965 54.830 304.295 55.210 ;
        RECT 304.765 55.050 305.395 55.300 ;
        RECT 305.575 54.830 305.995 55.210 ;
        RECT 306.195 55.090 306.435 55.380 ;
        RECT 306.665 54.830 306.995 55.520 ;
        RECT 307.165 55.090 307.335 55.700 ;
        RECT 307.685 55.550 307.935 56.140 ;
        RECT 308.655 55.810 308.835 56.670 ;
        RECT 309.840 56.630 311.050 57.380 ;
        RECT 307.605 55.040 307.935 55.550 ;
        RECT 308.115 54.830 308.400 55.630 ;
        RECT 308.580 55.340 308.835 55.810 ;
        RECT 309.840 55.920 310.360 56.460 ;
        RECT 310.530 56.090 311.050 56.630 ;
        RECT 308.580 55.170 308.920 55.340 ;
        RECT 308.580 55.140 308.835 55.170 ;
        RECT 309.840 54.830 311.050 55.920 ;
        RECT 162.095 54.660 311.135 54.830 ;
        RECT 162.180 53.570 163.390 54.660 ;
        RECT 163.560 53.570 165.230 54.660 ;
        RECT 165.865 53.990 166.120 54.490 ;
        RECT 166.290 54.160 166.620 54.660 ;
        RECT 165.865 53.820 166.615 53.990 ;
        RECT 162.180 52.860 162.700 53.400 ;
        RECT 162.870 53.030 163.390 53.570 ;
        RECT 163.560 52.880 164.310 53.400 ;
        RECT 164.480 53.050 165.230 53.570 ;
        RECT 165.865 53.000 166.215 53.650 ;
        RECT 162.180 52.110 163.390 52.860 ;
        RECT 163.560 52.110 165.230 52.880 ;
        RECT 166.385 52.830 166.615 53.820 ;
        RECT 165.865 52.660 166.615 52.830 ;
        RECT 165.865 52.370 166.120 52.660 ;
        RECT 166.290 52.110 166.620 52.490 ;
        RECT 166.790 52.370 166.960 54.490 ;
        RECT 167.130 53.690 167.455 54.475 ;
        RECT 167.625 54.200 167.875 54.660 ;
        RECT 168.045 54.160 168.295 54.490 ;
        RECT 168.510 54.160 169.190 54.490 ;
        RECT 168.045 54.030 168.215 54.160 ;
        RECT 167.820 53.860 168.215 54.030 ;
        RECT 167.190 52.640 167.650 53.690 ;
        RECT 167.820 52.500 167.990 53.860 ;
        RECT 168.385 53.600 168.850 53.990 ;
        RECT 168.160 52.790 168.510 53.410 ;
        RECT 168.680 53.010 168.850 53.600 ;
        RECT 169.020 53.380 169.190 54.160 ;
        RECT 169.360 54.060 169.530 54.400 ;
        RECT 169.765 54.230 170.095 54.660 ;
        RECT 170.265 54.060 170.435 54.400 ;
        RECT 170.730 54.200 171.100 54.660 ;
        RECT 169.360 53.890 170.435 54.060 ;
        RECT 171.270 54.030 171.440 54.490 ;
        RECT 171.675 54.150 172.545 54.490 ;
        RECT 172.715 54.200 172.965 54.660 ;
        RECT 170.880 53.860 171.440 54.030 ;
        RECT 170.880 53.720 171.050 53.860 ;
        RECT 169.550 53.550 171.050 53.720 ;
        RECT 171.745 53.690 172.205 53.980 ;
        RECT 169.020 53.210 170.710 53.380 ;
        RECT 168.680 52.790 169.035 53.010 ;
        RECT 169.205 52.500 169.375 53.210 ;
        RECT 169.580 52.790 170.370 53.040 ;
        RECT 170.540 53.030 170.710 53.210 ;
        RECT 170.880 52.860 171.050 53.550 ;
        RECT 167.320 52.110 167.650 52.470 ;
        RECT 167.820 52.330 168.315 52.500 ;
        RECT 168.520 52.330 169.375 52.500 ;
        RECT 170.250 52.110 170.580 52.570 ;
        RECT 170.790 52.470 171.050 52.860 ;
        RECT 171.240 53.680 172.205 53.690 ;
        RECT 172.375 53.770 172.545 54.150 ;
        RECT 173.135 54.110 173.305 54.400 ;
        RECT 173.485 54.280 173.815 54.660 ;
        RECT 173.135 53.940 173.935 54.110 ;
        RECT 171.240 53.520 171.915 53.680 ;
        RECT 172.375 53.600 173.595 53.770 ;
        RECT 171.240 52.730 171.450 53.520 ;
        RECT 172.375 53.510 172.545 53.600 ;
        RECT 171.620 52.730 171.970 53.350 ;
        RECT 172.140 53.340 172.545 53.510 ;
        RECT 172.140 52.560 172.310 53.340 ;
        RECT 172.480 52.890 172.700 53.170 ;
        RECT 172.880 53.060 173.420 53.430 ;
        RECT 173.765 53.350 173.935 53.940 ;
        RECT 174.155 53.520 174.460 54.660 ;
        RECT 174.630 53.470 174.885 54.350 ;
        RECT 175.060 53.495 175.350 54.660 ;
        RECT 175.520 53.690 175.830 54.490 ;
        RECT 176.000 53.860 176.310 54.660 ;
        RECT 176.480 54.030 176.740 54.490 ;
        RECT 176.910 54.200 177.165 54.660 ;
        RECT 177.340 54.030 177.600 54.490 ;
        RECT 176.480 53.860 177.600 54.030 ;
        RECT 176.960 53.810 177.130 53.860 ;
        RECT 175.520 53.520 176.550 53.690 ;
        RECT 173.765 53.320 174.505 53.350 ;
        RECT 172.480 52.720 173.010 52.890 ;
        RECT 170.790 52.300 171.140 52.470 ;
        RECT 171.360 52.280 172.310 52.560 ;
        RECT 172.480 52.110 172.670 52.550 ;
        RECT 172.840 52.490 173.010 52.720 ;
        RECT 173.180 52.660 173.420 53.060 ;
        RECT 173.590 53.020 174.505 53.320 ;
        RECT 173.590 52.845 173.915 53.020 ;
        RECT 173.590 52.490 173.910 52.845 ;
        RECT 174.675 52.820 174.885 53.470 ;
        RECT 172.840 52.320 173.910 52.490 ;
        RECT 174.155 52.110 174.460 52.570 ;
        RECT 174.630 52.290 174.885 52.820 ;
        RECT 175.060 52.110 175.350 52.835 ;
        RECT 175.520 52.610 175.690 53.520 ;
        RECT 175.860 52.780 176.210 53.350 ;
        RECT 176.380 53.270 176.550 53.520 ;
        RECT 177.340 53.610 177.600 53.860 ;
        RECT 177.770 53.790 178.055 54.660 ;
        RECT 178.280 54.225 183.625 54.660 ;
        RECT 184.265 54.280 184.600 54.660 ;
        RECT 177.340 53.440 178.095 53.610 ;
        RECT 176.380 53.100 177.520 53.270 ;
        RECT 177.690 52.930 178.095 53.440 ;
        RECT 176.445 52.760 178.095 52.930 ;
        RECT 175.520 52.280 175.820 52.610 ;
        RECT 175.990 52.110 176.265 52.590 ;
        RECT 176.445 52.370 176.740 52.760 ;
        RECT 176.910 52.110 177.165 52.590 ;
        RECT 177.340 52.370 177.600 52.760 ;
        RECT 179.865 52.655 180.205 53.485 ;
        RECT 181.685 52.975 182.035 54.225 ;
        RECT 184.260 52.790 184.500 54.100 ;
        RECT 184.770 53.690 185.020 54.490 ;
        RECT 185.240 53.940 185.570 54.660 ;
        RECT 185.755 53.690 186.005 54.490 ;
        RECT 186.470 53.860 186.800 54.660 ;
        RECT 186.970 54.230 187.310 54.490 ;
        RECT 184.670 53.520 186.860 53.690 ;
        RECT 177.770 52.110 178.050 52.590 ;
        RECT 178.280 52.110 183.625 52.655 ;
        RECT 184.670 52.610 184.840 53.520 ;
        RECT 186.545 53.350 186.860 53.520 ;
        RECT 184.345 52.280 184.840 52.610 ;
        RECT 185.060 52.385 185.410 53.350 ;
        RECT 185.590 52.380 185.890 53.350 ;
        RECT 186.070 52.380 186.350 53.350 ;
        RECT 186.545 53.100 186.875 53.350 ;
        RECT 186.530 52.110 186.800 52.910 ;
        RECT 187.050 52.830 187.310 54.230 ;
        RECT 187.480 54.150 187.740 54.660 ;
        RECT 187.480 53.100 187.820 53.980 ;
        RECT 187.990 53.270 188.160 54.490 ;
        RECT 188.400 54.155 189.015 54.660 ;
        RECT 188.400 53.620 188.650 53.985 ;
        RECT 188.820 53.980 189.015 54.155 ;
        RECT 189.185 54.150 189.660 54.490 ;
        RECT 189.830 54.115 190.045 54.660 ;
        RECT 188.820 53.790 189.150 53.980 ;
        RECT 189.370 53.620 190.085 53.915 ;
        RECT 190.255 53.790 190.530 54.490 ;
        RECT 191.000 54.020 191.330 54.450 ;
        RECT 188.400 53.450 190.190 53.620 ;
        RECT 187.990 53.020 188.785 53.270 ;
        RECT 187.990 52.930 188.240 53.020 ;
        RECT 186.970 52.320 187.310 52.830 ;
        RECT 187.480 52.110 187.740 52.930 ;
        RECT 187.910 52.510 188.240 52.930 ;
        RECT 188.955 52.595 189.210 53.450 ;
        RECT 188.420 52.330 189.210 52.595 ;
        RECT 189.380 52.750 189.790 53.270 ;
        RECT 189.960 53.020 190.190 53.450 ;
        RECT 190.360 52.760 190.530 53.790 ;
        RECT 189.380 52.330 189.580 52.750 ;
        RECT 189.770 52.110 190.100 52.570 ;
        RECT 190.270 52.280 190.530 52.760 ;
        RECT 190.875 53.850 191.330 54.020 ;
        RECT 191.510 54.020 191.760 54.440 ;
        RECT 191.990 54.190 192.320 54.660 ;
        RECT 192.550 54.020 192.800 54.440 ;
        RECT 191.510 53.850 192.800 54.020 ;
        RECT 190.875 52.850 191.045 53.850 ;
        RECT 191.215 53.020 191.460 53.680 ;
        RECT 191.675 53.020 191.940 53.680 ;
        RECT 192.135 53.020 192.420 53.680 ;
        RECT 192.595 53.350 192.810 53.680 ;
        RECT 192.990 53.520 193.240 54.660 ;
        RECT 193.410 53.600 193.740 54.450 ;
        RECT 195.040 53.990 195.320 54.660 ;
        RECT 195.490 53.770 195.790 54.320 ;
        RECT 195.990 53.940 196.320 54.660 ;
        RECT 196.510 53.940 196.970 54.490 ;
        RECT 193.520 53.470 193.740 53.600 ;
        RECT 192.595 53.020 192.900 53.350 ;
        RECT 193.070 53.020 193.380 53.350 ;
        RECT 193.070 52.850 193.240 53.020 ;
        RECT 190.875 52.680 193.240 52.850 ;
        RECT 193.550 52.835 193.740 53.470 ;
        RECT 194.855 53.350 195.120 53.710 ;
        RECT 195.490 53.600 196.430 53.770 ;
        RECT 196.260 53.350 196.430 53.600 ;
        RECT 194.855 53.100 195.530 53.350 ;
        RECT 195.750 53.100 196.090 53.350 ;
        RECT 196.260 53.020 196.550 53.350 ;
        RECT 196.260 52.930 196.430 53.020 ;
        RECT 191.030 52.110 191.360 52.510 ;
        RECT 191.530 52.340 191.860 52.680 ;
        RECT 192.910 52.110 193.240 52.510 ;
        RECT 193.410 52.325 193.740 52.835 ;
        RECT 195.040 52.740 196.430 52.930 ;
        RECT 195.040 52.380 195.370 52.740 ;
        RECT 196.720 52.570 196.970 53.940 ;
        RECT 197.140 53.520 197.400 54.660 ;
        RECT 197.570 53.690 197.900 54.490 ;
        RECT 198.070 53.860 198.240 54.660 ;
        RECT 198.410 53.690 198.740 54.490 ;
        RECT 198.910 53.860 199.165 54.660 ;
        RECT 197.570 53.520 199.270 53.690 ;
        RECT 199.440 53.570 200.650 54.660 ;
        RECT 197.140 53.100 197.900 53.350 ;
        RECT 198.070 53.100 198.820 53.350 ;
        RECT 198.990 52.930 199.270 53.520 ;
        RECT 195.990 52.110 196.240 52.570 ;
        RECT 196.410 52.280 196.970 52.570 ;
        RECT 197.140 52.740 198.240 52.910 ;
        RECT 197.140 52.280 197.480 52.740 ;
        RECT 197.650 52.110 197.820 52.570 ;
        RECT 197.990 52.490 198.240 52.740 ;
        RECT 198.410 52.680 199.270 52.930 ;
        RECT 199.440 52.860 199.960 53.400 ;
        RECT 200.130 53.030 200.650 53.570 ;
        RECT 200.820 53.495 201.110 54.660 ;
        RECT 201.280 53.570 202.490 54.660 ;
        RECT 201.280 52.860 201.800 53.400 ;
        RECT 201.970 53.030 202.490 53.570 ;
        RECT 202.845 53.690 203.235 53.865 ;
        RECT 203.720 53.860 204.050 54.660 ;
        RECT 204.220 53.870 204.755 54.490 ;
        RECT 202.845 53.520 204.270 53.690 ;
        RECT 198.830 52.490 199.160 52.510 ;
        RECT 197.990 52.280 199.160 52.490 ;
        RECT 199.440 52.110 200.650 52.860 ;
        RECT 200.820 52.110 201.110 52.835 ;
        RECT 201.280 52.110 202.490 52.860 ;
        RECT 202.720 52.790 203.075 53.350 ;
        RECT 203.245 52.620 203.415 53.520 ;
        RECT 203.585 52.790 203.850 53.350 ;
        RECT 204.100 53.020 204.270 53.520 ;
        RECT 204.440 52.850 204.755 53.870 ;
        RECT 204.960 53.570 208.470 54.660 ;
        RECT 202.825 52.110 203.065 52.620 ;
        RECT 203.245 52.290 203.525 52.620 ;
        RECT 203.755 52.110 203.970 52.620 ;
        RECT 204.140 52.280 204.755 52.850 ;
        RECT 204.960 52.880 206.610 53.400 ;
        RECT 206.780 53.050 208.470 53.570 ;
        RECT 208.825 53.690 209.215 53.865 ;
        RECT 209.700 53.860 210.030 54.660 ;
        RECT 210.200 53.870 210.735 54.490 ;
        RECT 208.825 53.520 210.250 53.690 ;
        RECT 204.960 52.110 208.470 52.880 ;
        RECT 208.700 52.790 209.055 53.350 ;
        RECT 209.225 52.620 209.395 53.520 ;
        RECT 209.565 52.790 209.830 53.350 ;
        RECT 210.080 53.020 210.250 53.520 ;
        RECT 210.420 52.850 210.735 53.870 ;
        RECT 210.945 53.990 211.200 54.490 ;
        RECT 211.370 54.160 211.700 54.660 ;
        RECT 210.945 53.820 211.695 53.990 ;
        RECT 210.945 53.000 211.295 53.650 ;
        RECT 208.805 52.110 209.045 52.620 ;
        RECT 209.225 52.290 209.505 52.620 ;
        RECT 209.735 52.110 209.950 52.620 ;
        RECT 210.120 52.280 210.735 52.850 ;
        RECT 211.465 52.830 211.695 53.820 ;
        RECT 210.945 52.660 211.695 52.830 ;
        RECT 210.945 52.370 211.200 52.660 ;
        RECT 211.370 52.110 211.700 52.490 ;
        RECT 211.870 52.370 212.040 54.490 ;
        RECT 212.210 53.690 212.535 54.475 ;
        RECT 212.705 54.200 212.955 54.660 ;
        RECT 213.125 54.160 213.375 54.490 ;
        RECT 213.590 54.160 214.270 54.490 ;
        RECT 213.125 54.030 213.295 54.160 ;
        RECT 212.900 53.860 213.295 54.030 ;
        RECT 212.270 52.640 212.730 53.690 ;
        RECT 212.900 52.500 213.070 53.860 ;
        RECT 213.465 53.600 213.930 53.990 ;
        RECT 213.240 52.790 213.590 53.410 ;
        RECT 213.760 53.010 213.930 53.600 ;
        RECT 214.100 53.380 214.270 54.160 ;
        RECT 214.440 54.060 214.610 54.400 ;
        RECT 214.845 54.230 215.175 54.660 ;
        RECT 215.345 54.060 215.515 54.400 ;
        RECT 215.810 54.200 216.180 54.660 ;
        RECT 214.440 53.890 215.515 54.060 ;
        RECT 216.350 54.030 216.520 54.490 ;
        RECT 216.755 54.150 217.625 54.490 ;
        RECT 217.795 54.200 218.045 54.660 ;
        RECT 215.960 53.860 216.520 54.030 ;
        RECT 215.960 53.720 216.130 53.860 ;
        RECT 214.630 53.550 216.130 53.720 ;
        RECT 216.825 53.690 217.285 53.980 ;
        RECT 214.100 53.210 215.790 53.380 ;
        RECT 213.760 52.790 214.115 53.010 ;
        RECT 214.285 52.500 214.455 53.210 ;
        RECT 214.660 52.790 215.450 53.040 ;
        RECT 215.620 53.030 215.790 53.210 ;
        RECT 215.960 52.860 216.130 53.550 ;
        RECT 212.400 52.110 212.730 52.470 ;
        RECT 212.900 52.330 213.395 52.500 ;
        RECT 213.600 52.330 214.455 52.500 ;
        RECT 215.330 52.110 215.660 52.570 ;
        RECT 215.870 52.470 216.130 52.860 ;
        RECT 216.320 53.680 217.285 53.690 ;
        RECT 217.455 53.770 217.625 54.150 ;
        RECT 218.215 54.110 218.385 54.400 ;
        RECT 218.565 54.280 218.895 54.660 ;
        RECT 218.215 53.940 219.015 54.110 ;
        RECT 216.320 53.520 216.995 53.680 ;
        RECT 217.455 53.600 218.675 53.770 ;
        RECT 216.320 52.730 216.530 53.520 ;
        RECT 217.455 53.510 217.625 53.600 ;
        RECT 216.700 52.730 217.050 53.350 ;
        RECT 217.220 53.340 217.625 53.510 ;
        RECT 217.220 52.560 217.390 53.340 ;
        RECT 217.560 52.890 217.780 53.170 ;
        RECT 217.960 53.060 218.500 53.430 ;
        RECT 218.845 53.350 219.015 53.940 ;
        RECT 219.235 53.520 219.540 54.660 ;
        RECT 219.710 53.470 219.965 54.350 ;
        RECT 220.140 53.570 221.350 54.660 ;
        RECT 221.770 53.930 222.065 54.660 ;
        RECT 222.235 53.760 222.495 54.485 ;
        RECT 222.665 53.930 222.925 54.660 ;
        RECT 223.095 53.760 223.355 54.485 ;
        RECT 223.525 53.930 223.785 54.660 ;
        RECT 223.955 53.760 224.215 54.485 ;
        RECT 224.385 53.930 224.645 54.660 ;
        RECT 224.815 53.760 225.075 54.485 ;
        RECT 218.845 53.320 219.585 53.350 ;
        RECT 217.560 52.720 218.090 52.890 ;
        RECT 215.870 52.300 216.220 52.470 ;
        RECT 216.440 52.280 217.390 52.560 ;
        RECT 217.560 52.110 217.750 52.550 ;
        RECT 217.920 52.490 218.090 52.720 ;
        RECT 218.260 52.660 218.500 53.060 ;
        RECT 218.670 53.020 219.585 53.320 ;
        RECT 218.670 52.845 218.995 53.020 ;
        RECT 218.670 52.490 218.990 52.845 ;
        RECT 219.755 52.820 219.965 53.470 ;
        RECT 217.920 52.320 218.990 52.490 ;
        RECT 219.235 52.110 219.540 52.570 ;
        RECT 219.710 52.290 219.965 52.820 ;
        RECT 220.140 52.860 220.660 53.400 ;
        RECT 220.830 53.030 221.350 53.570 ;
        RECT 221.765 53.520 225.075 53.760 ;
        RECT 225.245 53.550 225.505 54.660 ;
        RECT 221.765 52.930 222.735 53.520 ;
        RECT 225.675 53.350 225.925 54.485 ;
        RECT 226.105 53.550 226.400 54.660 ;
        RECT 226.580 53.495 226.870 54.660 ;
        RECT 227.050 53.550 227.345 54.660 ;
        RECT 227.525 53.350 227.775 54.485 ;
        RECT 227.945 53.550 228.205 54.660 ;
        RECT 228.375 53.760 228.635 54.485 ;
        RECT 228.805 53.930 229.065 54.660 ;
        RECT 229.235 53.760 229.495 54.485 ;
        RECT 229.665 53.930 229.925 54.660 ;
        RECT 230.095 53.760 230.355 54.485 ;
        RECT 230.525 53.930 230.785 54.660 ;
        RECT 230.955 53.760 231.215 54.485 ;
        RECT 231.385 53.930 231.680 54.660 ;
        RECT 228.375 53.520 231.685 53.760 ;
        RECT 232.285 53.690 232.675 53.865 ;
        RECT 233.160 53.860 233.490 54.660 ;
        RECT 233.660 53.870 234.195 54.490 ;
        RECT 232.285 53.520 233.710 53.690 ;
        RECT 222.905 53.100 225.925 53.350 ;
        RECT 220.140 52.110 221.350 52.860 ;
        RECT 221.765 52.760 225.075 52.930 ;
        RECT 221.765 52.110 222.065 52.590 ;
        RECT 222.235 52.305 222.495 52.760 ;
        RECT 222.665 52.110 222.925 52.590 ;
        RECT 223.095 52.305 223.355 52.760 ;
        RECT 223.525 52.110 223.785 52.590 ;
        RECT 223.955 52.305 224.215 52.760 ;
        RECT 224.385 52.110 224.645 52.590 ;
        RECT 224.815 52.305 225.075 52.760 ;
        RECT 225.245 52.110 225.505 52.635 ;
        RECT 225.675 52.290 225.925 53.100 ;
        RECT 226.095 52.740 226.410 53.350 ;
        RECT 226.105 52.110 226.350 52.570 ;
        RECT 226.580 52.110 226.870 52.835 ;
        RECT 227.040 52.740 227.355 53.350 ;
        RECT 227.525 53.100 230.545 53.350 ;
        RECT 227.100 52.110 227.345 52.570 ;
        RECT 227.525 52.290 227.775 53.100 ;
        RECT 230.715 52.930 231.685 53.520 ;
        RECT 228.375 52.760 231.685 52.930 ;
        RECT 232.160 52.790 232.515 53.350 ;
        RECT 227.945 52.110 228.205 52.635 ;
        RECT 228.375 52.305 228.635 52.760 ;
        RECT 228.805 52.110 229.065 52.590 ;
        RECT 229.235 52.305 229.495 52.760 ;
        RECT 229.665 52.110 229.925 52.590 ;
        RECT 230.095 52.305 230.355 52.760 ;
        RECT 230.525 52.110 230.785 52.590 ;
        RECT 230.955 52.305 231.215 52.760 ;
        RECT 232.685 52.620 232.855 53.520 ;
        RECT 233.025 52.790 233.290 53.350 ;
        RECT 233.540 53.020 233.710 53.520 ;
        RECT 233.880 52.850 234.195 53.870 ;
        RECT 231.385 52.110 231.685 52.590 ;
        RECT 232.265 52.110 232.505 52.620 ;
        RECT 232.685 52.290 232.965 52.620 ;
        RECT 233.195 52.110 233.410 52.620 ;
        RECT 233.580 52.280 234.195 52.850 ;
        RECT 235.320 53.900 235.985 54.490 ;
        RECT 235.320 52.930 235.570 53.900 ;
        RECT 236.155 53.820 236.485 54.660 ;
        RECT 236.995 54.070 237.800 54.490 ;
        RECT 236.655 53.900 238.220 54.070 ;
        RECT 236.655 53.650 236.825 53.900 ;
        RECT 235.905 53.480 236.825 53.650 ;
        RECT 235.905 53.310 236.075 53.480 ;
        RECT 236.995 53.310 237.370 53.730 ;
        RECT 235.740 53.100 236.075 53.310 ;
        RECT 236.245 53.100 236.695 53.310 ;
        RECT 236.885 53.300 237.370 53.310 ;
        RECT 237.560 53.350 237.880 53.730 ;
        RECT 238.050 53.650 238.220 53.900 ;
        RECT 238.390 53.820 238.640 54.660 ;
        RECT 238.835 53.650 239.135 54.490 ;
        RECT 238.050 53.480 239.135 53.650 ;
        RECT 239.460 53.570 240.670 54.660 ;
        RECT 236.885 53.130 237.390 53.300 ;
        RECT 236.885 53.100 237.370 53.130 ;
        RECT 237.560 53.100 237.940 53.350 ;
        RECT 238.120 53.100 238.450 53.310 ;
        RECT 235.320 52.290 236.005 52.930 ;
        RECT 236.175 52.110 236.345 52.930 ;
        RECT 236.515 52.760 238.215 52.930 ;
        RECT 236.515 52.295 236.845 52.760 ;
        RECT 237.830 52.670 238.215 52.760 ;
        RECT 238.620 52.850 238.790 53.480 ;
        RECT 238.960 53.020 239.290 53.310 ;
        RECT 239.460 52.860 239.980 53.400 ;
        RECT 240.150 53.030 240.670 53.570 ;
        RECT 240.840 53.520 241.225 54.490 ;
        RECT 241.395 54.200 241.720 54.660 ;
        RECT 242.240 54.030 242.520 54.490 ;
        RECT 241.395 53.810 242.520 54.030 ;
        RECT 238.620 52.670 239.130 52.850 ;
        RECT 237.015 52.110 237.185 52.580 ;
        RECT 237.445 52.330 238.630 52.500 ;
        RECT 238.800 52.280 239.130 52.670 ;
        RECT 239.460 52.110 240.670 52.860 ;
        RECT 240.840 52.850 241.120 53.520 ;
        RECT 241.395 53.350 241.845 53.810 ;
        RECT 242.710 53.640 243.110 54.490 ;
        RECT 243.510 54.200 243.780 54.660 ;
        RECT 243.950 54.030 244.235 54.490 ;
        RECT 244.620 54.200 244.790 54.660 ;
        RECT 241.290 53.020 241.845 53.350 ;
        RECT 242.015 53.080 243.110 53.640 ;
        RECT 241.395 52.910 241.845 53.020 ;
        RECT 240.840 52.280 241.225 52.850 ;
        RECT 241.395 52.740 242.520 52.910 ;
        RECT 241.395 52.110 241.720 52.570 ;
        RECT 242.240 52.280 242.520 52.740 ;
        RECT 242.710 52.280 243.110 53.080 ;
        RECT 243.280 53.810 244.235 54.030 ;
        RECT 243.280 52.910 243.490 53.810 ;
        RECT 244.960 53.710 245.290 54.490 ;
        RECT 245.460 53.860 245.630 54.660 ;
        RECT 244.520 53.690 245.290 53.710 ;
        RECT 245.800 53.690 246.130 54.490 ;
        RECT 246.300 53.860 246.470 54.660 ;
        RECT 246.640 53.690 246.970 54.490 ;
        RECT 243.660 53.080 244.350 53.640 ;
        RECT 244.520 53.520 246.970 53.690 ;
        RECT 247.230 53.520 247.525 54.660 ;
        RECT 247.855 54.030 248.140 54.490 ;
        RECT 248.310 54.200 248.580 54.660 ;
        RECT 247.855 53.810 248.810 54.030 ;
        RECT 244.520 52.930 244.870 53.520 ;
        RECT 245.040 53.100 247.550 53.350 ;
        RECT 247.740 53.080 248.430 53.640 ;
        RECT 243.280 52.740 244.235 52.910 ;
        RECT 244.520 52.750 246.890 52.930 ;
        RECT 248.600 52.910 248.810 53.810 ;
        RECT 243.510 52.110 243.780 52.570 ;
        RECT 243.950 52.280 244.235 52.740 ;
        RECT 244.620 52.110 244.870 52.575 ;
        RECT 245.040 52.280 245.210 52.750 ;
        RECT 245.460 52.110 245.630 52.570 ;
        RECT 245.880 52.280 246.050 52.750 ;
        RECT 246.300 52.110 246.470 52.570 ;
        RECT 246.720 52.280 246.890 52.750 ;
        RECT 247.855 52.740 248.810 52.910 ;
        RECT 248.980 53.640 249.380 54.490 ;
        RECT 249.570 54.030 249.850 54.490 ;
        RECT 250.370 54.200 250.695 54.660 ;
        RECT 249.570 53.810 250.695 54.030 ;
        RECT 248.980 53.080 250.075 53.640 ;
        RECT 250.245 53.350 250.695 53.810 ;
        RECT 250.865 53.520 251.250 54.490 ;
        RECT 247.260 52.110 247.525 52.570 ;
        RECT 247.855 52.280 248.140 52.740 ;
        RECT 248.310 52.110 248.580 52.570 ;
        RECT 248.980 52.280 249.380 53.080 ;
        RECT 250.245 53.020 250.800 53.350 ;
        RECT 250.245 52.910 250.695 53.020 ;
        RECT 249.570 52.740 250.695 52.910 ;
        RECT 250.970 52.850 251.250 53.520 ;
        RECT 252.340 53.495 252.630 54.660 ;
        RECT 252.835 53.870 253.370 54.490 ;
        RECT 249.570 52.280 249.850 52.740 ;
        RECT 250.370 52.110 250.695 52.570 ;
        RECT 250.865 52.280 251.250 52.850 ;
        RECT 252.835 52.850 253.150 53.870 ;
        RECT 253.540 53.860 253.870 54.660 ;
        RECT 254.355 53.690 254.745 53.865 ;
        RECT 253.320 53.520 254.745 53.690 ;
        RECT 255.110 53.550 255.405 54.660 ;
        RECT 253.320 53.020 253.490 53.520 ;
        RECT 252.340 52.110 252.630 52.835 ;
        RECT 252.835 52.280 253.450 52.850 ;
        RECT 253.740 52.790 254.005 53.350 ;
        RECT 254.175 52.620 254.345 53.520 ;
        RECT 255.585 53.350 255.835 54.485 ;
        RECT 256.005 53.550 256.265 54.660 ;
        RECT 256.435 53.760 256.695 54.485 ;
        RECT 256.865 53.930 257.125 54.660 ;
        RECT 257.295 53.760 257.555 54.485 ;
        RECT 257.725 53.930 257.985 54.660 ;
        RECT 258.155 53.760 258.415 54.485 ;
        RECT 258.585 53.930 258.845 54.660 ;
        RECT 259.015 53.760 259.275 54.485 ;
        RECT 259.445 53.930 259.740 54.660 ;
        RECT 256.435 53.520 259.745 53.760 ;
        RECT 254.515 52.790 254.870 53.350 ;
        RECT 255.100 52.740 255.415 53.350 ;
        RECT 255.585 53.100 258.605 53.350 ;
        RECT 253.620 52.110 253.835 52.620 ;
        RECT 254.065 52.290 254.345 52.620 ;
        RECT 254.525 52.110 254.765 52.620 ;
        RECT 255.160 52.110 255.405 52.570 ;
        RECT 255.585 52.290 255.835 53.100 ;
        RECT 258.775 52.930 259.745 53.520 ;
        RECT 256.435 52.760 259.745 52.930 ;
        RECT 261.085 53.470 261.340 54.350 ;
        RECT 261.510 53.520 261.815 54.660 ;
        RECT 262.155 54.280 262.485 54.660 ;
        RECT 262.665 54.110 262.835 54.400 ;
        RECT 263.005 54.200 263.255 54.660 ;
        RECT 262.035 53.940 262.835 54.110 ;
        RECT 263.425 54.150 264.295 54.490 ;
        RECT 261.085 52.820 261.295 53.470 ;
        RECT 262.035 53.350 262.205 53.940 ;
        RECT 263.425 53.770 263.595 54.150 ;
        RECT 264.530 54.030 264.700 54.490 ;
        RECT 264.870 54.200 265.240 54.660 ;
        RECT 265.535 54.060 265.705 54.400 ;
        RECT 265.875 54.230 266.205 54.660 ;
        RECT 266.440 54.060 266.610 54.400 ;
        RECT 262.375 53.600 263.595 53.770 ;
        RECT 263.765 53.690 264.225 53.980 ;
        RECT 264.530 53.860 265.090 54.030 ;
        RECT 265.535 53.890 266.610 54.060 ;
        RECT 266.780 54.160 267.460 54.490 ;
        RECT 267.675 54.160 267.925 54.490 ;
        RECT 268.095 54.200 268.345 54.660 ;
        RECT 264.920 53.720 265.090 53.860 ;
        RECT 263.765 53.680 264.730 53.690 ;
        RECT 263.425 53.510 263.595 53.600 ;
        RECT 264.055 53.520 264.730 53.680 ;
        RECT 261.465 53.320 262.205 53.350 ;
        RECT 261.465 53.020 262.380 53.320 ;
        RECT 262.055 52.845 262.380 53.020 ;
        RECT 256.005 52.110 256.265 52.635 ;
        RECT 256.435 52.305 256.695 52.760 ;
        RECT 256.865 52.110 257.125 52.590 ;
        RECT 257.295 52.305 257.555 52.760 ;
        RECT 257.725 52.110 257.985 52.590 ;
        RECT 258.155 52.305 258.415 52.760 ;
        RECT 258.585 52.110 258.845 52.590 ;
        RECT 259.015 52.305 259.275 52.760 ;
        RECT 259.445 52.110 259.745 52.590 ;
        RECT 261.085 52.290 261.340 52.820 ;
        RECT 261.510 52.110 261.815 52.570 ;
        RECT 262.060 52.490 262.380 52.845 ;
        RECT 262.550 53.060 263.090 53.430 ;
        RECT 263.425 53.340 263.830 53.510 ;
        RECT 262.550 52.660 262.790 53.060 ;
        RECT 263.270 52.890 263.490 53.170 ;
        RECT 262.960 52.720 263.490 52.890 ;
        RECT 262.960 52.490 263.130 52.720 ;
        RECT 263.660 52.560 263.830 53.340 ;
        RECT 264.000 52.730 264.350 53.350 ;
        RECT 264.520 52.730 264.730 53.520 ;
        RECT 264.920 53.550 266.420 53.720 ;
        RECT 264.920 52.860 265.090 53.550 ;
        RECT 266.780 53.380 266.950 54.160 ;
        RECT 267.755 54.030 267.925 54.160 ;
        RECT 265.260 53.210 266.950 53.380 ;
        RECT 267.120 53.600 267.585 53.990 ;
        RECT 267.755 53.860 268.150 54.030 ;
        RECT 265.260 53.030 265.430 53.210 ;
        RECT 262.060 52.320 263.130 52.490 ;
        RECT 263.300 52.110 263.490 52.550 ;
        RECT 263.660 52.280 264.610 52.560 ;
        RECT 264.920 52.470 265.180 52.860 ;
        RECT 265.600 52.790 266.390 53.040 ;
        RECT 264.830 52.300 265.180 52.470 ;
        RECT 265.390 52.110 265.720 52.570 ;
        RECT 266.595 52.500 266.765 53.210 ;
        RECT 267.120 53.010 267.290 53.600 ;
        RECT 266.935 52.790 267.290 53.010 ;
        RECT 267.460 52.790 267.810 53.410 ;
        RECT 267.980 52.500 268.150 53.860 ;
        RECT 268.515 53.690 268.840 54.475 ;
        RECT 268.320 52.640 268.780 53.690 ;
        RECT 266.595 52.330 267.450 52.500 ;
        RECT 267.655 52.330 268.150 52.500 ;
        RECT 268.320 52.110 268.650 52.470 ;
        RECT 269.010 52.370 269.180 54.490 ;
        RECT 269.350 54.160 269.680 54.660 ;
        RECT 269.850 53.990 270.105 54.490 ;
        RECT 269.355 53.820 270.105 53.990 ;
        RECT 269.355 52.830 269.585 53.820 ;
        RECT 269.755 53.000 270.105 53.650 ;
        RECT 270.280 53.520 270.665 54.490 ;
        RECT 270.835 54.200 271.160 54.660 ;
        RECT 271.680 54.030 271.960 54.490 ;
        RECT 270.835 53.810 271.960 54.030 ;
        RECT 270.280 52.850 270.560 53.520 ;
        RECT 270.835 53.350 271.285 53.810 ;
        RECT 272.150 53.640 272.550 54.490 ;
        RECT 272.950 54.200 273.220 54.660 ;
        RECT 273.390 54.030 273.675 54.490 ;
        RECT 270.730 53.020 271.285 53.350 ;
        RECT 271.455 53.080 272.550 53.640 ;
        RECT 270.835 52.910 271.285 53.020 ;
        RECT 269.355 52.660 270.105 52.830 ;
        RECT 269.350 52.110 269.680 52.490 ;
        RECT 269.850 52.370 270.105 52.660 ;
        RECT 270.280 52.280 270.665 52.850 ;
        RECT 270.835 52.740 271.960 52.910 ;
        RECT 270.835 52.110 271.160 52.570 ;
        RECT 271.680 52.280 271.960 52.740 ;
        RECT 272.150 52.280 272.550 53.080 ;
        RECT 272.720 53.810 273.675 54.030 ;
        RECT 272.720 52.910 272.930 53.810 ;
        RECT 273.100 53.080 273.790 53.640 ;
        RECT 273.960 53.570 277.470 54.660 ;
        RECT 272.720 52.740 273.675 52.910 ;
        RECT 272.950 52.110 273.220 52.570 ;
        RECT 273.390 52.280 273.675 52.740 ;
        RECT 273.960 52.880 275.610 53.400 ;
        RECT 275.780 53.050 277.470 53.570 ;
        RECT 278.100 53.495 278.390 54.660 ;
        RECT 278.560 53.570 281.150 54.660 ;
        RECT 278.560 52.880 279.770 53.400 ;
        RECT 279.940 53.050 281.150 53.570 ;
        RECT 281.325 53.520 281.660 54.490 ;
        RECT 281.830 53.520 282.000 54.660 ;
        RECT 282.170 54.320 284.200 54.490 ;
        RECT 273.960 52.110 277.470 52.880 ;
        RECT 278.100 52.110 278.390 52.835 ;
        RECT 278.560 52.110 281.150 52.880 ;
        RECT 281.325 52.850 281.495 53.520 ;
        RECT 282.170 53.350 282.340 54.320 ;
        RECT 281.665 53.020 281.920 53.350 ;
        RECT 282.145 53.020 282.340 53.350 ;
        RECT 282.510 53.980 283.635 54.150 ;
        RECT 281.750 52.850 281.920 53.020 ;
        RECT 282.510 52.850 282.680 53.980 ;
        RECT 281.325 52.280 281.580 52.850 ;
        RECT 281.750 52.680 282.680 52.850 ;
        RECT 282.850 53.640 283.860 53.810 ;
        RECT 282.850 52.840 283.020 53.640 ;
        RECT 282.505 52.645 282.680 52.680 ;
        RECT 281.750 52.110 282.080 52.510 ;
        RECT 282.505 52.280 283.035 52.645 ;
        RECT 283.225 52.620 283.500 53.440 ;
        RECT 283.220 52.450 283.500 52.620 ;
        RECT 283.225 52.280 283.500 52.450 ;
        RECT 283.670 52.280 283.860 53.640 ;
        RECT 284.030 53.655 284.200 54.320 ;
        RECT 284.370 53.900 284.540 54.660 ;
        RECT 284.775 53.900 285.290 54.310 ;
        RECT 284.030 53.465 284.780 53.655 ;
        RECT 284.950 53.090 285.290 53.900 ;
        RECT 285.470 53.640 285.800 54.490 ;
        RECT 285.970 53.810 286.140 54.660 ;
        RECT 286.310 53.640 286.640 54.490 ;
        RECT 286.810 53.810 286.980 54.660 ;
        RECT 287.150 53.640 287.480 54.490 ;
        RECT 287.650 53.860 287.820 54.660 ;
        RECT 287.990 53.640 288.320 54.490 ;
        RECT 288.490 53.860 288.660 54.660 ;
        RECT 288.830 53.640 289.160 54.490 ;
        RECT 289.330 53.860 289.500 54.660 ;
        RECT 289.670 53.640 290.000 54.490 ;
        RECT 290.170 53.860 290.340 54.660 ;
        RECT 290.510 53.640 290.840 54.490 ;
        RECT 291.010 53.860 291.180 54.660 ;
        RECT 291.350 53.640 291.680 54.490 ;
        RECT 291.850 53.860 292.020 54.660 ;
        RECT 292.190 53.640 292.520 54.490 ;
        RECT 292.690 53.860 292.860 54.660 ;
        RECT 293.030 53.640 293.360 54.490 ;
        RECT 293.530 53.860 293.700 54.660 ;
        RECT 293.870 53.640 294.200 54.490 ;
        RECT 294.370 53.860 294.540 54.660 ;
        RECT 294.710 53.640 295.040 54.490 ;
        RECT 295.210 53.860 295.380 54.660 ;
        RECT 295.550 53.640 295.880 54.490 ;
        RECT 296.050 53.860 296.220 54.660 ;
        RECT 285.470 53.470 286.980 53.640 ;
        RECT 287.150 53.470 289.500 53.640 ;
        RECT 289.670 53.470 296.330 53.640 ;
        RECT 296.500 53.570 300.010 54.660 ;
        RECT 286.810 53.300 286.980 53.470 ;
        RECT 289.325 53.300 289.500 53.470 ;
        RECT 285.465 53.100 286.640 53.300 ;
        RECT 286.810 53.100 289.120 53.300 ;
        RECT 289.325 53.100 295.885 53.300 ;
        RECT 284.060 52.920 285.290 53.090 ;
        RECT 286.810 52.930 286.980 53.100 ;
        RECT 289.325 52.930 289.500 53.100 ;
        RECT 296.055 52.930 296.330 53.470 ;
        RECT 284.040 52.110 284.550 52.645 ;
        RECT 284.770 52.315 285.015 52.920 ;
        RECT 285.470 52.760 286.980 52.930 ;
        RECT 287.150 52.760 289.500 52.930 ;
        RECT 289.670 52.760 296.330 52.930 ;
        RECT 296.500 52.880 298.150 53.400 ;
        RECT 298.320 53.050 300.010 53.570 ;
        RECT 301.100 53.690 301.410 54.490 ;
        RECT 301.580 53.860 301.890 54.660 ;
        RECT 302.060 54.030 302.320 54.490 ;
        RECT 302.490 54.200 302.745 54.660 ;
        RECT 302.920 54.030 303.180 54.490 ;
        RECT 302.060 53.860 303.180 54.030 ;
        RECT 301.100 53.520 302.130 53.690 ;
        RECT 285.470 52.285 285.800 52.760 ;
        RECT 285.970 52.110 286.140 52.590 ;
        RECT 286.310 52.285 286.640 52.760 ;
        RECT 286.810 52.110 286.980 52.590 ;
        RECT 287.150 52.285 287.480 52.760 ;
        RECT 287.650 52.110 287.820 52.590 ;
        RECT 287.990 52.285 288.320 52.760 ;
        RECT 288.490 52.110 288.660 52.590 ;
        RECT 288.830 52.285 289.160 52.760 ;
        RECT 289.330 52.110 289.500 52.590 ;
        RECT 289.670 52.285 290.000 52.760 ;
        RECT 289.670 52.280 289.920 52.285 ;
        RECT 290.170 52.110 290.340 52.590 ;
        RECT 290.510 52.285 290.840 52.760 ;
        RECT 290.590 52.280 290.760 52.285 ;
        RECT 291.010 52.110 291.180 52.590 ;
        RECT 291.350 52.285 291.680 52.760 ;
        RECT 291.430 52.280 291.600 52.285 ;
        RECT 291.850 52.110 292.020 52.590 ;
        RECT 292.190 52.285 292.520 52.760 ;
        RECT 292.690 52.110 292.860 52.590 ;
        RECT 293.030 52.285 293.360 52.760 ;
        RECT 293.530 52.110 293.700 52.590 ;
        RECT 293.870 52.285 294.200 52.760 ;
        RECT 294.370 52.110 294.540 52.590 ;
        RECT 294.710 52.285 295.040 52.760 ;
        RECT 295.210 52.110 295.380 52.590 ;
        RECT 295.550 52.285 295.880 52.760 ;
        RECT 296.050 52.110 296.220 52.590 ;
        RECT 296.500 52.110 300.010 52.880 ;
        RECT 301.100 52.610 301.270 53.520 ;
        RECT 301.440 52.780 301.790 53.350 ;
        RECT 301.960 53.270 302.130 53.520 ;
        RECT 302.920 53.610 303.180 53.860 ;
        RECT 303.350 53.790 303.635 54.660 ;
        RECT 302.920 53.440 303.675 53.610 ;
        RECT 303.860 53.495 304.150 54.660 ;
        RECT 304.780 53.585 305.050 54.490 ;
        RECT 305.220 53.900 305.550 54.660 ;
        RECT 305.730 53.730 305.900 54.490 ;
        RECT 301.960 53.100 303.100 53.270 ;
        RECT 303.270 52.930 303.675 53.440 ;
        RECT 302.025 52.760 303.675 52.930 ;
        RECT 301.100 52.280 301.400 52.610 ;
        RECT 301.570 52.110 301.845 52.590 ;
        RECT 302.025 52.370 302.320 52.760 ;
        RECT 302.490 52.110 302.745 52.590 ;
        RECT 302.920 52.370 303.180 52.760 ;
        RECT 303.350 52.110 303.630 52.590 ;
        RECT 303.860 52.110 304.150 52.835 ;
        RECT 304.780 52.785 304.950 53.585 ;
        RECT 305.235 53.560 305.900 53.730 ;
        RECT 305.235 53.415 305.405 53.560 ;
        RECT 305.120 53.085 305.405 53.415 ;
        RECT 306.160 53.520 306.545 54.490 ;
        RECT 306.715 54.200 307.040 54.660 ;
        RECT 307.560 54.030 307.840 54.490 ;
        RECT 306.715 53.810 307.840 54.030 ;
        RECT 305.235 52.830 305.405 53.085 ;
        RECT 305.640 53.010 305.970 53.380 ;
        RECT 306.160 52.850 306.440 53.520 ;
        RECT 306.715 53.350 307.165 53.810 ;
        RECT 308.030 53.640 308.430 54.490 ;
        RECT 308.830 54.200 309.100 54.660 ;
        RECT 309.270 54.030 309.555 54.490 ;
        RECT 306.610 53.020 307.165 53.350 ;
        RECT 307.335 53.080 308.430 53.640 ;
        RECT 306.715 52.910 307.165 53.020 ;
        RECT 304.780 52.280 305.040 52.785 ;
        RECT 305.235 52.660 305.900 52.830 ;
        RECT 305.220 52.110 305.550 52.490 ;
        RECT 305.730 52.280 305.900 52.660 ;
        RECT 306.160 52.280 306.545 52.850 ;
        RECT 306.715 52.740 307.840 52.910 ;
        RECT 306.715 52.110 307.040 52.570 ;
        RECT 307.560 52.280 307.840 52.740 ;
        RECT 308.030 52.280 308.430 53.080 ;
        RECT 308.600 53.810 309.555 54.030 ;
        RECT 308.600 52.910 308.810 53.810 ;
        RECT 308.980 53.080 309.670 53.640 ;
        RECT 309.840 53.570 311.050 54.660 ;
        RECT 309.840 53.030 310.360 53.570 ;
        RECT 308.600 52.740 309.555 52.910 ;
        RECT 310.530 52.860 311.050 53.400 ;
        RECT 308.830 52.110 309.100 52.570 ;
        RECT 309.270 52.280 309.555 52.740 ;
        RECT 309.840 52.110 311.050 52.860 ;
        RECT 162.095 51.940 311.135 52.110 ;
        RECT 162.180 51.190 163.390 51.940 ;
        RECT 162.180 50.650 162.700 51.190 ;
        RECT 163.560 51.170 166.150 51.940 ;
        RECT 166.325 51.390 166.580 51.680 ;
        RECT 166.750 51.560 167.080 51.940 ;
        RECT 166.325 51.220 167.075 51.390 ;
        RECT 162.870 50.480 163.390 51.020 ;
        RECT 163.560 50.650 164.770 51.170 ;
        RECT 164.940 50.480 166.150 51.000 ;
        RECT 162.180 49.390 163.390 50.480 ;
        RECT 163.560 49.390 166.150 50.480 ;
        RECT 166.325 50.400 166.675 51.050 ;
        RECT 166.845 50.230 167.075 51.220 ;
        RECT 166.325 50.060 167.075 50.230 ;
        RECT 166.325 49.560 166.580 50.060 ;
        RECT 166.750 49.390 167.080 49.890 ;
        RECT 167.250 49.560 167.420 51.680 ;
        RECT 167.780 51.580 168.110 51.940 ;
        RECT 168.280 51.550 168.775 51.720 ;
        RECT 168.980 51.550 169.835 51.720 ;
        RECT 167.650 50.360 168.110 51.410 ;
        RECT 167.590 49.575 167.915 50.360 ;
        RECT 168.280 50.190 168.450 51.550 ;
        RECT 168.620 50.640 168.970 51.260 ;
        RECT 169.140 51.040 169.495 51.260 ;
        RECT 169.140 50.450 169.310 51.040 ;
        RECT 169.665 50.840 169.835 51.550 ;
        RECT 170.710 51.480 171.040 51.940 ;
        RECT 171.250 51.580 171.600 51.750 ;
        RECT 170.040 51.010 170.830 51.260 ;
        RECT 171.250 51.190 171.510 51.580 ;
        RECT 171.820 51.490 172.770 51.770 ;
        RECT 172.940 51.500 173.130 51.940 ;
        RECT 173.300 51.560 174.370 51.730 ;
        RECT 171.000 50.840 171.170 51.020 ;
        RECT 168.280 50.020 168.675 50.190 ;
        RECT 168.845 50.060 169.310 50.450 ;
        RECT 169.480 50.670 171.170 50.840 ;
        RECT 168.505 49.890 168.675 50.020 ;
        RECT 169.480 49.890 169.650 50.670 ;
        RECT 171.340 50.500 171.510 51.190 ;
        RECT 170.010 50.330 171.510 50.500 ;
        RECT 171.700 50.530 171.910 51.320 ;
        RECT 172.080 50.700 172.430 51.320 ;
        RECT 172.600 50.710 172.770 51.490 ;
        RECT 173.300 51.330 173.470 51.560 ;
        RECT 172.940 51.160 173.470 51.330 ;
        RECT 172.940 50.880 173.160 51.160 ;
        RECT 173.640 50.990 173.880 51.390 ;
        RECT 172.600 50.540 173.005 50.710 ;
        RECT 173.340 50.620 173.880 50.990 ;
        RECT 174.050 51.205 174.370 51.560 ;
        RECT 174.615 51.480 174.920 51.940 ;
        RECT 175.090 51.230 175.345 51.760 ;
        RECT 174.050 51.030 174.375 51.205 ;
        RECT 174.050 50.730 174.965 51.030 ;
        RECT 174.225 50.700 174.965 50.730 ;
        RECT 171.700 50.370 172.375 50.530 ;
        RECT 172.835 50.450 173.005 50.540 ;
        RECT 171.700 50.360 172.665 50.370 ;
        RECT 171.340 50.190 171.510 50.330 ;
        RECT 168.085 49.390 168.335 49.850 ;
        RECT 168.505 49.560 168.755 49.890 ;
        RECT 168.970 49.560 169.650 49.890 ;
        RECT 169.820 49.990 170.895 50.160 ;
        RECT 171.340 50.020 171.900 50.190 ;
        RECT 172.205 50.070 172.665 50.360 ;
        RECT 172.835 50.280 174.055 50.450 ;
        RECT 169.820 49.650 169.990 49.990 ;
        RECT 170.225 49.390 170.555 49.820 ;
        RECT 170.725 49.650 170.895 49.990 ;
        RECT 171.190 49.390 171.560 49.850 ;
        RECT 171.730 49.560 171.900 50.020 ;
        RECT 172.835 49.900 173.005 50.280 ;
        RECT 174.225 50.110 174.395 50.700 ;
        RECT 175.135 50.580 175.345 51.230 ;
        RECT 172.135 49.560 173.005 49.900 ;
        RECT 173.595 49.940 174.395 50.110 ;
        RECT 173.175 49.390 173.425 49.850 ;
        RECT 173.595 49.650 173.765 49.940 ;
        RECT 173.945 49.390 174.275 49.770 ;
        RECT 174.615 49.390 174.920 50.530 ;
        RECT 175.090 49.700 175.345 50.580 ;
        RECT 175.520 51.440 175.820 51.770 ;
        RECT 175.990 51.460 176.265 51.940 ;
        RECT 175.520 50.530 175.690 51.440 ;
        RECT 176.445 51.290 176.740 51.680 ;
        RECT 176.910 51.460 177.165 51.940 ;
        RECT 177.340 51.290 177.600 51.680 ;
        RECT 177.770 51.460 178.050 51.940 ;
        RECT 175.860 50.700 176.210 51.270 ;
        RECT 176.445 51.120 178.095 51.290 ;
        RECT 176.380 50.780 177.520 50.950 ;
        RECT 176.380 50.530 176.550 50.780 ;
        RECT 177.690 50.610 178.095 51.120 ;
        RECT 178.280 51.170 181.790 51.940 ;
        RECT 178.280 50.650 179.930 51.170 ;
        RECT 182.890 51.130 183.160 51.940 ;
        RECT 183.330 51.130 183.660 51.770 ;
        RECT 183.830 51.130 184.070 51.940 ;
        RECT 184.265 51.685 184.600 51.730 ;
        RECT 184.260 51.220 184.600 51.685 ;
        RECT 184.770 51.560 185.100 51.940 ;
        RECT 175.520 50.360 176.550 50.530 ;
        RECT 177.340 50.440 178.095 50.610 ;
        RECT 180.100 50.480 181.790 51.000 ;
        RECT 182.880 50.700 183.230 50.950 ;
        RECT 183.400 50.530 183.570 51.130 ;
        RECT 183.740 50.700 184.090 50.950 ;
        RECT 184.260 50.530 184.430 51.220 ;
        RECT 184.600 50.700 184.860 51.030 ;
        RECT 175.520 49.560 175.830 50.360 ;
        RECT 177.340 50.190 177.600 50.440 ;
        RECT 176.000 49.390 176.310 50.190 ;
        RECT 176.480 50.020 177.600 50.190 ;
        RECT 176.480 49.560 176.740 50.020 ;
        RECT 176.910 49.390 177.165 49.850 ;
        RECT 177.340 49.560 177.600 50.020 ;
        RECT 177.770 49.390 178.055 50.260 ;
        RECT 178.280 49.390 181.790 50.480 ;
        RECT 182.890 49.390 183.220 50.530 ;
        RECT 183.400 50.360 184.080 50.530 ;
        RECT 183.750 49.575 184.080 50.360 ;
        RECT 184.260 49.560 184.520 50.530 ;
        RECT 184.690 50.150 184.860 50.700 ;
        RECT 185.030 50.330 185.370 51.360 ;
        RECT 185.560 50.580 185.830 51.605 ;
        RECT 185.560 50.410 185.870 50.580 ;
        RECT 185.560 50.330 185.830 50.410 ;
        RECT 186.055 50.330 186.335 51.605 ;
        RECT 186.535 51.440 186.765 51.770 ;
        RECT 187.010 51.560 187.340 51.940 ;
        RECT 186.535 50.150 186.705 51.440 ;
        RECT 187.510 51.370 187.685 51.770 ;
        RECT 187.055 51.200 187.685 51.370 ;
        RECT 187.940 51.215 188.230 51.940 ;
        RECT 187.055 51.030 187.225 51.200 ;
        RECT 188.440 51.120 188.670 51.940 ;
        RECT 188.840 51.140 189.170 51.770 ;
        RECT 186.875 50.700 187.225 51.030 ;
        RECT 184.690 49.980 186.705 50.150 ;
        RECT 187.055 50.180 187.225 50.700 ;
        RECT 187.405 50.350 187.770 51.030 ;
        RECT 188.420 50.700 188.750 50.950 ;
        RECT 187.055 50.010 187.685 50.180 ;
        RECT 184.715 49.390 185.045 49.800 ;
        RECT 185.245 49.560 185.415 49.980 ;
        RECT 185.630 49.390 186.300 49.800 ;
        RECT 186.535 49.560 186.705 49.980 ;
        RECT 187.010 49.390 187.340 49.830 ;
        RECT 187.510 49.560 187.685 50.010 ;
        RECT 187.940 49.390 188.230 50.555 ;
        RECT 188.920 50.540 189.170 51.140 ;
        RECT 189.340 51.120 189.550 51.940 ;
        RECT 190.300 51.480 190.545 51.940 ;
        RECT 190.240 50.700 190.555 51.310 ;
        RECT 190.725 50.950 190.975 51.760 ;
        RECT 191.145 51.415 191.405 51.940 ;
        RECT 191.575 51.290 191.835 51.745 ;
        RECT 192.005 51.460 192.265 51.940 ;
        RECT 192.435 51.290 192.695 51.745 ;
        RECT 192.865 51.460 193.125 51.940 ;
        RECT 193.295 51.290 193.555 51.745 ;
        RECT 193.725 51.460 193.985 51.940 ;
        RECT 194.155 51.290 194.415 51.745 ;
        RECT 194.585 51.460 194.885 51.940 ;
        RECT 195.305 51.390 195.560 51.680 ;
        RECT 195.730 51.560 196.060 51.940 ;
        RECT 191.575 51.120 194.885 51.290 ;
        RECT 195.305 51.220 196.055 51.390 ;
        RECT 190.725 50.700 193.745 50.950 ;
        RECT 188.440 49.390 188.670 50.530 ;
        RECT 188.840 49.560 189.170 50.540 ;
        RECT 189.340 49.390 189.550 50.530 ;
        RECT 190.250 49.390 190.545 50.500 ;
        RECT 190.725 49.565 190.975 50.700 ;
        RECT 193.915 50.530 194.885 51.120 ;
        RECT 191.145 49.390 191.405 50.500 ;
        RECT 191.575 50.290 194.885 50.530 ;
        RECT 195.305 50.400 195.655 51.050 ;
        RECT 191.575 49.565 191.835 50.290 ;
        RECT 192.005 49.390 192.265 50.120 ;
        RECT 192.435 49.565 192.695 50.290 ;
        RECT 192.865 49.390 193.125 50.120 ;
        RECT 193.295 49.565 193.555 50.290 ;
        RECT 193.725 49.390 193.985 50.120 ;
        RECT 194.155 49.565 194.415 50.290 ;
        RECT 195.825 50.230 196.055 51.220 ;
        RECT 194.585 49.390 194.880 50.120 ;
        RECT 195.305 50.060 196.055 50.230 ;
        RECT 195.305 49.560 195.560 50.060 ;
        RECT 195.730 49.390 196.060 49.890 ;
        RECT 196.230 49.560 196.400 51.680 ;
        RECT 196.760 51.580 197.090 51.940 ;
        RECT 197.260 51.550 197.755 51.720 ;
        RECT 197.960 51.550 198.815 51.720 ;
        RECT 196.630 50.360 197.090 51.410 ;
        RECT 196.570 49.575 196.895 50.360 ;
        RECT 197.260 50.190 197.430 51.550 ;
        RECT 197.600 50.640 197.950 51.260 ;
        RECT 198.120 51.040 198.475 51.260 ;
        RECT 198.120 50.450 198.290 51.040 ;
        RECT 198.645 50.840 198.815 51.550 ;
        RECT 199.690 51.480 200.020 51.940 ;
        RECT 200.230 51.580 200.580 51.750 ;
        RECT 199.020 51.010 199.810 51.260 ;
        RECT 200.230 51.190 200.490 51.580 ;
        RECT 200.800 51.490 201.750 51.770 ;
        RECT 201.920 51.500 202.110 51.940 ;
        RECT 202.280 51.560 203.350 51.730 ;
        RECT 199.980 50.840 200.150 51.020 ;
        RECT 197.260 50.020 197.655 50.190 ;
        RECT 197.825 50.060 198.290 50.450 ;
        RECT 198.460 50.670 200.150 50.840 ;
        RECT 197.485 49.890 197.655 50.020 ;
        RECT 198.460 49.890 198.630 50.670 ;
        RECT 200.320 50.500 200.490 51.190 ;
        RECT 198.990 50.330 200.490 50.500 ;
        RECT 200.680 50.530 200.890 51.320 ;
        RECT 201.060 50.700 201.410 51.320 ;
        RECT 201.580 50.710 201.750 51.490 ;
        RECT 202.280 51.330 202.450 51.560 ;
        RECT 201.920 51.160 202.450 51.330 ;
        RECT 201.920 50.880 202.140 51.160 ;
        RECT 202.620 50.990 202.860 51.390 ;
        RECT 201.580 50.540 201.985 50.710 ;
        RECT 202.320 50.620 202.860 50.990 ;
        RECT 203.030 51.205 203.350 51.560 ;
        RECT 203.595 51.480 203.900 51.940 ;
        RECT 204.070 51.230 204.325 51.760 ;
        RECT 203.030 51.030 203.355 51.205 ;
        RECT 203.030 50.730 203.945 51.030 ;
        RECT 203.205 50.700 203.945 50.730 ;
        RECT 200.680 50.370 201.355 50.530 ;
        RECT 201.815 50.450 201.985 50.540 ;
        RECT 200.680 50.360 201.645 50.370 ;
        RECT 200.320 50.190 200.490 50.330 ;
        RECT 197.065 49.390 197.315 49.850 ;
        RECT 197.485 49.560 197.735 49.890 ;
        RECT 197.950 49.560 198.630 49.890 ;
        RECT 198.800 49.990 199.875 50.160 ;
        RECT 200.320 50.020 200.880 50.190 ;
        RECT 201.185 50.070 201.645 50.360 ;
        RECT 201.815 50.280 203.035 50.450 ;
        RECT 198.800 49.650 198.970 49.990 ;
        RECT 199.205 49.390 199.535 49.820 ;
        RECT 199.705 49.650 199.875 49.990 ;
        RECT 200.170 49.390 200.540 49.850 ;
        RECT 200.710 49.560 200.880 50.020 ;
        RECT 201.815 49.900 201.985 50.280 ;
        RECT 203.205 50.110 203.375 50.700 ;
        RECT 204.115 50.580 204.325 51.230 ;
        RECT 204.505 51.390 204.760 51.680 ;
        RECT 204.930 51.560 205.260 51.940 ;
        RECT 204.505 51.220 205.255 51.390 ;
        RECT 201.115 49.560 201.985 49.900 ;
        RECT 202.575 49.940 203.375 50.110 ;
        RECT 202.155 49.390 202.405 49.850 ;
        RECT 202.575 49.650 202.745 49.940 ;
        RECT 202.925 49.390 203.255 49.770 ;
        RECT 203.595 49.390 203.900 50.530 ;
        RECT 204.070 49.700 204.325 50.580 ;
        RECT 204.505 50.400 204.855 51.050 ;
        RECT 205.025 50.230 205.255 51.220 ;
        RECT 204.505 50.060 205.255 50.230 ;
        RECT 204.505 49.560 204.760 50.060 ;
        RECT 204.930 49.390 205.260 49.890 ;
        RECT 205.430 49.560 205.600 51.680 ;
        RECT 205.960 51.580 206.290 51.940 ;
        RECT 206.460 51.550 206.955 51.720 ;
        RECT 207.160 51.550 208.015 51.720 ;
        RECT 205.830 50.360 206.290 51.410 ;
        RECT 205.770 49.575 206.095 50.360 ;
        RECT 206.460 50.190 206.630 51.550 ;
        RECT 206.800 50.640 207.150 51.260 ;
        RECT 207.320 51.040 207.675 51.260 ;
        RECT 207.320 50.450 207.490 51.040 ;
        RECT 207.845 50.840 208.015 51.550 ;
        RECT 208.890 51.480 209.220 51.940 ;
        RECT 209.430 51.580 209.780 51.750 ;
        RECT 208.220 51.010 209.010 51.260 ;
        RECT 209.430 51.190 209.690 51.580 ;
        RECT 210.000 51.490 210.950 51.770 ;
        RECT 211.120 51.500 211.310 51.940 ;
        RECT 211.480 51.560 212.550 51.730 ;
        RECT 209.180 50.840 209.350 51.020 ;
        RECT 206.460 50.020 206.855 50.190 ;
        RECT 207.025 50.060 207.490 50.450 ;
        RECT 207.660 50.670 209.350 50.840 ;
        RECT 206.685 49.890 206.855 50.020 ;
        RECT 207.660 49.890 207.830 50.670 ;
        RECT 209.520 50.500 209.690 51.190 ;
        RECT 208.190 50.330 209.690 50.500 ;
        RECT 209.880 50.530 210.090 51.320 ;
        RECT 210.260 50.700 210.610 51.320 ;
        RECT 210.780 50.710 210.950 51.490 ;
        RECT 211.480 51.330 211.650 51.560 ;
        RECT 211.120 51.160 211.650 51.330 ;
        RECT 211.120 50.880 211.340 51.160 ;
        RECT 211.820 50.990 212.060 51.390 ;
        RECT 210.780 50.540 211.185 50.710 ;
        RECT 211.520 50.620 212.060 50.990 ;
        RECT 212.230 51.205 212.550 51.560 ;
        RECT 212.795 51.480 213.100 51.940 ;
        RECT 213.270 51.230 213.525 51.760 ;
        RECT 212.230 51.030 212.555 51.205 ;
        RECT 212.230 50.730 213.145 51.030 ;
        RECT 212.405 50.700 213.145 50.730 ;
        RECT 209.880 50.370 210.555 50.530 ;
        RECT 211.015 50.450 211.185 50.540 ;
        RECT 209.880 50.360 210.845 50.370 ;
        RECT 209.520 50.190 209.690 50.330 ;
        RECT 206.265 49.390 206.515 49.850 ;
        RECT 206.685 49.560 206.935 49.890 ;
        RECT 207.150 49.560 207.830 49.890 ;
        RECT 208.000 49.990 209.075 50.160 ;
        RECT 209.520 50.020 210.080 50.190 ;
        RECT 210.385 50.070 210.845 50.360 ;
        RECT 211.015 50.280 212.235 50.450 ;
        RECT 208.000 49.650 208.170 49.990 ;
        RECT 208.405 49.390 208.735 49.820 ;
        RECT 208.905 49.650 209.075 49.990 ;
        RECT 209.370 49.390 209.740 49.850 ;
        RECT 209.910 49.560 210.080 50.020 ;
        RECT 211.015 49.900 211.185 50.280 ;
        RECT 212.405 50.110 212.575 50.700 ;
        RECT 213.315 50.580 213.525 51.230 ;
        RECT 213.700 51.215 213.990 51.940 ;
        RECT 214.160 51.170 217.670 51.940 ;
        RECT 217.900 51.480 218.145 51.940 ;
        RECT 214.160 50.650 215.810 51.170 ;
        RECT 210.315 49.560 211.185 49.900 ;
        RECT 211.775 49.940 212.575 50.110 ;
        RECT 211.355 49.390 211.605 49.850 ;
        RECT 211.775 49.650 211.945 49.940 ;
        RECT 212.125 49.390 212.455 49.770 ;
        RECT 212.795 49.390 213.100 50.530 ;
        RECT 213.270 49.700 213.525 50.580 ;
        RECT 213.700 49.390 213.990 50.555 ;
        RECT 215.980 50.480 217.670 51.000 ;
        RECT 217.840 50.700 218.155 51.310 ;
        RECT 218.325 50.950 218.575 51.760 ;
        RECT 218.745 51.415 219.005 51.940 ;
        RECT 219.175 51.290 219.435 51.745 ;
        RECT 219.605 51.460 219.865 51.940 ;
        RECT 220.035 51.290 220.295 51.745 ;
        RECT 220.465 51.460 220.725 51.940 ;
        RECT 220.895 51.290 221.155 51.745 ;
        RECT 221.325 51.460 221.585 51.940 ;
        RECT 221.755 51.290 222.015 51.745 ;
        RECT 222.185 51.460 222.485 51.940 ;
        RECT 222.910 51.290 223.240 51.765 ;
        RECT 223.410 51.460 223.580 51.940 ;
        RECT 223.750 51.290 224.080 51.765 ;
        RECT 224.250 51.460 224.420 51.940 ;
        RECT 224.590 51.290 224.920 51.765 ;
        RECT 225.090 51.460 225.260 51.940 ;
        RECT 225.430 51.290 225.760 51.765 ;
        RECT 225.930 51.460 226.100 51.940 ;
        RECT 226.270 51.290 226.600 51.765 ;
        RECT 226.770 51.460 226.940 51.940 ;
        RECT 227.110 51.765 227.360 51.770 ;
        RECT 227.110 51.290 227.440 51.765 ;
        RECT 227.610 51.460 227.780 51.940 ;
        RECT 228.030 51.765 228.200 51.770 ;
        RECT 227.950 51.290 228.280 51.765 ;
        RECT 228.450 51.460 228.620 51.940 ;
        RECT 228.870 51.765 229.040 51.770 ;
        RECT 228.790 51.290 229.120 51.765 ;
        RECT 229.290 51.460 229.460 51.940 ;
        RECT 229.630 51.290 229.960 51.765 ;
        RECT 230.130 51.460 230.300 51.940 ;
        RECT 230.470 51.290 230.800 51.765 ;
        RECT 230.970 51.460 231.140 51.940 ;
        RECT 231.310 51.290 231.640 51.765 ;
        RECT 231.810 51.460 231.980 51.940 ;
        RECT 232.150 51.290 232.480 51.765 ;
        RECT 232.650 51.460 232.820 51.940 ;
        RECT 232.990 51.290 233.320 51.765 ;
        RECT 233.490 51.460 233.660 51.940 ;
        RECT 219.175 51.120 222.485 51.290 ;
        RECT 222.910 51.120 224.420 51.290 ;
        RECT 224.590 51.120 226.940 51.290 ;
        RECT 227.110 51.120 233.770 51.290 ;
        RECT 218.325 50.700 221.345 50.950 ;
        RECT 214.160 49.390 217.670 50.480 ;
        RECT 217.850 49.390 218.145 50.500 ;
        RECT 218.325 49.565 218.575 50.700 ;
        RECT 221.515 50.530 222.485 51.120 ;
        RECT 224.250 50.950 224.420 51.120 ;
        RECT 226.765 50.950 226.940 51.120 ;
        RECT 222.905 50.750 224.080 50.950 ;
        RECT 224.250 50.750 226.560 50.950 ;
        RECT 226.765 50.750 233.325 50.950 ;
        RECT 224.250 50.580 224.420 50.750 ;
        RECT 226.765 50.580 226.940 50.750 ;
        RECT 233.495 50.580 233.770 51.120 ;
        RECT 233.940 51.170 235.610 51.940 ;
        RECT 235.780 51.200 236.165 51.770 ;
        RECT 236.335 51.480 236.660 51.940 ;
        RECT 237.180 51.310 237.460 51.770 ;
        RECT 233.940 50.650 234.690 51.170 ;
        RECT 218.745 49.390 219.005 50.500 ;
        RECT 219.175 50.290 222.485 50.530 ;
        RECT 222.910 50.410 224.420 50.580 ;
        RECT 224.590 50.410 226.940 50.580 ;
        RECT 227.110 50.410 233.770 50.580 ;
        RECT 234.860 50.480 235.610 51.000 ;
        RECT 219.175 49.565 219.435 50.290 ;
        RECT 219.605 49.390 219.865 50.120 ;
        RECT 220.035 49.565 220.295 50.290 ;
        RECT 220.465 49.390 220.725 50.120 ;
        RECT 220.895 49.565 221.155 50.290 ;
        RECT 221.325 49.390 221.585 50.120 ;
        RECT 221.755 49.565 222.015 50.290 ;
        RECT 222.185 49.390 222.480 50.120 ;
        RECT 222.910 49.560 223.240 50.410 ;
        RECT 223.410 49.390 223.580 50.240 ;
        RECT 223.750 49.560 224.080 50.410 ;
        RECT 224.250 49.390 224.420 50.240 ;
        RECT 224.590 49.560 224.920 50.410 ;
        RECT 225.090 49.390 225.260 50.190 ;
        RECT 225.430 49.560 225.760 50.410 ;
        RECT 225.930 49.390 226.100 50.190 ;
        RECT 226.270 49.560 226.600 50.410 ;
        RECT 226.770 49.390 226.940 50.190 ;
        RECT 227.110 49.560 227.440 50.410 ;
        RECT 227.610 49.390 227.780 50.190 ;
        RECT 227.950 49.560 228.280 50.410 ;
        RECT 228.450 49.390 228.620 50.190 ;
        RECT 228.790 49.560 229.120 50.410 ;
        RECT 229.290 49.390 229.460 50.190 ;
        RECT 229.630 49.560 229.960 50.410 ;
        RECT 230.130 49.390 230.300 50.190 ;
        RECT 230.470 49.560 230.800 50.410 ;
        RECT 230.970 49.390 231.140 50.190 ;
        RECT 231.310 49.560 231.640 50.410 ;
        RECT 231.810 49.390 231.980 50.190 ;
        RECT 232.150 49.560 232.480 50.410 ;
        RECT 232.650 49.390 232.820 50.190 ;
        RECT 232.990 49.560 233.320 50.410 ;
        RECT 233.490 49.390 233.660 50.190 ;
        RECT 233.940 49.390 235.610 50.480 ;
        RECT 235.780 50.530 236.060 51.200 ;
        RECT 236.335 51.140 237.460 51.310 ;
        RECT 236.335 51.030 236.785 51.140 ;
        RECT 236.230 50.700 236.785 51.030 ;
        RECT 237.650 50.970 238.050 51.770 ;
        RECT 238.450 51.480 238.720 51.940 ;
        RECT 238.890 51.310 239.175 51.770 ;
        RECT 235.780 49.560 236.165 50.530 ;
        RECT 236.335 50.240 236.785 50.700 ;
        RECT 236.955 50.410 238.050 50.970 ;
        RECT 236.335 50.020 237.460 50.240 ;
        RECT 236.335 49.390 236.660 49.850 ;
        RECT 237.180 49.560 237.460 50.020 ;
        RECT 237.650 49.560 238.050 50.410 ;
        RECT 238.220 51.140 239.175 51.310 ;
        RECT 239.460 51.215 239.750 51.940 ;
        RECT 239.920 51.170 241.590 51.940 ;
        RECT 241.760 51.200 242.145 51.770 ;
        RECT 242.315 51.480 242.640 51.940 ;
        RECT 243.160 51.310 243.440 51.770 ;
        RECT 238.220 50.240 238.430 51.140 ;
        RECT 238.600 50.410 239.290 50.970 ;
        RECT 239.920 50.650 240.670 51.170 ;
        RECT 238.220 50.020 239.175 50.240 ;
        RECT 238.450 49.390 238.720 49.850 ;
        RECT 238.890 49.560 239.175 50.020 ;
        RECT 239.460 49.390 239.750 50.555 ;
        RECT 240.840 50.480 241.590 51.000 ;
        RECT 239.920 49.390 241.590 50.480 ;
        RECT 241.760 50.530 242.040 51.200 ;
        RECT 242.315 51.140 243.440 51.310 ;
        RECT 242.315 51.030 242.765 51.140 ;
        RECT 242.210 50.700 242.765 51.030 ;
        RECT 243.630 50.970 244.030 51.770 ;
        RECT 244.430 51.480 244.700 51.940 ;
        RECT 244.870 51.310 245.155 51.770 ;
        RECT 241.760 49.560 242.145 50.530 ;
        RECT 242.315 50.240 242.765 50.700 ;
        RECT 242.935 50.410 244.030 50.970 ;
        RECT 242.315 50.020 243.440 50.240 ;
        RECT 242.315 49.390 242.640 49.850 ;
        RECT 243.160 49.560 243.440 50.020 ;
        RECT 243.630 49.560 244.030 50.410 ;
        RECT 244.200 51.140 245.155 51.310 ;
        RECT 245.440 51.190 246.650 51.940 ;
        RECT 244.200 50.240 244.410 51.140 ;
        RECT 244.580 50.410 245.270 50.970 ;
        RECT 245.440 50.650 245.960 51.190 ;
        RECT 246.820 51.120 247.505 51.760 ;
        RECT 247.675 51.120 247.845 51.940 ;
        RECT 248.015 51.290 248.345 51.755 ;
        RECT 248.515 51.470 248.685 51.940 ;
        RECT 248.945 51.550 250.130 51.720 ;
        RECT 250.300 51.380 250.630 51.770 ;
        RECT 249.330 51.290 249.715 51.380 ;
        RECT 248.015 51.120 249.715 51.290 ;
        RECT 250.120 51.200 250.630 51.380 ;
        RECT 246.130 50.480 246.650 51.020 ;
        RECT 244.200 50.020 245.155 50.240 ;
        RECT 244.430 49.390 244.700 49.850 ;
        RECT 244.870 49.560 245.155 50.020 ;
        RECT 245.440 49.390 246.650 50.480 ;
        RECT 246.820 50.150 247.070 51.120 ;
        RECT 247.240 50.740 247.575 50.950 ;
        RECT 247.745 50.740 248.195 50.950 ;
        RECT 248.385 50.740 248.870 50.950 ;
        RECT 247.405 50.570 247.575 50.740 ;
        RECT 248.495 50.580 248.870 50.740 ;
        RECT 249.060 50.700 249.440 50.950 ;
        RECT 249.620 50.740 249.950 50.950 ;
        RECT 247.405 50.400 248.325 50.570 ;
        RECT 246.820 49.560 247.485 50.150 ;
        RECT 247.655 49.390 247.985 50.230 ;
        RECT 248.155 50.150 248.325 50.400 ;
        RECT 248.495 50.410 248.890 50.580 ;
        RECT 248.495 50.320 248.870 50.410 ;
        RECT 249.060 50.320 249.380 50.700 ;
        RECT 250.120 50.570 250.290 51.200 ;
        RECT 251.880 51.120 252.565 51.760 ;
        RECT 252.735 51.120 252.905 51.940 ;
        RECT 253.075 51.290 253.405 51.755 ;
        RECT 253.575 51.470 253.745 51.940 ;
        RECT 254.005 51.550 255.190 51.720 ;
        RECT 255.360 51.380 255.690 51.770 ;
        RECT 256.080 51.480 256.325 51.940 ;
        RECT 254.390 51.290 254.775 51.380 ;
        RECT 253.075 51.120 254.775 51.290 ;
        RECT 255.180 51.200 255.690 51.380 ;
        RECT 250.460 50.740 250.790 51.030 ;
        RECT 249.550 50.400 250.635 50.570 ;
        RECT 249.550 50.150 249.720 50.400 ;
        RECT 248.155 49.980 249.720 50.150 ;
        RECT 248.495 49.560 249.300 49.980 ;
        RECT 249.890 49.390 250.140 50.230 ;
        RECT 250.335 49.560 250.635 50.400 ;
        RECT 251.880 50.150 252.130 51.120 ;
        RECT 252.300 50.740 252.635 50.950 ;
        RECT 252.805 50.740 253.255 50.950 ;
        RECT 253.445 50.920 253.930 50.950 ;
        RECT 253.445 50.750 253.950 50.920 ;
        RECT 253.445 50.740 253.930 50.750 ;
        RECT 252.465 50.570 252.635 50.740 ;
        RECT 252.465 50.400 253.385 50.570 ;
        RECT 251.880 49.560 252.545 50.150 ;
        RECT 252.715 49.390 253.045 50.230 ;
        RECT 253.215 50.150 253.385 50.400 ;
        RECT 253.555 50.320 253.930 50.740 ;
        RECT 254.120 50.700 254.500 50.950 ;
        RECT 254.680 50.740 255.010 50.950 ;
        RECT 254.120 50.320 254.440 50.700 ;
        RECT 255.180 50.570 255.350 51.200 ;
        RECT 255.520 50.740 255.850 51.030 ;
        RECT 256.020 50.700 256.335 51.310 ;
        RECT 256.505 50.950 256.755 51.760 ;
        RECT 256.925 51.415 257.185 51.940 ;
        RECT 257.355 51.290 257.615 51.745 ;
        RECT 257.785 51.460 258.045 51.940 ;
        RECT 258.215 51.290 258.475 51.745 ;
        RECT 258.645 51.460 258.905 51.940 ;
        RECT 259.075 51.290 259.335 51.745 ;
        RECT 259.505 51.460 259.765 51.940 ;
        RECT 259.935 51.290 260.195 51.745 ;
        RECT 260.365 51.460 260.665 51.940 ;
        RECT 257.355 51.120 260.665 51.290 ;
        RECT 256.505 50.700 259.525 50.950 ;
        RECT 254.610 50.400 255.695 50.570 ;
        RECT 254.610 50.150 254.780 50.400 ;
        RECT 253.215 49.980 254.780 50.150 ;
        RECT 253.555 49.560 254.360 49.980 ;
        RECT 254.950 49.390 255.200 50.230 ;
        RECT 255.395 49.560 255.695 50.400 ;
        RECT 256.030 49.390 256.325 50.500 ;
        RECT 256.505 49.565 256.755 50.700 ;
        RECT 259.695 50.530 260.665 51.120 ;
        RECT 256.925 49.390 257.185 50.500 ;
        RECT 257.355 50.290 260.665 50.530 ;
        RECT 261.080 51.200 261.465 51.770 ;
        RECT 261.635 51.480 261.960 51.940 ;
        RECT 262.480 51.310 262.760 51.770 ;
        RECT 261.080 50.530 261.360 51.200 ;
        RECT 261.635 51.140 262.760 51.310 ;
        RECT 261.635 51.030 262.085 51.140 ;
        RECT 261.530 50.700 262.085 51.030 ;
        RECT 262.950 50.970 263.350 51.770 ;
        RECT 263.750 51.480 264.020 51.940 ;
        RECT 264.190 51.310 264.475 51.770 ;
        RECT 257.355 49.565 257.615 50.290 ;
        RECT 257.785 49.390 258.045 50.120 ;
        RECT 258.215 49.565 258.475 50.290 ;
        RECT 258.645 49.390 258.905 50.120 ;
        RECT 259.075 49.565 259.335 50.290 ;
        RECT 259.505 49.390 259.765 50.120 ;
        RECT 259.935 49.565 260.195 50.290 ;
        RECT 260.365 49.390 260.660 50.120 ;
        RECT 261.080 49.560 261.465 50.530 ;
        RECT 261.635 50.240 262.085 50.700 ;
        RECT 262.255 50.410 263.350 50.970 ;
        RECT 261.635 50.020 262.760 50.240 ;
        RECT 261.635 49.390 261.960 49.850 ;
        RECT 262.480 49.560 262.760 50.020 ;
        RECT 262.950 49.560 263.350 50.410 ;
        RECT 263.520 51.140 264.475 51.310 ;
        RECT 265.220 51.215 265.510 51.940 ;
        RECT 263.520 50.240 263.730 51.140 ;
        RECT 265.740 51.120 265.950 51.940 ;
        RECT 266.120 51.140 266.450 51.770 ;
        RECT 263.900 50.410 264.590 50.970 ;
        RECT 263.520 50.020 264.475 50.240 ;
        RECT 263.750 49.390 264.020 49.850 ;
        RECT 264.190 49.560 264.475 50.020 ;
        RECT 265.220 49.390 265.510 50.555 ;
        RECT 266.120 50.540 266.370 51.140 ;
        RECT 266.620 51.120 266.850 51.940 ;
        RECT 267.985 51.390 268.240 51.680 ;
        RECT 268.410 51.560 268.740 51.940 ;
        RECT 267.985 51.220 268.735 51.390 ;
        RECT 266.540 50.700 266.870 50.950 ;
        RECT 265.740 49.390 265.950 50.530 ;
        RECT 266.120 49.560 266.450 50.540 ;
        RECT 266.620 49.390 266.850 50.530 ;
        RECT 267.985 50.400 268.335 51.050 ;
        RECT 268.505 50.230 268.735 51.220 ;
        RECT 267.985 50.060 268.735 50.230 ;
        RECT 267.985 49.560 268.240 50.060 ;
        RECT 268.410 49.390 268.740 49.890 ;
        RECT 268.910 49.560 269.080 51.680 ;
        RECT 269.440 51.580 269.770 51.940 ;
        RECT 269.940 51.550 270.435 51.720 ;
        RECT 270.640 51.550 271.495 51.720 ;
        RECT 269.310 50.360 269.770 51.410 ;
        RECT 269.250 49.575 269.575 50.360 ;
        RECT 269.940 50.190 270.110 51.550 ;
        RECT 270.280 50.640 270.630 51.260 ;
        RECT 270.800 51.040 271.155 51.260 ;
        RECT 270.800 50.450 270.970 51.040 ;
        RECT 271.325 50.840 271.495 51.550 ;
        RECT 272.370 51.480 272.700 51.940 ;
        RECT 272.910 51.580 273.260 51.750 ;
        RECT 271.700 51.010 272.490 51.260 ;
        RECT 272.910 51.190 273.170 51.580 ;
        RECT 273.480 51.490 274.430 51.770 ;
        RECT 274.600 51.500 274.790 51.940 ;
        RECT 274.960 51.560 276.030 51.730 ;
        RECT 272.660 50.840 272.830 51.020 ;
        RECT 269.940 50.020 270.335 50.190 ;
        RECT 270.505 50.060 270.970 50.450 ;
        RECT 271.140 50.670 272.830 50.840 ;
        RECT 270.165 49.890 270.335 50.020 ;
        RECT 271.140 49.890 271.310 50.670 ;
        RECT 273.000 50.500 273.170 51.190 ;
        RECT 271.670 50.330 273.170 50.500 ;
        RECT 273.360 50.530 273.570 51.320 ;
        RECT 273.740 50.700 274.090 51.320 ;
        RECT 274.260 50.710 274.430 51.490 ;
        RECT 274.960 51.330 275.130 51.560 ;
        RECT 274.600 51.160 275.130 51.330 ;
        RECT 274.600 50.880 274.820 51.160 ;
        RECT 275.300 50.990 275.540 51.390 ;
        RECT 274.260 50.540 274.665 50.710 ;
        RECT 275.000 50.620 275.540 50.990 ;
        RECT 275.710 51.205 276.030 51.560 ;
        RECT 276.275 51.480 276.580 51.940 ;
        RECT 276.750 51.230 277.005 51.760 ;
        RECT 275.710 51.030 276.035 51.205 ;
        RECT 275.710 50.730 276.625 51.030 ;
        RECT 275.885 50.700 276.625 50.730 ;
        RECT 273.360 50.370 274.035 50.530 ;
        RECT 274.495 50.450 274.665 50.540 ;
        RECT 273.360 50.360 274.325 50.370 ;
        RECT 273.000 50.190 273.170 50.330 ;
        RECT 269.745 49.390 269.995 49.850 ;
        RECT 270.165 49.560 270.415 49.890 ;
        RECT 270.630 49.560 271.310 49.890 ;
        RECT 271.480 49.990 272.555 50.160 ;
        RECT 273.000 50.020 273.560 50.190 ;
        RECT 273.865 50.070 274.325 50.360 ;
        RECT 274.495 50.280 275.715 50.450 ;
        RECT 271.480 49.650 271.650 49.990 ;
        RECT 271.885 49.390 272.215 49.820 ;
        RECT 272.385 49.650 272.555 49.990 ;
        RECT 272.850 49.390 273.220 49.850 ;
        RECT 273.390 49.560 273.560 50.020 ;
        RECT 274.495 49.900 274.665 50.280 ;
        RECT 275.885 50.110 276.055 50.700 ;
        RECT 276.795 50.580 277.005 51.230 ;
        RECT 277.180 51.170 278.850 51.940 ;
        RECT 279.025 51.390 279.280 51.680 ;
        RECT 279.450 51.560 279.780 51.940 ;
        RECT 279.025 51.220 279.775 51.390 ;
        RECT 277.180 50.650 277.930 51.170 ;
        RECT 273.795 49.560 274.665 49.900 ;
        RECT 275.255 49.940 276.055 50.110 ;
        RECT 274.835 49.390 275.085 49.850 ;
        RECT 275.255 49.650 275.425 49.940 ;
        RECT 275.605 49.390 275.935 49.770 ;
        RECT 276.275 49.390 276.580 50.530 ;
        RECT 276.750 49.700 277.005 50.580 ;
        RECT 278.100 50.480 278.850 51.000 ;
        RECT 277.180 49.390 278.850 50.480 ;
        RECT 279.025 50.400 279.375 51.050 ;
        RECT 279.545 50.230 279.775 51.220 ;
        RECT 279.025 50.060 279.775 50.230 ;
        RECT 279.025 49.560 279.280 50.060 ;
        RECT 279.450 49.390 279.780 49.890 ;
        RECT 279.950 49.560 280.120 51.680 ;
        RECT 280.480 51.580 280.810 51.940 ;
        RECT 280.980 51.550 281.475 51.720 ;
        RECT 281.680 51.550 282.535 51.720 ;
        RECT 280.350 50.360 280.810 51.410 ;
        RECT 280.290 49.575 280.615 50.360 ;
        RECT 280.980 50.190 281.150 51.550 ;
        RECT 281.320 50.640 281.670 51.260 ;
        RECT 281.840 51.040 282.195 51.260 ;
        RECT 281.840 50.450 282.010 51.040 ;
        RECT 282.365 50.840 282.535 51.550 ;
        RECT 283.410 51.480 283.740 51.940 ;
        RECT 283.950 51.580 284.300 51.750 ;
        RECT 282.740 51.010 283.530 51.260 ;
        RECT 283.950 51.190 284.210 51.580 ;
        RECT 284.520 51.490 285.470 51.770 ;
        RECT 285.640 51.500 285.830 51.940 ;
        RECT 286.000 51.560 287.070 51.730 ;
        RECT 283.700 50.840 283.870 51.020 ;
        RECT 280.980 50.020 281.375 50.190 ;
        RECT 281.545 50.060 282.010 50.450 ;
        RECT 282.180 50.670 283.870 50.840 ;
        RECT 281.205 49.890 281.375 50.020 ;
        RECT 282.180 49.890 282.350 50.670 ;
        RECT 284.040 50.500 284.210 51.190 ;
        RECT 282.710 50.330 284.210 50.500 ;
        RECT 284.400 50.530 284.610 51.320 ;
        RECT 284.780 50.700 285.130 51.320 ;
        RECT 285.300 50.710 285.470 51.490 ;
        RECT 286.000 51.330 286.170 51.560 ;
        RECT 285.640 51.160 286.170 51.330 ;
        RECT 285.640 50.880 285.860 51.160 ;
        RECT 286.340 50.990 286.580 51.390 ;
        RECT 285.300 50.540 285.705 50.710 ;
        RECT 286.040 50.620 286.580 50.990 ;
        RECT 286.750 51.205 287.070 51.560 ;
        RECT 287.315 51.480 287.620 51.940 ;
        RECT 287.790 51.230 288.045 51.760 ;
        RECT 288.230 51.450 288.560 51.940 ;
        RECT 288.730 51.345 289.350 51.770 ;
        RECT 286.750 51.030 287.075 51.205 ;
        RECT 286.750 50.730 287.665 51.030 ;
        RECT 286.925 50.700 287.665 50.730 ;
        RECT 284.400 50.370 285.075 50.530 ;
        RECT 285.535 50.450 285.705 50.540 ;
        RECT 284.400 50.360 285.365 50.370 ;
        RECT 284.040 50.190 284.210 50.330 ;
        RECT 280.785 49.390 281.035 49.850 ;
        RECT 281.205 49.560 281.455 49.890 ;
        RECT 281.670 49.560 282.350 49.890 ;
        RECT 282.520 49.990 283.595 50.160 ;
        RECT 284.040 50.020 284.600 50.190 ;
        RECT 284.905 50.070 285.365 50.360 ;
        RECT 285.535 50.280 286.755 50.450 ;
        RECT 282.520 49.650 282.690 49.990 ;
        RECT 282.925 49.390 283.255 49.820 ;
        RECT 283.425 49.650 283.595 49.990 ;
        RECT 283.890 49.390 284.260 49.850 ;
        RECT 284.430 49.560 284.600 50.020 ;
        RECT 285.535 49.900 285.705 50.280 ;
        RECT 286.925 50.110 287.095 50.700 ;
        RECT 287.835 50.580 288.045 51.230 ;
        RECT 288.220 50.700 288.560 51.280 ;
        RECT 288.730 51.010 289.090 51.345 ;
        RECT 289.810 51.250 290.140 51.940 ;
        RECT 290.980 51.215 291.270 51.940 ;
        RECT 291.440 51.395 296.785 51.940 ;
        RECT 288.730 50.730 290.150 51.010 ;
        RECT 284.835 49.560 285.705 49.900 ;
        RECT 286.295 49.940 287.095 50.110 ;
        RECT 285.875 49.390 286.125 49.850 ;
        RECT 286.295 49.650 286.465 49.940 ;
        RECT 286.645 49.390 286.975 49.770 ;
        RECT 287.315 49.390 287.620 50.530 ;
        RECT 287.790 49.700 288.045 50.580 ;
        RECT 288.230 49.390 288.560 50.530 ;
        RECT 288.730 49.560 289.090 50.730 ;
        RECT 289.290 49.390 289.620 50.560 ;
        RECT 289.820 49.560 290.150 50.730 ;
        RECT 293.025 50.565 293.365 51.395 ;
        RECT 296.960 51.170 299.550 51.940 ;
        RECT 299.720 51.430 299.990 51.940 ;
        RECT 300.160 51.260 300.405 51.760 ;
        RECT 299.720 51.200 300.405 51.260 ;
        RECT 300.575 51.200 300.905 51.940 ;
        RECT 299.720 51.170 300.320 51.200 ;
        RECT 290.350 49.390 290.680 50.560 ;
        RECT 290.980 49.390 291.270 50.555 ;
        RECT 294.845 49.825 295.195 51.075 ;
        RECT 296.960 50.650 298.170 51.170 ;
        RECT 299.720 51.130 300.305 51.170 ;
        RECT 298.340 50.480 299.550 51.000 ;
        RECT 291.440 49.390 296.785 49.825 ;
        RECT 296.960 49.390 299.550 50.480 ;
        RECT 299.720 50.580 300.275 51.130 ;
        RECT 301.075 51.030 301.245 51.680 ;
        RECT 300.445 50.700 301.245 51.030 ;
        RECT 299.720 50.530 300.320 50.580 ;
        RECT 299.720 50.410 300.485 50.530 ;
        RECT 299.720 49.390 299.985 50.240 ;
        RECT 300.155 49.565 300.485 50.410 ;
        RECT 300.655 49.390 300.825 50.530 ;
        RECT 300.995 50.110 301.245 50.700 ;
        RECT 301.415 51.345 301.765 51.675 ;
        RECT 301.965 51.460 302.605 51.940 ;
        RECT 302.805 51.550 303.655 51.720 ;
        RECT 301.415 50.450 301.605 51.345 ;
        RECT 301.955 51.020 302.635 51.290 ;
        RECT 302.285 50.960 302.635 51.020 ;
        RECT 301.805 50.790 302.155 50.850 ;
        RECT 302.805 50.790 302.975 51.550 ;
        RECT 304.215 51.480 304.535 51.940 ;
        RECT 304.735 51.300 304.985 51.730 ;
        RECT 305.275 51.500 305.685 51.940 ;
        RECT 305.855 51.560 306.870 51.760 ;
        RECT 303.145 51.130 304.415 51.300 ;
        RECT 303.145 51.010 303.495 51.130 ;
        RECT 301.805 50.620 303.725 50.790 ;
        RECT 301.415 50.280 303.385 50.450 ;
        RECT 301.415 50.260 301.785 50.280 ;
        RECT 300.995 49.600 301.325 50.110 ;
        RECT 301.615 49.650 301.785 50.260 ;
        RECT 303.555 50.110 303.725 50.620 ;
        RECT 303.895 50.550 304.075 50.960 ;
        RECT 304.245 50.370 304.415 51.130 ;
        RECT 301.955 49.390 302.285 50.080 ;
        RECT 302.515 49.940 303.725 50.110 ;
        RECT 303.895 50.060 304.415 50.370 ;
        RECT 304.585 50.960 304.985 51.300 ;
        RECT 305.275 50.960 305.685 51.290 ;
        RECT 304.585 50.190 304.755 50.960 ;
        RECT 305.855 50.830 306.025 51.560 ;
        RECT 307.170 51.390 307.340 51.720 ;
        RECT 307.510 51.560 307.840 51.940 ;
        RECT 308.060 51.460 308.280 51.680 ;
        RECT 308.450 51.560 308.780 51.940 ;
        RECT 306.195 51.010 306.545 51.380 ;
        RECT 305.855 50.790 306.275 50.830 ;
        RECT 304.925 50.620 306.275 50.790 ;
        RECT 304.925 50.460 305.175 50.620 ;
        RECT 305.685 50.190 305.935 50.450 ;
        RECT 304.585 49.940 305.935 50.190 ;
        RECT 302.515 49.650 302.755 49.940 ;
        RECT 303.555 49.860 303.725 49.940 ;
        RECT 302.955 49.390 303.375 49.770 ;
        RECT 303.555 49.610 304.185 49.860 ;
        RECT 304.635 49.390 304.965 49.770 ;
        RECT 305.135 49.650 305.305 49.940 ;
        RECT 306.105 49.775 306.275 50.620 ;
        RECT 306.725 50.450 306.945 51.320 ;
        RECT 307.170 51.200 307.865 51.390 ;
        RECT 306.445 50.070 306.945 50.450 ;
        RECT 307.115 50.400 307.525 51.020 ;
        RECT 307.695 50.230 307.865 51.200 ;
        RECT 307.170 50.060 307.865 50.230 ;
        RECT 305.485 49.390 305.865 49.770 ;
        RECT 306.105 49.605 306.935 49.775 ;
        RECT 307.170 49.560 307.340 50.060 ;
        RECT 308.060 49.980 308.290 51.460 ;
        RECT 308.950 51.390 309.210 51.680 ;
        RECT 308.460 51.220 309.210 51.390 ;
        RECT 308.460 50.230 308.690 51.220 ;
        RECT 309.840 51.190 311.050 51.940 ;
        RECT 308.860 50.400 309.210 51.050 ;
        RECT 309.840 50.480 310.360 51.020 ;
        RECT 310.530 50.650 311.050 51.190 ;
        RECT 308.460 50.060 309.210 50.230 ;
        RECT 307.510 49.390 307.840 49.890 ;
        RECT 308.060 49.560 308.280 49.980 ;
        RECT 308.450 49.390 308.780 49.890 ;
        RECT 308.950 49.560 309.210 50.060 ;
        RECT 309.840 49.390 311.050 50.480 ;
        RECT 162.095 49.220 311.135 49.390 ;
        RECT 162.180 48.130 163.390 49.220 ;
        RECT 163.560 48.785 168.905 49.220 ;
        RECT 162.180 47.420 162.700 47.960 ;
        RECT 162.870 47.590 163.390 48.130 ;
        RECT 162.180 46.670 163.390 47.420 ;
        RECT 165.145 47.215 165.485 48.045 ;
        RECT 166.965 47.535 167.315 48.785 ;
        RECT 169.080 48.130 170.750 49.220 ;
        RECT 169.080 47.440 169.830 47.960 ;
        RECT 170.000 47.610 170.750 48.130 ;
        RECT 170.925 48.080 171.260 49.050 ;
        RECT 171.430 48.080 171.600 49.220 ;
        RECT 171.770 48.880 173.800 49.050 ;
        RECT 163.560 46.670 168.905 47.215 ;
        RECT 169.080 46.670 170.750 47.440 ;
        RECT 170.925 47.410 171.095 48.080 ;
        RECT 171.770 47.910 171.940 48.880 ;
        RECT 171.265 47.580 171.520 47.910 ;
        RECT 171.745 47.580 171.940 47.910 ;
        RECT 172.110 48.540 173.235 48.710 ;
        RECT 171.350 47.410 171.520 47.580 ;
        RECT 172.110 47.410 172.280 48.540 ;
        RECT 170.925 46.840 171.180 47.410 ;
        RECT 171.350 47.240 172.280 47.410 ;
        RECT 172.450 48.200 173.460 48.370 ;
        RECT 172.450 47.400 172.620 48.200 ;
        RECT 172.105 47.205 172.280 47.240 ;
        RECT 171.350 46.670 171.680 47.070 ;
        RECT 172.105 46.840 172.635 47.205 ;
        RECT 172.825 47.180 173.100 48.000 ;
        RECT 172.820 47.010 173.100 47.180 ;
        RECT 172.825 46.840 173.100 47.010 ;
        RECT 173.270 46.840 173.460 48.200 ;
        RECT 173.630 48.215 173.800 48.880 ;
        RECT 173.970 48.460 174.140 49.220 ;
        RECT 174.375 48.460 174.890 48.870 ;
        RECT 173.630 48.025 174.380 48.215 ;
        RECT 174.550 47.650 174.890 48.460 ;
        RECT 175.060 48.055 175.350 49.220 ;
        RECT 175.520 48.130 176.730 49.220 ;
        RECT 173.660 47.480 174.890 47.650 ;
        RECT 173.640 46.670 174.150 47.205 ;
        RECT 174.370 46.875 174.615 47.480 ;
        RECT 175.520 47.420 176.040 47.960 ;
        RECT 176.210 47.590 176.730 48.130 ;
        RECT 176.905 48.080 177.240 49.050 ;
        RECT 177.410 48.080 177.580 49.220 ;
        RECT 177.750 48.880 179.780 49.050 ;
        RECT 175.060 46.670 175.350 47.395 ;
        RECT 175.520 46.670 176.730 47.420 ;
        RECT 176.905 47.410 177.075 48.080 ;
        RECT 177.750 47.910 177.920 48.880 ;
        RECT 177.245 47.580 177.500 47.910 ;
        RECT 177.725 47.580 177.920 47.910 ;
        RECT 178.090 48.540 179.215 48.710 ;
        RECT 177.330 47.410 177.500 47.580 ;
        RECT 178.090 47.410 178.260 48.540 ;
        RECT 176.905 46.840 177.160 47.410 ;
        RECT 177.330 47.240 178.260 47.410 ;
        RECT 178.430 48.200 179.440 48.370 ;
        RECT 178.430 47.400 178.600 48.200 ;
        RECT 178.805 47.520 179.080 48.000 ;
        RECT 178.800 47.350 179.080 47.520 ;
        RECT 178.085 47.205 178.260 47.240 ;
        RECT 177.330 46.670 177.660 47.070 ;
        RECT 178.085 46.840 178.615 47.205 ;
        RECT 178.805 46.840 179.080 47.350 ;
        RECT 179.250 46.840 179.440 48.200 ;
        RECT 179.610 48.215 179.780 48.880 ;
        RECT 179.950 48.460 180.120 49.220 ;
        RECT 180.355 48.460 180.870 48.870 ;
        RECT 179.610 48.025 180.360 48.215 ;
        RECT 180.530 47.650 180.870 48.460 ;
        RECT 181.155 48.590 181.440 49.050 ;
        RECT 181.610 48.760 181.880 49.220 ;
        RECT 181.155 48.370 182.110 48.590 ;
        RECT 179.640 47.480 180.870 47.650 ;
        RECT 181.040 47.640 181.730 48.200 ;
        RECT 179.620 46.670 180.130 47.205 ;
        RECT 180.350 46.875 180.595 47.480 ;
        RECT 181.900 47.470 182.110 48.370 ;
        RECT 181.155 47.300 182.110 47.470 ;
        RECT 182.280 48.200 182.680 49.050 ;
        RECT 182.870 48.590 183.150 49.050 ;
        RECT 183.670 48.760 183.995 49.220 ;
        RECT 182.870 48.370 183.995 48.590 ;
        RECT 182.280 47.640 183.375 48.200 ;
        RECT 183.545 47.910 183.995 48.370 ;
        RECT 184.165 48.080 184.550 49.050 ;
        RECT 184.720 48.785 190.065 49.220 ;
        RECT 181.155 46.840 181.440 47.300 ;
        RECT 181.610 46.670 181.880 47.130 ;
        RECT 182.280 46.840 182.680 47.640 ;
        RECT 183.545 47.580 184.100 47.910 ;
        RECT 183.545 47.470 183.995 47.580 ;
        RECT 182.870 47.300 183.995 47.470 ;
        RECT 184.270 47.410 184.550 48.080 ;
        RECT 182.870 46.840 183.150 47.300 ;
        RECT 183.670 46.670 183.995 47.130 ;
        RECT 184.165 46.840 184.550 47.410 ;
        RECT 186.305 47.215 186.645 48.045 ;
        RECT 188.125 47.535 188.475 48.785 ;
        RECT 190.240 48.130 192.830 49.220 ;
        RECT 190.240 47.440 191.450 47.960 ;
        RECT 191.620 47.610 192.830 48.130 ;
        RECT 193.070 48.215 193.325 49.020 ;
        RECT 193.495 48.385 193.755 49.220 ;
        RECT 193.925 48.215 194.185 49.020 ;
        RECT 194.355 48.385 194.610 49.220 ;
        RECT 195.090 48.490 195.385 49.220 ;
        RECT 195.555 48.320 195.815 49.045 ;
        RECT 195.985 48.490 196.245 49.220 ;
        RECT 196.415 48.320 196.675 49.045 ;
        RECT 196.845 48.490 197.105 49.220 ;
        RECT 197.275 48.320 197.535 49.045 ;
        RECT 197.705 48.490 197.965 49.220 ;
        RECT 198.135 48.320 198.395 49.045 ;
        RECT 193.070 48.045 194.670 48.215 ;
        RECT 193.000 47.650 194.220 47.875 ;
        RECT 194.390 47.480 194.670 48.045 ;
        RECT 184.720 46.670 190.065 47.215 ;
        RECT 190.240 46.670 192.830 47.440 ;
        RECT 193.940 47.310 194.670 47.480 ;
        RECT 195.085 48.080 198.395 48.320 ;
        RECT 198.565 48.110 198.825 49.220 ;
        RECT 195.085 47.490 196.055 48.080 ;
        RECT 198.995 47.910 199.245 49.045 ;
        RECT 199.425 48.110 199.720 49.220 ;
        RECT 200.820 48.055 201.110 49.220 ;
        RECT 201.280 48.130 204.790 49.220 ;
        RECT 196.225 47.660 199.245 47.910 ;
        RECT 195.085 47.320 198.395 47.490 ;
        RECT 193.475 46.670 193.770 47.195 ;
        RECT 193.940 46.865 194.165 47.310 ;
        RECT 194.335 46.670 194.665 47.140 ;
        RECT 195.085 46.670 195.385 47.150 ;
        RECT 195.555 46.865 195.815 47.320 ;
        RECT 195.985 46.670 196.245 47.150 ;
        RECT 196.415 46.865 196.675 47.320 ;
        RECT 196.845 46.670 197.105 47.150 ;
        RECT 197.275 46.865 197.535 47.320 ;
        RECT 197.705 46.670 197.965 47.150 ;
        RECT 198.135 46.865 198.395 47.320 ;
        RECT 198.565 46.670 198.825 47.195 ;
        RECT 198.995 46.850 199.245 47.660 ;
        RECT 199.415 47.300 199.730 47.910 ;
        RECT 201.280 47.440 202.930 47.960 ;
        RECT 203.100 47.610 204.790 48.130 ;
        RECT 204.965 48.030 205.220 48.910 ;
        RECT 205.390 48.080 205.695 49.220 ;
        RECT 206.035 48.840 206.365 49.220 ;
        RECT 206.545 48.670 206.715 48.960 ;
        RECT 206.885 48.760 207.135 49.220 ;
        RECT 205.915 48.500 206.715 48.670 ;
        RECT 207.305 48.710 208.175 49.050 ;
        RECT 199.425 46.670 199.670 47.130 ;
        RECT 200.820 46.670 201.110 47.395 ;
        RECT 201.280 46.670 204.790 47.440 ;
        RECT 204.965 47.380 205.175 48.030 ;
        RECT 205.915 47.910 206.085 48.500 ;
        RECT 207.305 48.330 207.475 48.710 ;
        RECT 208.410 48.590 208.580 49.050 ;
        RECT 208.750 48.760 209.120 49.220 ;
        RECT 209.415 48.620 209.585 48.960 ;
        RECT 209.755 48.790 210.085 49.220 ;
        RECT 210.320 48.620 210.490 48.960 ;
        RECT 206.255 48.160 207.475 48.330 ;
        RECT 207.645 48.250 208.105 48.540 ;
        RECT 208.410 48.420 208.970 48.590 ;
        RECT 209.415 48.450 210.490 48.620 ;
        RECT 210.660 48.720 211.340 49.050 ;
        RECT 211.555 48.720 211.805 49.050 ;
        RECT 211.975 48.760 212.225 49.220 ;
        RECT 208.800 48.280 208.970 48.420 ;
        RECT 207.645 48.240 208.610 48.250 ;
        RECT 207.305 48.070 207.475 48.160 ;
        RECT 207.935 48.080 208.610 48.240 ;
        RECT 205.345 47.880 206.085 47.910 ;
        RECT 205.345 47.580 206.260 47.880 ;
        RECT 205.935 47.405 206.260 47.580 ;
        RECT 204.965 46.850 205.220 47.380 ;
        RECT 205.390 46.670 205.695 47.130 ;
        RECT 205.940 47.050 206.260 47.405 ;
        RECT 206.430 47.620 206.970 47.990 ;
        RECT 207.305 47.900 207.710 48.070 ;
        RECT 206.430 47.220 206.670 47.620 ;
        RECT 207.150 47.450 207.370 47.730 ;
        RECT 206.840 47.280 207.370 47.450 ;
        RECT 206.840 47.050 207.010 47.280 ;
        RECT 207.540 47.120 207.710 47.900 ;
        RECT 207.880 47.290 208.230 47.910 ;
        RECT 208.400 47.290 208.610 48.080 ;
        RECT 208.800 48.110 210.300 48.280 ;
        RECT 208.800 47.420 208.970 48.110 ;
        RECT 210.660 47.940 210.830 48.720 ;
        RECT 211.635 48.590 211.805 48.720 ;
        RECT 209.140 47.770 210.830 47.940 ;
        RECT 211.000 48.160 211.465 48.550 ;
        RECT 211.635 48.420 212.030 48.590 ;
        RECT 209.140 47.590 209.310 47.770 ;
        RECT 205.940 46.880 207.010 47.050 ;
        RECT 207.180 46.670 207.370 47.110 ;
        RECT 207.540 46.840 208.490 47.120 ;
        RECT 208.800 47.030 209.060 47.420 ;
        RECT 209.480 47.350 210.270 47.600 ;
        RECT 208.710 46.860 209.060 47.030 ;
        RECT 209.270 46.670 209.600 47.130 ;
        RECT 210.475 47.060 210.645 47.770 ;
        RECT 211.000 47.570 211.170 48.160 ;
        RECT 210.815 47.350 211.170 47.570 ;
        RECT 211.340 47.350 211.690 47.970 ;
        RECT 211.860 47.060 212.030 48.420 ;
        RECT 212.395 48.250 212.720 49.035 ;
        RECT 212.200 47.200 212.660 48.250 ;
        RECT 210.475 46.890 211.330 47.060 ;
        RECT 211.535 46.890 212.030 47.060 ;
        RECT 212.200 46.670 212.530 47.030 ;
        RECT 212.890 46.930 213.060 49.050 ;
        RECT 213.230 48.720 213.560 49.220 ;
        RECT 213.730 48.550 213.985 49.050 ;
        RECT 213.235 48.380 213.985 48.550 ;
        RECT 214.165 48.550 214.420 49.050 ;
        RECT 214.590 48.720 214.920 49.220 ;
        RECT 214.165 48.380 214.915 48.550 ;
        RECT 213.235 47.390 213.465 48.380 ;
        RECT 213.635 47.560 213.985 48.210 ;
        RECT 214.165 47.560 214.515 48.210 ;
        RECT 214.685 47.390 214.915 48.380 ;
        RECT 213.235 47.220 213.985 47.390 ;
        RECT 213.230 46.670 213.560 47.050 ;
        RECT 213.730 46.930 213.985 47.220 ;
        RECT 214.165 47.220 214.915 47.390 ;
        RECT 214.165 46.930 214.420 47.220 ;
        RECT 214.590 46.670 214.920 47.050 ;
        RECT 215.090 46.930 215.260 49.050 ;
        RECT 215.430 48.250 215.755 49.035 ;
        RECT 215.925 48.760 216.175 49.220 ;
        RECT 216.345 48.720 216.595 49.050 ;
        RECT 216.810 48.720 217.490 49.050 ;
        RECT 216.345 48.590 216.515 48.720 ;
        RECT 216.120 48.420 216.515 48.590 ;
        RECT 215.490 47.200 215.950 48.250 ;
        RECT 216.120 47.060 216.290 48.420 ;
        RECT 216.685 48.160 217.150 48.550 ;
        RECT 216.460 47.350 216.810 47.970 ;
        RECT 216.980 47.570 217.150 48.160 ;
        RECT 217.320 47.940 217.490 48.720 ;
        RECT 217.660 48.620 217.830 48.960 ;
        RECT 218.065 48.790 218.395 49.220 ;
        RECT 218.565 48.620 218.735 48.960 ;
        RECT 219.030 48.760 219.400 49.220 ;
        RECT 217.660 48.450 218.735 48.620 ;
        RECT 219.570 48.590 219.740 49.050 ;
        RECT 219.975 48.710 220.845 49.050 ;
        RECT 221.015 48.760 221.265 49.220 ;
        RECT 219.180 48.420 219.740 48.590 ;
        RECT 219.180 48.280 219.350 48.420 ;
        RECT 217.850 48.110 219.350 48.280 ;
        RECT 220.045 48.250 220.505 48.540 ;
        RECT 217.320 47.770 219.010 47.940 ;
        RECT 216.980 47.350 217.335 47.570 ;
        RECT 217.505 47.060 217.675 47.770 ;
        RECT 217.880 47.350 218.670 47.600 ;
        RECT 218.840 47.590 219.010 47.770 ;
        RECT 219.180 47.420 219.350 48.110 ;
        RECT 215.620 46.670 215.950 47.030 ;
        RECT 216.120 46.890 216.615 47.060 ;
        RECT 216.820 46.890 217.675 47.060 ;
        RECT 218.550 46.670 218.880 47.130 ;
        RECT 219.090 47.030 219.350 47.420 ;
        RECT 219.540 48.240 220.505 48.250 ;
        RECT 220.675 48.330 220.845 48.710 ;
        RECT 221.435 48.670 221.605 48.960 ;
        RECT 221.785 48.840 222.115 49.220 ;
        RECT 221.435 48.500 222.235 48.670 ;
        RECT 219.540 48.080 220.215 48.240 ;
        RECT 220.675 48.160 221.895 48.330 ;
        RECT 219.540 47.290 219.750 48.080 ;
        RECT 220.675 48.070 220.845 48.160 ;
        RECT 219.920 47.290 220.270 47.910 ;
        RECT 220.440 47.900 220.845 48.070 ;
        RECT 220.440 47.120 220.610 47.900 ;
        RECT 220.780 47.450 221.000 47.730 ;
        RECT 221.180 47.620 221.720 47.990 ;
        RECT 222.065 47.910 222.235 48.500 ;
        RECT 222.455 48.080 222.760 49.220 ;
        RECT 222.930 48.030 223.185 48.910 ;
        RECT 223.360 48.130 225.950 49.220 ;
        RECT 222.065 47.880 222.805 47.910 ;
        RECT 220.780 47.280 221.310 47.450 ;
        RECT 219.090 46.860 219.440 47.030 ;
        RECT 219.660 46.840 220.610 47.120 ;
        RECT 220.780 46.670 220.970 47.110 ;
        RECT 221.140 47.050 221.310 47.280 ;
        RECT 221.480 47.220 221.720 47.620 ;
        RECT 221.890 47.580 222.805 47.880 ;
        RECT 221.890 47.405 222.215 47.580 ;
        RECT 221.890 47.050 222.210 47.405 ;
        RECT 222.975 47.380 223.185 48.030 ;
        RECT 221.140 46.880 222.210 47.050 ;
        RECT 222.455 46.670 222.760 47.130 ;
        RECT 222.930 46.850 223.185 47.380 ;
        RECT 223.360 47.440 224.570 47.960 ;
        RECT 224.740 47.610 225.950 48.130 ;
        RECT 226.580 48.055 226.870 49.220 ;
        RECT 227.040 48.130 229.630 49.220 ;
        RECT 230.265 48.550 230.520 49.050 ;
        RECT 230.690 48.720 231.020 49.220 ;
        RECT 230.265 48.380 231.015 48.550 ;
        RECT 227.040 47.440 228.250 47.960 ;
        RECT 228.420 47.610 229.630 48.130 ;
        RECT 230.265 47.560 230.615 48.210 ;
        RECT 223.360 46.670 225.950 47.440 ;
        RECT 226.580 46.670 226.870 47.395 ;
        RECT 227.040 46.670 229.630 47.440 ;
        RECT 230.785 47.390 231.015 48.380 ;
        RECT 230.265 47.220 231.015 47.390 ;
        RECT 230.265 46.930 230.520 47.220 ;
        RECT 230.690 46.670 231.020 47.050 ;
        RECT 231.190 46.930 231.360 49.050 ;
        RECT 231.530 48.250 231.855 49.035 ;
        RECT 232.025 48.760 232.275 49.220 ;
        RECT 232.445 48.720 232.695 49.050 ;
        RECT 232.910 48.720 233.590 49.050 ;
        RECT 232.445 48.590 232.615 48.720 ;
        RECT 232.220 48.420 232.615 48.590 ;
        RECT 231.590 47.200 232.050 48.250 ;
        RECT 232.220 47.060 232.390 48.420 ;
        RECT 232.785 48.160 233.250 48.550 ;
        RECT 232.560 47.350 232.910 47.970 ;
        RECT 233.080 47.570 233.250 48.160 ;
        RECT 233.420 47.940 233.590 48.720 ;
        RECT 233.760 48.620 233.930 48.960 ;
        RECT 234.165 48.790 234.495 49.220 ;
        RECT 234.665 48.620 234.835 48.960 ;
        RECT 235.130 48.760 235.500 49.220 ;
        RECT 233.760 48.450 234.835 48.620 ;
        RECT 235.670 48.590 235.840 49.050 ;
        RECT 236.075 48.710 236.945 49.050 ;
        RECT 237.115 48.760 237.365 49.220 ;
        RECT 235.280 48.420 235.840 48.590 ;
        RECT 235.280 48.280 235.450 48.420 ;
        RECT 233.950 48.110 235.450 48.280 ;
        RECT 236.145 48.250 236.605 48.540 ;
        RECT 233.420 47.770 235.110 47.940 ;
        RECT 233.080 47.350 233.435 47.570 ;
        RECT 233.605 47.060 233.775 47.770 ;
        RECT 233.980 47.350 234.770 47.600 ;
        RECT 234.940 47.590 235.110 47.770 ;
        RECT 235.280 47.420 235.450 48.110 ;
        RECT 231.720 46.670 232.050 47.030 ;
        RECT 232.220 46.890 232.715 47.060 ;
        RECT 232.920 46.890 233.775 47.060 ;
        RECT 234.650 46.670 234.980 47.130 ;
        RECT 235.190 47.030 235.450 47.420 ;
        RECT 235.640 48.240 236.605 48.250 ;
        RECT 236.775 48.330 236.945 48.710 ;
        RECT 237.535 48.670 237.705 48.960 ;
        RECT 237.885 48.840 238.215 49.220 ;
        RECT 237.535 48.500 238.335 48.670 ;
        RECT 235.640 48.080 236.315 48.240 ;
        RECT 236.775 48.160 237.995 48.330 ;
        RECT 235.640 47.290 235.850 48.080 ;
        RECT 236.775 48.070 236.945 48.160 ;
        RECT 236.020 47.290 236.370 47.910 ;
        RECT 236.540 47.900 236.945 48.070 ;
        RECT 236.540 47.120 236.710 47.900 ;
        RECT 236.880 47.450 237.100 47.730 ;
        RECT 237.280 47.620 237.820 47.990 ;
        RECT 238.165 47.910 238.335 48.500 ;
        RECT 238.555 48.080 238.860 49.220 ;
        RECT 239.030 48.030 239.285 48.910 ;
        RECT 239.460 48.130 241.130 49.220 ;
        RECT 241.305 48.550 241.560 49.050 ;
        RECT 241.730 48.720 242.060 49.220 ;
        RECT 241.305 48.380 242.055 48.550 ;
        RECT 238.165 47.880 238.905 47.910 ;
        RECT 236.880 47.280 237.410 47.450 ;
        RECT 235.190 46.860 235.540 47.030 ;
        RECT 235.760 46.840 236.710 47.120 ;
        RECT 236.880 46.670 237.070 47.110 ;
        RECT 237.240 47.050 237.410 47.280 ;
        RECT 237.580 47.220 237.820 47.620 ;
        RECT 237.990 47.580 238.905 47.880 ;
        RECT 237.990 47.405 238.315 47.580 ;
        RECT 237.990 47.050 238.310 47.405 ;
        RECT 239.075 47.380 239.285 48.030 ;
        RECT 237.240 46.880 238.310 47.050 ;
        RECT 238.555 46.670 238.860 47.130 ;
        RECT 239.030 46.850 239.285 47.380 ;
        RECT 239.460 47.440 240.210 47.960 ;
        RECT 240.380 47.610 241.130 48.130 ;
        RECT 241.305 47.560 241.655 48.210 ;
        RECT 239.460 46.670 241.130 47.440 ;
        RECT 241.825 47.390 242.055 48.380 ;
        RECT 241.305 47.220 242.055 47.390 ;
        RECT 241.305 46.930 241.560 47.220 ;
        RECT 241.730 46.670 242.060 47.050 ;
        RECT 242.230 46.930 242.400 49.050 ;
        RECT 242.570 48.250 242.895 49.035 ;
        RECT 243.065 48.760 243.315 49.220 ;
        RECT 243.485 48.720 243.735 49.050 ;
        RECT 243.950 48.720 244.630 49.050 ;
        RECT 243.485 48.590 243.655 48.720 ;
        RECT 243.260 48.420 243.655 48.590 ;
        RECT 242.630 47.200 243.090 48.250 ;
        RECT 243.260 47.060 243.430 48.420 ;
        RECT 243.825 48.160 244.290 48.550 ;
        RECT 243.600 47.350 243.950 47.970 ;
        RECT 244.120 47.570 244.290 48.160 ;
        RECT 244.460 47.940 244.630 48.720 ;
        RECT 244.800 48.620 244.970 48.960 ;
        RECT 245.205 48.790 245.535 49.220 ;
        RECT 245.705 48.620 245.875 48.960 ;
        RECT 246.170 48.760 246.540 49.220 ;
        RECT 244.800 48.450 245.875 48.620 ;
        RECT 246.710 48.590 246.880 49.050 ;
        RECT 247.115 48.710 247.985 49.050 ;
        RECT 248.155 48.760 248.405 49.220 ;
        RECT 246.320 48.420 246.880 48.590 ;
        RECT 246.320 48.280 246.490 48.420 ;
        RECT 244.990 48.110 246.490 48.280 ;
        RECT 247.185 48.250 247.645 48.540 ;
        RECT 244.460 47.770 246.150 47.940 ;
        RECT 244.120 47.350 244.475 47.570 ;
        RECT 244.645 47.060 244.815 47.770 ;
        RECT 245.020 47.350 245.810 47.600 ;
        RECT 245.980 47.590 246.150 47.770 ;
        RECT 246.320 47.420 246.490 48.110 ;
        RECT 242.760 46.670 243.090 47.030 ;
        RECT 243.260 46.890 243.755 47.060 ;
        RECT 243.960 46.890 244.815 47.060 ;
        RECT 245.690 46.670 246.020 47.130 ;
        RECT 246.230 47.030 246.490 47.420 ;
        RECT 246.680 48.240 247.645 48.250 ;
        RECT 247.815 48.330 247.985 48.710 ;
        RECT 248.575 48.670 248.745 48.960 ;
        RECT 248.925 48.840 249.255 49.220 ;
        RECT 248.575 48.500 249.375 48.670 ;
        RECT 246.680 48.080 247.355 48.240 ;
        RECT 247.815 48.160 249.035 48.330 ;
        RECT 246.680 47.290 246.890 48.080 ;
        RECT 247.815 48.070 247.985 48.160 ;
        RECT 247.060 47.290 247.410 47.910 ;
        RECT 247.580 47.900 247.985 48.070 ;
        RECT 247.580 47.120 247.750 47.900 ;
        RECT 247.920 47.450 248.140 47.730 ;
        RECT 248.320 47.620 248.860 47.990 ;
        RECT 249.205 47.910 249.375 48.500 ;
        RECT 249.595 48.080 249.900 49.220 ;
        RECT 250.070 48.030 250.325 48.910 ;
        RECT 250.500 48.130 252.170 49.220 ;
        RECT 249.205 47.880 249.945 47.910 ;
        RECT 247.920 47.280 248.450 47.450 ;
        RECT 246.230 46.860 246.580 47.030 ;
        RECT 246.800 46.840 247.750 47.120 ;
        RECT 247.920 46.670 248.110 47.110 ;
        RECT 248.280 47.050 248.450 47.280 ;
        RECT 248.620 47.220 248.860 47.620 ;
        RECT 249.030 47.580 249.945 47.880 ;
        RECT 249.030 47.405 249.355 47.580 ;
        RECT 249.030 47.050 249.350 47.405 ;
        RECT 250.115 47.380 250.325 48.030 ;
        RECT 248.280 46.880 249.350 47.050 ;
        RECT 249.595 46.670 249.900 47.130 ;
        RECT 250.070 46.850 250.325 47.380 ;
        RECT 250.500 47.440 251.250 47.960 ;
        RECT 251.420 47.610 252.170 48.130 ;
        RECT 252.340 48.055 252.630 49.220 ;
        RECT 252.800 48.130 254.470 49.220 ;
        RECT 254.645 48.550 254.900 49.050 ;
        RECT 255.070 48.720 255.400 49.220 ;
        RECT 254.645 48.380 255.395 48.550 ;
        RECT 252.800 47.440 253.550 47.960 ;
        RECT 253.720 47.610 254.470 48.130 ;
        RECT 254.645 47.560 254.995 48.210 ;
        RECT 250.500 46.670 252.170 47.440 ;
        RECT 252.340 46.670 252.630 47.395 ;
        RECT 252.800 46.670 254.470 47.440 ;
        RECT 255.165 47.390 255.395 48.380 ;
        RECT 254.645 47.220 255.395 47.390 ;
        RECT 254.645 46.930 254.900 47.220 ;
        RECT 255.070 46.670 255.400 47.050 ;
        RECT 255.570 46.930 255.740 49.050 ;
        RECT 255.910 48.250 256.235 49.035 ;
        RECT 256.405 48.760 256.655 49.220 ;
        RECT 256.825 48.720 257.075 49.050 ;
        RECT 257.290 48.720 257.970 49.050 ;
        RECT 256.825 48.590 256.995 48.720 ;
        RECT 256.600 48.420 256.995 48.590 ;
        RECT 255.970 47.200 256.430 48.250 ;
        RECT 256.600 47.060 256.770 48.420 ;
        RECT 257.165 48.160 257.630 48.550 ;
        RECT 256.940 47.350 257.290 47.970 ;
        RECT 257.460 47.570 257.630 48.160 ;
        RECT 257.800 47.940 257.970 48.720 ;
        RECT 258.140 48.620 258.310 48.960 ;
        RECT 258.545 48.790 258.875 49.220 ;
        RECT 259.045 48.620 259.215 48.960 ;
        RECT 259.510 48.760 259.880 49.220 ;
        RECT 258.140 48.450 259.215 48.620 ;
        RECT 260.050 48.590 260.220 49.050 ;
        RECT 260.455 48.710 261.325 49.050 ;
        RECT 261.495 48.760 261.745 49.220 ;
        RECT 259.660 48.420 260.220 48.590 ;
        RECT 259.660 48.280 259.830 48.420 ;
        RECT 258.330 48.110 259.830 48.280 ;
        RECT 260.525 48.250 260.985 48.540 ;
        RECT 257.800 47.770 259.490 47.940 ;
        RECT 257.460 47.350 257.815 47.570 ;
        RECT 257.985 47.060 258.155 47.770 ;
        RECT 258.360 47.350 259.150 47.600 ;
        RECT 259.320 47.590 259.490 47.770 ;
        RECT 259.660 47.420 259.830 48.110 ;
        RECT 256.100 46.670 256.430 47.030 ;
        RECT 256.600 46.890 257.095 47.060 ;
        RECT 257.300 46.890 258.155 47.060 ;
        RECT 259.030 46.670 259.360 47.130 ;
        RECT 259.570 47.030 259.830 47.420 ;
        RECT 260.020 48.240 260.985 48.250 ;
        RECT 261.155 48.330 261.325 48.710 ;
        RECT 261.915 48.670 262.085 48.960 ;
        RECT 262.265 48.840 262.595 49.220 ;
        RECT 261.915 48.500 262.715 48.670 ;
        RECT 260.020 48.080 260.695 48.240 ;
        RECT 261.155 48.160 262.375 48.330 ;
        RECT 260.020 47.290 260.230 48.080 ;
        RECT 261.155 48.070 261.325 48.160 ;
        RECT 260.400 47.290 260.750 47.910 ;
        RECT 260.920 47.900 261.325 48.070 ;
        RECT 260.920 47.120 261.090 47.900 ;
        RECT 261.260 47.450 261.480 47.730 ;
        RECT 261.660 47.620 262.200 47.990 ;
        RECT 262.545 47.910 262.715 48.500 ;
        RECT 262.935 48.080 263.240 49.220 ;
        RECT 263.410 48.030 263.665 48.910 ;
        RECT 262.545 47.880 263.285 47.910 ;
        RECT 261.260 47.280 261.790 47.450 ;
        RECT 259.570 46.860 259.920 47.030 ;
        RECT 260.140 46.840 261.090 47.120 ;
        RECT 261.260 46.670 261.450 47.110 ;
        RECT 261.620 47.050 261.790 47.280 ;
        RECT 261.960 47.220 262.200 47.620 ;
        RECT 262.370 47.580 263.285 47.880 ;
        RECT 262.370 47.405 262.695 47.580 ;
        RECT 262.370 47.050 262.690 47.405 ;
        RECT 263.455 47.380 263.665 48.030 ;
        RECT 261.620 46.880 262.690 47.050 ;
        RECT 262.935 46.670 263.240 47.130 ;
        RECT 263.410 46.850 263.665 47.380 ;
        RECT 263.840 48.080 264.225 49.050 ;
        RECT 264.395 48.760 264.720 49.220 ;
        RECT 265.240 48.590 265.520 49.050 ;
        RECT 264.395 48.370 265.520 48.590 ;
        RECT 263.840 47.410 264.120 48.080 ;
        RECT 264.395 47.910 264.845 48.370 ;
        RECT 265.710 48.200 266.110 49.050 ;
        RECT 266.510 48.760 266.780 49.220 ;
        RECT 266.950 48.590 267.235 49.050 ;
        RECT 264.290 47.580 264.845 47.910 ;
        RECT 265.015 47.640 266.110 48.200 ;
        RECT 264.395 47.470 264.845 47.580 ;
        RECT 263.840 46.840 264.225 47.410 ;
        RECT 264.395 47.300 265.520 47.470 ;
        RECT 264.395 46.670 264.720 47.130 ;
        RECT 265.240 46.840 265.520 47.300 ;
        RECT 265.710 46.840 266.110 47.640 ;
        RECT 266.280 48.370 267.235 48.590 ;
        RECT 266.280 47.470 266.490 48.370 ;
        RECT 267.610 48.210 267.780 49.050 ;
        RECT 267.950 48.880 269.120 49.050 ;
        RECT 267.950 48.380 268.280 48.880 ;
        RECT 268.790 48.840 269.120 48.880 ;
        RECT 269.310 48.800 269.665 49.220 ;
        RECT 268.450 48.620 268.680 48.710 ;
        RECT 269.835 48.620 270.085 49.050 ;
        RECT 268.450 48.380 270.085 48.620 ;
        RECT 270.255 48.460 270.585 49.220 ;
        RECT 270.755 48.380 271.010 49.050 ;
        RECT 266.660 47.640 267.350 48.200 ;
        RECT 267.610 48.040 270.670 48.210 ;
        RECT 267.525 47.660 267.875 47.870 ;
        RECT 268.045 47.660 268.490 47.860 ;
        RECT 268.660 47.660 269.135 47.860 ;
        RECT 266.280 47.300 267.235 47.470 ;
        RECT 266.510 46.670 266.780 47.130 ;
        RECT 266.950 46.840 267.235 47.300 ;
        RECT 267.610 47.320 268.675 47.490 ;
        RECT 267.610 46.840 267.780 47.320 ;
        RECT 267.950 46.670 268.280 47.150 ;
        RECT 268.505 47.090 268.675 47.320 ;
        RECT 268.855 47.260 269.135 47.660 ;
        RECT 269.405 47.660 269.735 47.860 ;
        RECT 269.905 47.660 270.270 47.860 ;
        RECT 269.405 47.260 269.690 47.660 ;
        RECT 270.500 47.490 270.670 48.040 ;
        RECT 269.870 47.320 270.670 47.490 ;
        RECT 269.870 47.090 270.040 47.320 ;
        RECT 270.840 47.250 271.010 48.380 ;
        RECT 271.200 48.130 273.790 49.220 ;
        RECT 270.825 47.170 271.010 47.250 ;
        RECT 268.505 46.840 270.040 47.090 ;
        RECT 270.210 46.670 270.540 47.150 ;
        RECT 270.755 46.840 271.010 47.170 ;
        RECT 271.200 47.440 272.410 47.960 ;
        RECT 272.580 47.610 273.790 48.130 ;
        RECT 274.420 48.080 274.805 49.050 ;
        RECT 274.975 48.760 275.300 49.220 ;
        RECT 275.820 48.590 276.100 49.050 ;
        RECT 274.975 48.370 276.100 48.590 ;
        RECT 271.200 46.670 273.790 47.440 ;
        RECT 274.420 47.410 274.700 48.080 ;
        RECT 274.975 47.910 275.425 48.370 ;
        RECT 276.290 48.200 276.690 49.050 ;
        RECT 277.090 48.760 277.360 49.220 ;
        RECT 277.530 48.590 277.815 49.050 ;
        RECT 274.870 47.580 275.425 47.910 ;
        RECT 275.595 47.640 276.690 48.200 ;
        RECT 274.975 47.470 275.425 47.580 ;
        RECT 274.420 46.840 274.805 47.410 ;
        RECT 274.975 47.300 276.100 47.470 ;
        RECT 274.975 46.670 275.300 47.130 ;
        RECT 275.820 46.840 276.100 47.300 ;
        RECT 276.290 46.840 276.690 47.640 ;
        RECT 276.860 48.370 277.815 48.590 ;
        RECT 276.860 47.470 277.070 48.370 ;
        RECT 277.240 47.640 277.930 48.200 ;
        RECT 278.100 48.055 278.390 49.220 ;
        RECT 278.565 48.030 278.820 48.910 ;
        RECT 278.990 48.080 279.295 49.220 ;
        RECT 279.635 48.840 279.965 49.220 ;
        RECT 280.145 48.670 280.315 48.960 ;
        RECT 280.485 48.760 280.735 49.220 ;
        RECT 279.515 48.500 280.315 48.670 ;
        RECT 280.905 48.710 281.775 49.050 ;
        RECT 276.860 47.300 277.815 47.470 ;
        RECT 277.090 46.670 277.360 47.130 ;
        RECT 277.530 46.840 277.815 47.300 ;
        RECT 278.100 46.670 278.390 47.395 ;
        RECT 278.565 47.380 278.775 48.030 ;
        RECT 279.515 47.910 279.685 48.500 ;
        RECT 280.905 48.330 281.075 48.710 ;
        RECT 282.010 48.590 282.180 49.050 ;
        RECT 282.350 48.760 282.720 49.220 ;
        RECT 283.015 48.620 283.185 48.960 ;
        RECT 283.355 48.790 283.685 49.220 ;
        RECT 283.920 48.620 284.090 48.960 ;
        RECT 279.855 48.160 281.075 48.330 ;
        RECT 281.245 48.250 281.705 48.540 ;
        RECT 282.010 48.420 282.570 48.590 ;
        RECT 283.015 48.450 284.090 48.620 ;
        RECT 284.260 48.720 284.940 49.050 ;
        RECT 285.155 48.720 285.405 49.050 ;
        RECT 285.575 48.760 285.825 49.220 ;
        RECT 282.400 48.280 282.570 48.420 ;
        RECT 281.245 48.240 282.210 48.250 ;
        RECT 280.905 48.070 281.075 48.160 ;
        RECT 281.535 48.080 282.210 48.240 ;
        RECT 278.945 47.880 279.685 47.910 ;
        RECT 278.945 47.580 279.860 47.880 ;
        RECT 279.535 47.405 279.860 47.580 ;
        RECT 278.565 46.850 278.820 47.380 ;
        RECT 278.990 46.670 279.295 47.130 ;
        RECT 279.540 47.050 279.860 47.405 ;
        RECT 280.030 47.620 280.570 47.990 ;
        RECT 280.905 47.900 281.310 48.070 ;
        RECT 280.030 47.220 280.270 47.620 ;
        RECT 280.750 47.450 280.970 47.730 ;
        RECT 280.440 47.280 280.970 47.450 ;
        RECT 280.440 47.050 280.610 47.280 ;
        RECT 281.140 47.120 281.310 47.900 ;
        RECT 281.480 47.290 281.830 47.910 ;
        RECT 282.000 47.290 282.210 48.080 ;
        RECT 282.400 48.110 283.900 48.280 ;
        RECT 282.400 47.420 282.570 48.110 ;
        RECT 284.260 47.940 284.430 48.720 ;
        RECT 285.235 48.590 285.405 48.720 ;
        RECT 282.740 47.770 284.430 47.940 ;
        RECT 284.600 48.160 285.065 48.550 ;
        RECT 285.235 48.420 285.630 48.590 ;
        RECT 282.740 47.590 282.910 47.770 ;
        RECT 279.540 46.880 280.610 47.050 ;
        RECT 280.780 46.670 280.970 47.110 ;
        RECT 281.140 46.840 282.090 47.120 ;
        RECT 282.400 47.030 282.660 47.420 ;
        RECT 283.080 47.350 283.870 47.600 ;
        RECT 282.310 46.860 282.660 47.030 ;
        RECT 282.870 46.670 283.200 47.130 ;
        RECT 284.075 47.060 284.245 47.770 ;
        RECT 284.600 47.570 284.770 48.160 ;
        RECT 284.415 47.350 284.770 47.570 ;
        RECT 284.940 47.350 285.290 47.970 ;
        RECT 285.460 47.060 285.630 48.420 ;
        RECT 285.995 48.250 286.320 49.035 ;
        RECT 285.800 47.200 286.260 48.250 ;
        RECT 284.075 46.890 284.930 47.060 ;
        RECT 285.135 46.890 285.630 47.060 ;
        RECT 285.800 46.670 286.130 47.030 ;
        RECT 286.490 46.930 286.660 49.050 ;
        RECT 286.830 48.720 287.160 49.220 ;
        RECT 287.330 48.550 287.585 49.050 ;
        RECT 286.835 48.380 287.585 48.550 ;
        RECT 287.765 48.550 288.020 49.050 ;
        RECT 288.190 48.720 288.520 49.220 ;
        RECT 287.765 48.380 288.515 48.550 ;
        RECT 286.835 47.390 287.065 48.380 ;
        RECT 287.235 47.560 287.585 48.210 ;
        RECT 287.765 47.560 288.115 48.210 ;
        RECT 288.285 47.390 288.515 48.380 ;
        RECT 286.835 47.220 287.585 47.390 ;
        RECT 286.830 46.670 287.160 47.050 ;
        RECT 287.330 46.930 287.585 47.220 ;
        RECT 287.765 47.220 288.515 47.390 ;
        RECT 287.765 46.930 288.020 47.220 ;
        RECT 288.190 46.670 288.520 47.050 ;
        RECT 288.690 46.930 288.860 49.050 ;
        RECT 289.030 48.250 289.355 49.035 ;
        RECT 289.525 48.760 289.775 49.220 ;
        RECT 289.945 48.720 290.195 49.050 ;
        RECT 290.410 48.720 291.090 49.050 ;
        RECT 289.945 48.590 290.115 48.720 ;
        RECT 289.720 48.420 290.115 48.590 ;
        RECT 289.090 47.200 289.550 48.250 ;
        RECT 289.720 47.060 289.890 48.420 ;
        RECT 290.285 48.160 290.750 48.550 ;
        RECT 290.060 47.350 290.410 47.970 ;
        RECT 290.580 47.570 290.750 48.160 ;
        RECT 290.920 47.940 291.090 48.720 ;
        RECT 291.260 48.620 291.430 48.960 ;
        RECT 291.665 48.790 291.995 49.220 ;
        RECT 292.165 48.620 292.335 48.960 ;
        RECT 292.630 48.760 293.000 49.220 ;
        RECT 291.260 48.450 292.335 48.620 ;
        RECT 293.170 48.590 293.340 49.050 ;
        RECT 293.575 48.710 294.445 49.050 ;
        RECT 294.615 48.760 294.865 49.220 ;
        RECT 292.780 48.420 293.340 48.590 ;
        RECT 292.780 48.280 292.950 48.420 ;
        RECT 291.450 48.110 292.950 48.280 ;
        RECT 293.645 48.250 294.105 48.540 ;
        RECT 290.920 47.770 292.610 47.940 ;
        RECT 290.580 47.350 290.935 47.570 ;
        RECT 291.105 47.060 291.275 47.770 ;
        RECT 291.480 47.350 292.270 47.600 ;
        RECT 292.440 47.590 292.610 47.770 ;
        RECT 292.780 47.420 292.950 48.110 ;
        RECT 289.220 46.670 289.550 47.030 ;
        RECT 289.720 46.890 290.215 47.060 ;
        RECT 290.420 46.890 291.275 47.060 ;
        RECT 292.150 46.670 292.480 47.130 ;
        RECT 292.690 47.030 292.950 47.420 ;
        RECT 293.140 48.240 294.105 48.250 ;
        RECT 294.275 48.330 294.445 48.710 ;
        RECT 295.035 48.670 295.205 48.960 ;
        RECT 295.385 48.840 295.715 49.220 ;
        RECT 295.035 48.500 295.835 48.670 ;
        RECT 293.140 48.080 293.815 48.240 ;
        RECT 294.275 48.160 295.495 48.330 ;
        RECT 293.140 47.290 293.350 48.080 ;
        RECT 294.275 48.070 294.445 48.160 ;
        RECT 293.520 47.290 293.870 47.910 ;
        RECT 294.040 47.900 294.445 48.070 ;
        RECT 294.040 47.120 294.210 47.900 ;
        RECT 294.380 47.450 294.600 47.730 ;
        RECT 294.780 47.620 295.320 47.990 ;
        RECT 295.665 47.910 295.835 48.500 ;
        RECT 296.055 48.080 296.360 49.220 ;
        RECT 296.530 48.030 296.785 48.910 ;
        RECT 297.995 48.590 298.280 49.050 ;
        RECT 298.450 48.760 298.720 49.220 ;
        RECT 297.995 48.370 298.950 48.590 ;
        RECT 295.665 47.880 296.405 47.910 ;
        RECT 294.380 47.280 294.910 47.450 ;
        RECT 292.690 46.860 293.040 47.030 ;
        RECT 293.260 46.840 294.210 47.120 ;
        RECT 294.380 46.670 294.570 47.110 ;
        RECT 294.740 47.050 294.910 47.280 ;
        RECT 295.080 47.220 295.320 47.620 ;
        RECT 295.490 47.580 296.405 47.880 ;
        RECT 295.490 47.405 295.815 47.580 ;
        RECT 295.490 47.050 295.810 47.405 ;
        RECT 296.575 47.380 296.785 48.030 ;
        RECT 297.880 47.640 298.570 48.200 ;
        RECT 298.740 47.470 298.950 48.370 ;
        RECT 294.740 46.880 295.810 47.050 ;
        RECT 296.055 46.670 296.360 47.130 ;
        RECT 296.530 46.850 296.785 47.380 ;
        RECT 297.995 47.300 298.950 47.470 ;
        RECT 299.120 48.200 299.520 49.050 ;
        RECT 299.710 48.590 299.990 49.050 ;
        RECT 300.510 48.760 300.835 49.220 ;
        RECT 299.710 48.370 300.835 48.590 ;
        RECT 299.120 47.640 300.215 48.200 ;
        RECT 300.385 47.910 300.835 48.370 ;
        RECT 301.005 48.080 301.390 49.050 ;
        RECT 301.560 48.130 303.230 49.220 ;
        RECT 297.995 46.840 298.280 47.300 ;
        RECT 298.450 46.670 298.720 47.130 ;
        RECT 299.120 46.840 299.520 47.640 ;
        RECT 300.385 47.580 300.940 47.910 ;
        RECT 300.385 47.470 300.835 47.580 ;
        RECT 299.710 47.300 300.835 47.470 ;
        RECT 301.110 47.410 301.390 48.080 ;
        RECT 299.710 46.840 299.990 47.300 ;
        RECT 300.510 46.670 300.835 47.130 ;
        RECT 301.005 46.840 301.390 47.410 ;
        RECT 301.560 47.440 302.310 47.960 ;
        RECT 302.480 47.610 303.230 48.130 ;
        RECT 303.860 48.055 304.150 49.220 ;
        RECT 304.320 48.785 309.665 49.220 ;
        RECT 301.560 46.670 303.230 47.440 ;
        RECT 303.860 46.670 304.150 47.395 ;
        RECT 305.905 47.215 306.245 48.045 ;
        RECT 307.725 47.535 308.075 48.785 ;
        RECT 309.840 48.130 311.050 49.220 ;
        RECT 309.840 47.590 310.360 48.130 ;
        RECT 310.530 47.420 311.050 47.960 ;
        RECT 304.320 46.670 309.665 47.215 ;
        RECT 309.840 46.670 311.050 47.420 ;
        RECT 162.095 46.500 311.135 46.670 ;
        RECT 162.180 45.750 163.390 46.500 ;
        RECT 163.560 45.955 168.905 46.500 ;
        RECT 162.180 45.210 162.700 45.750 ;
        RECT 162.870 45.040 163.390 45.580 ;
        RECT 165.145 45.125 165.485 45.955 ;
        RECT 169.080 45.730 171.670 46.500 ;
        RECT 171.845 45.950 172.100 46.240 ;
        RECT 172.270 46.120 172.600 46.500 ;
        RECT 171.845 45.780 172.595 45.950 ;
        RECT 162.180 43.950 163.390 45.040 ;
        RECT 166.965 44.385 167.315 45.635 ;
        RECT 169.080 45.210 170.290 45.730 ;
        RECT 170.460 45.040 171.670 45.560 ;
        RECT 163.560 43.950 168.905 44.385 ;
        RECT 169.080 43.950 171.670 45.040 ;
        RECT 171.845 44.960 172.195 45.610 ;
        RECT 172.365 44.790 172.595 45.780 ;
        RECT 171.845 44.620 172.595 44.790 ;
        RECT 171.845 44.120 172.100 44.620 ;
        RECT 172.270 43.950 172.600 44.450 ;
        RECT 172.770 44.120 172.940 46.240 ;
        RECT 173.300 46.140 173.630 46.500 ;
        RECT 173.800 46.110 174.295 46.280 ;
        RECT 174.500 46.110 175.355 46.280 ;
        RECT 173.170 44.920 173.630 45.970 ;
        RECT 173.110 44.135 173.435 44.920 ;
        RECT 173.800 44.750 173.970 46.110 ;
        RECT 174.140 45.200 174.490 45.820 ;
        RECT 174.660 45.600 175.015 45.820 ;
        RECT 174.660 45.010 174.830 45.600 ;
        RECT 175.185 45.400 175.355 46.110 ;
        RECT 176.230 46.040 176.560 46.500 ;
        RECT 176.770 46.140 177.120 46.310 ;
        RECT 175.560 45.570 176.350 45.820 ;
        RECT 176.770 45.750 177.030 46.140 ;
        RECT 177.340 46.050 178.290 46.330 ;
        RECT 178.460 46.060 178.650 46.500 ;
        RECT 178.820 46.120 179.890 46.290 ;
        RECT 176.520 45.400 176.690 45.580 ;
        RECT 173.800 44.580 174.195 44.750 ;
        RECT 174.365 44.620 174.830 45.010 ;
        RECT 175.000 45.230 176.690 45.400 ;
        RECT 174.025 44.450 174.195 44.580 ;
        RECT 175.000 44.450 175.170 45.230 ;
        RECT 176.860 45.060 177.030 45.750 ;
        RECT 175.530 44.890 177.030 45.060 ;
        RECT 177.220 45.090 177.430 45.880 ;
        RECT 177.600 45.260 177.950 45.880 ;
        RECT 178.120 45.270 178.290 46.050 ;
        RECT 178.820 45.890 178.990 46.120 ;
        RECT 178.460 45.720 178.990 45.890 ;
        RECT 178.460 45.440 178.680 45.720 ;
        RECT 179.160 45.550 179.400 45.950 ;
        RECT 178.120 45.100 178.525 45.270 ;
        RECT 178.860 45.180 179.400 45.550 ;
        RECT 179.570 45.765 179.890 46.120 ;
        RECT 180.135 46.040 180.440 46.500 ;
        RECT 180.610 45.790 180.860 46.320 ;
        RECT 179.570 45.590 179.895 45.765 ;
        RECT 179.570 45.290 180.485 45.590 ;
        RECT 179.745 45.260 180.485 45.290 ;
        RECT 177.220 44.930 177.895 45.090 ;
        RECT 178.355 45.010 178.525 45.100 ;
        RECT 177.220 44.920 178.185 44.930 ;
        RECT 176.860 44.750 177.030 44.890 ;
        RECT 173.605 43.950 173.855 44.410 ;
        RECT 174.025 44.120 174.275 44.450 ;
        RECT 174.490 44.120 175.170 44.450 ;
        RECT 175.340 44.550 176.415 44.720 ;
        RECT 176.860 44.580 177.420 44.750 ;
        RECT 177.725 44.630 178.185 44.920 ;
        RECT 178.355 44.840 179.575 45.010 ;
        RECT 175.340 44.210 175.510 44.550 ;
        RECT 175.745 43.950 176.075 44.380 ;
        RECT 176.245 44.210 176.415 44.550 ;
        RECT 176.710 43.950 177.080 44.410 ;
        RECT 177.250 44.120 177.420 44.580 ;
        RECT 178.355 44.460 178.525 44.840 ;
        RECT 179.745 44.670 179.915 45.260 ;
        RECT 180.655 45.140 180.860 45.790 ;
        RECT 181.030 45.745 181.280 46.500 ;
        RECT 181.505 45.760 181.760 46.330 ;
        RECT 181.930 46.100 182.260 46.500 ;
        RECT 182.685 45.965 183.215 46.330 ;
        RECT 183.405 46.160 183.680 46.330 ;
        RECT 183.400 45.990 183.680 46.160 ;
        RECT 182.685 45.930 182.860 45.965 ;
        RECT 181.930 45.760 182.860 45.930 ;
        RECT 177.655 44.120 178.525 44.460 ;
        RECT 179.115 44.500 179.915 44.670 ;
        RECT 178.695 43.950 178.945 44.410 ;
        RECT 179.115 44.210 179.285 44.500 ;
        RECT 179.465 43.950 179.795 44.330 ;
        RECT 180.135 43.950 180.440 45.090 ;
        RECT 180.610 44.260 180.860 45.140 ;
        RECT 181.505 45.090 181.675 45.760 ;
        RECT 181.930 45.590 182.100 45.760 ;
        RECT 181.845 45.260 182.100 45.590 ;
        RECT 182.325 45.260 182.520 45.590 ;
        RECT 181.030 43.950 181.280 45.090 ;
        RECT 181.505 44.120 181.840 45.090 ;
        RECT 182.010 43.950 182.180 45.090 ;
        RECT 182.350 44.290 182.520 45.260 ;
        RECT 182.690 44.630 182.860 45.760 ;
        RECT 183.030 44.970 183.200 45.770 ;
        RECT 183.405 45.170 183.680 45.990 ;
        RECT 183.850 44.970 184.040 46.330 ;
        RECT 184.220 45.965 184.730 46.500 ;
        RECT 184.950 45.690 185.195 46.295 ;
        RECT 185.640 45.730 187.310 46.500 ;
        RECT 187.940 45.775 188.230 46.500 ;
        RECT 189.325 45.950 189.580 46.240 ;
        RECT 189.750 46.120 190.080 46.500 ;
        RECT 189.325 45.780 190.075 45.950 ;
        RECT 184.240 45.520 185.470 45.690 ;
        RECT 183.030 44.800 184.040 44.970 ;
        RECT 184.210 44.955 184.960 45.145 ;
        RECT 182.690 44.460 183.815 44.630 ;
        RECT 184.210 44.290 184.380 44.955 ;
        RECT 185.130 44.710 185.470 45.520 ;
        RECT 185.640 45.210 186.390 45.730 ;
        RECT 186.560 45.040 187.310 45.560 ;
        RECT 182.350 44.120 184.380 44.290 ;
        RECT 184.550 43.950 184.720 44.710 ;
        RECT 184.955 44.300 185.470 44.710 ;
        RECT 185.640 43.950 187.310 45.040 ;
        RECT 187.940 43.950 188.230 45.115 ;
        RECT 189.325 44.960 189.675 45.610 ;
        RECT 189.845 44.790 190.075 45.780 ;
        RECT 189.325 44.620 190.075 44.790 ;
        RECT 189.325 44.120 189.580 44.620 ;
        RECT 189.750 43.950 190.080 44.450 ;
        RECT 190.250 44.120 190.420 46.240 ;
        RECT 190.780 46.140 191.110 46.500 ;
        RECT 191.280 46.110 191.775 46.280 ;
        RECT 191.980 46.110 192.835 46.280 ;
        RECT 190.650 44.920 191.110 45.970 ;
        RECT 190.590 44.135 190.915 44.920 ;
        RECT 191.280 44.750 191.450 46.110 ;
        RECT 191.620 45.200 191.970 45.820 ;
        RECT 192.140 45.600 192.495 45.820 ;
        RECT 192.140 45.010 192.310 45.600 ;
        RECT 192.665 45.400 192.835 46.110 ;
        RECT 193.710 46.040 194.040 46.500 ;
        RECT 194.250 46.140 194.600 46.310 ;
        RECT 193.040 45.570 193.830 45.820 ;
        RECT 194.250 45.750 194.510 46.140 ;
        RECT 194.820 46.050 195.770 46.330 ;
        RECT 195.940 46.060 196.130 46.500 ;
        RECT 196.300 46.120 197.370 46.290 ;
        RECT 194.000 45.400 194.170 45.580 ;
        RECT 191.280 44.580 191.675 44.750 ;
        RECT 191.845 44.620 192.310 45.010 ;
        RECT 192.480 45.230 194.170 45.400 ;
        RECT 191.505 44.450 191.675 44.580 ;
        RECT 192.480 44.450 192.650 45.230 ;
        RECT 194.340 45.060 194.510 45.750 ;
        RECT 193.010 44.890 194.510 45.060 ;
        RECT 194.700 45.090 194.910 45.880 ;
        RECT 195.080 45.260 195.430 45.880 ;
        RECT 195.600 45.270 195.770 46.050 ;
        RECT 196.300 45.890 196.470 46.120 ;
        RECT 195.940 45.720 196.470 45.890 ;
        RECT 195.940 45.440 196.160 45.720 ;
        RECT 196.640 45.550 196.880 45.950 ;
        RECT 195.600 45.100 196.005 45.270 ;
        RECT 196.340 45.180 196.880 45.550 ;
        RECT 197.050 45.765 197.370 46.120 ;
        RECT 197.615 46.040 197.920 46.500 ;
        RECT 198.090 45.790 198.340 46.320 ;
        RECT 197.050 45.590 197.375 45.765 ;
        RECT 197.050 45.290 197.965 45.590 ;
        RECT 197.225 45.260 197.965 45.290 ;
        RECT 194.700 44.930 195.375 45.090 ;
        RECT 195.835 45.010 196.005 45.100 ;
        RECT 194.700 44.920 195.665 44.930 ;
        RECT 194.340 44.750 194.510 44.890 ;
        RECT 191.085 43.950 191.335 44.410 ;
        RECT 191.505 44.120 191.755 44.450 ;
        RECT 191.970 44.120 192.650 44.450 ;
        RECT 192.820 44.550 193.895 44.720 ;
        RECT 194.340 44.580 194.900 44.750 ;
        RECT 195.205 44.630 195.665 44.920 ;
        RECT 195.835 44.840 197.055 45.010 ;
        RECT 192.820 44.210 192.990 44.550 ;
        RECT 193.225 43.950 193.555 44.380 ;
        RECT 193.725 44.210 193.895 44.550 ;
        RECT 194.190 43.950 194.560 44.410 ;
        RECT 194.730 44.120 194.900 44.580 ;
        RECT 195.835 44.460 196.005 44.840 ;
        RECT 197.225 44.670 197.395 45.260 ;
        RECT 198.135 45.140 198.340 45.790 ;
        RECT 198.510 45.745 198.760 46.500 ;
        RECT 200.015 45.870 200.300 46.330 ;
        RECT 200.470 46.040 200.740 46.500 ;
        RECT 200.015 45.700 200.970 45.870 ;
        RECT 195.135 44.120 196.005 44.460 ;
        RECT 196.595 44.500 197.395 44.670 ;
        RECT 196.175 43.950 196.425 44.410 ;
        RECT 196.595 44.210 196.765 44.500 ;
        RECT 196.945 43.950 197.275 44.330 ;
        RECT 197.615 43.950 197.920 45.090 ;
        RECT 198.090 44.260 198.340 45.140 ;
        RECT 198.510 43.950 198.760 45.090 ;
        RECT 199.900 44.970 200.590 45.530 ;
        RECT 200.760 44.800 200.970 45.700 ;
        RECT 200.015 44.580 200.970 44.800 ;
        RECT 201.140 45.530 201.540 46.330 ;
        RECT 201.730 45.870 202.010 46.330 ;
        RECT 202.530 46.040 202.855 46.500 ;
        RECT 201.730 45.700 202.855 45.870 ;
        RECT 203.025 45.760 203.410 46.330 ;
        RECT 202.405 45.590 202.855 45.700 ;
        RECT 201.140 44.970 202.235 45.530 ;
        RECT 202.405 45.260 202.960 45.590 ;
        RECT 200.015 44.120 200.300 44.580 ;
        RECT 200.470 43.950 200.740 44.410 ;
        RECT 201.140 44.120 201.540 44.970 ;
        RECT 202.405 44.800 202.855 45.260 ;
        RECT 203.130 45.090 203.410 45.760 ;
        RECT 201.730 44.580 202.855 44.800 ;
        RECT 201.730 44.120 202.010 44.580 ;
        RECT 202.530 43.950 202.855 44.410 ;
        RECT 203.025 44.120 203.410 45.090 ;
        RECT 203.585 45.760 203.840 46.330 ;
        RECT 204.010 46.100 204.340 46.500 ;
        RECT 204.765 45.965 205.295 46.330 ;
        RECT 204.765 45.930 204.940 45.965 ;
        RECT 204.010 45.760 204.940 45.930 ;
        RECT 203.585 45.090 203.755 45.760 ;
        RECT 204.010 45.590 204.180 45.760 ;
        RECT 203.925 45.260 204.180 45.590 ;
        RECT 204.405 45.260 204.600 45.590 ;
        RECT 203.585 44.120 203.920 45.090 ;
        RECT 204.090 43.950 204.260 45.090 ;
        RECT 204.430 44.290 204.600 45.260 ;
        RECT 204.770 44.630 204.940 45.760 ;
        RECT 205.110 44.970 205.280 45.770 ;
        RECT 205.485 45.480 205.760 46.330 ;
        RECT 205.480 45.310 205.760 45.480 ;
        RECT 205.485 45.170 205.760 45.310 ;
        RECT 205.930 44.970 206.120 46.330 ;
        RECT 206.300 45.965 206.810 46.500 ;
        RECT 207.030 45.690 207.275 46.295 ;
        RECT 207.720 45.730 209.390 46.500 ;
        RECT 206.320 45.520 207.550 45.690 ;
        RECT 205.110 44.800 206.120 44.970 ;
        RECT 206.290 44.955 207.040 45.145 ;
        RECT 204.770 44.460 205.895 44.630 ;
        RECT 206.290 44.290 206.460 44.955 ;
        RECT 207.210 44.710 207.550 45.520 ;
        RECT 207.720 45.210 208.470 45.730 ;
        RECT 209.835 45.690 210.080 46.295 ;
        RECT 210.300 45.965 210.810 46.500 ;
        RECT 208.640 45.040 209.390 45.560 ;
        RECT 204.430 44.120 206.460 44.290 ;
        RECT 206.630 43.950 206.800 44.710 ;
        RECT 207.035 44.300 207.550 44.710 ;
        RECT 207.720 43.950 209.390 45.040 ;
        RECT 209.560 45.520 210.790 45.690 ;
        RECT 209.560 44.710 209.900 45.520 ;
        RECT 210.070 44.955 210.820 45.145 ;
        RECT 209.560 44.300 210.075 44.710 ;
        RECT 210.310 43.950 210.480 44.710 ;
        RECT 210.650 44.290 210.820 44.955 ;
        RECT 210.990 44.970 211.180 46.330 ;
        RECT 211.350 45.480 211.625 46.330 ;
        RECT 211.815 45.965 212.345 46.330 ;
        RECT 212.770 46.100 213.100 46.500 ;
        RECT 212.170 45.930 212.345 45.965 ;
        RECT 211.350 45.310 211.630 45.480 ;
        RECT 211.350 45.170 211.625 45.310 ;
        RECT 211.830 44.970 212.000 45.770 ;
        RECT 210.990 44.800 212.000 44.970 ;
        RECT 212.170 45.760 213.100 45.930 ;
        RECT 213.270 45.760 213.525 46.330 ;
        RECT 213.700 45.775 213.990 46.500 ;
        RECT 212.170 44.630 212.340 45.760 ;
        RECT 212.930 45.590 213.100 45.760 ;
        RECT 211.215 44.460 212.340 44.630 ;
        RECT 212.510 45.260 212.705 45.590 ;
        RECT 212.930 45.260 213.185 45.590 ;
        RECT 212.510 44.290 212.680 45.260 ;
        RECT 213.355 45.090 213.525 45.760 ;
        RECT 214.160 45.730 215.830 46.500 ;
        RECT 216.465 45.950 216.720 46.240 ;
        RECT 216.890 46.120 217.220 46.500 ;
        RECT 216.465 45.780 217.215 45.950 ;
        RECT 214.160 45.210 214.910 45.730 ;
        RECT 210.650 44.120 212.680 44.290 ;
        RECT 212.850 43.950 213.020 45.090 ;
        RECT 213.190 44.120 213.525 45.090 ;
        RECT 213.700 43.950 213.990 45.115 ;
        RECT 215.080 45.040 215.830 45.560 ;
        RECT 214.160 43.950 215.830 45.040 ;
        RECT 216.465 44.960 216.815 45.610 ;
        RECT 216.985 44.790 217.215 45.780 ;
        RECT 216.465 44.620 217.215 44.790 ;
        RECT 216.465 44.120 216.720 44.620 ;
        RECT 216.890 43.950 217.220 44.450 ;
        RECT 217.390 44.120 217.560 46.240 ;
        RECT 217.920 46.140 218.250 46.500 ;
        RECT 218.420 46.110 218.915 46.280 ;
        RECT 219.120 46.110 219.975 46.280 ;
        RECT 217.790 44.920 218.250 45.970 ;
        RECT 217.730 44.135 218.055 44.920 ;
        RECT 218.420 44.750 218.590 46.110 ;
        RECT 218.760 45.200 219.110 45.820 ;
        RECT 219.280 45.600 219.635 45.820 ;
        RECT 219.280 45.010 219.450 45.600 ;
        RECT 219.805 45.400 219.975 46.110 ;
        RECT 220.850 46.040 221.180 46.500 ;
        RECT 221.390 46.140 221.740 46.310 ;
        RECT 220.180 45.570 220.970 45.820 ;
        RECT 221.390 45.750 221.650 46.140 ;
        RECT 221.960 46.050 222.910 46.330 ;
        RECT 223.080 46.060 223.270 46.500 ;
        RECT 223.440 46.120 224.510 46.290 ;
        RECT 221.140 45.400 221.310 45.580 ;
        RECT 218.420 44.580 218.815 44.750 ;
        RECT 218.985 44.620 219.450 45.010 ;
        RECT 219.620 45.230 221.310 45.400 ;
        RECT 218.645 44.450 218.815 44.580 ;
        RECT 219.620 44.450 219.790 45.230 ;
        RECT 221.480 45.060 221.650 45.750 ;
        RECT 220.150 44.890 221.650 45.060 ;
        RECT 221.840 45.090 222.050 45.880 ;
        RECT 222.220 45.260 222.570 45.880 ;
        RECT 222.740 45.270 222.910 46.050 ;
        RECT 223.440 45.890 223.610 46.120 ;
        RECT 223.080 45.720 223.610 45.890 ;
        RECT 223.080 45.440 223.300 45.720 ;
        RECT 223.780 45.550 224.020 45.950 ;
        RECT 222.740 45.100 223.145 45.270 ;
        RECT 223.480 45.180 224.020 45.550 ;
        RECT 224.190 45.765 224.510 46.120 ;
        RECT 224.755 46.040 225.060 46.500 ;
        RECT 225.230 45.790 225.485 46.320 ;
        RECT 224.190 45.590 224.515 45.765 ;
        RECT 224.190 45.290 225.105 45.590 ;
        RECT 224.365 45.260 225.105 45.290 ;
        RECT 221.840 44.930 222.515 45.090 ;
        RECT 222.975 45.010 223.145 45.100 ;
        RECT 221.840 44.920 222.805 44.930 ;
        RECT 221.480 44.750 221.650 44.890 ;
        RECT 218.225 43.950 218.475 44.410 ;
        RECT 218.645 44.120 218.895 44.450 ;
        RECT 219.110 44.120 219.790 44.450 ;
        RECT 219.960 44.550 221.035 44.720 ;
        RECT 221.480 44.580 222.040 44.750 ;
        RECT 222.345 44.630 222.805 44.920 ;
        RECT 222.975 44.840 224.195 45.010 ;
        RECT 219.960 44.210 220.130 44.550 ;
        RECT 220.365 43.950 220.695 44.380 ;
        RECT 220.865 44.210 221.035 44.550 ;
        RECT 221.330 43.950 221.700 44.410 ;
        RECT 221.870 44.120 222.040 44.580 ;
        RECT 222.975 44.460 223.145 44.840 ;
        RECT 224.365 44.670 224.535 45.260 ;
        RECT 225.275 45.140 225.485 45.790 ;
        RECT 222.275 44.120 223.145 44.460 ;
        RECT 223.735 44.500 224.535 44.670 ;
        RECT 223.315 43.950 223.565 44.410 ;
        RECT 223.735 44.210 223.905 44.500 ;
        RECT 224.085 43.950 224.415 44.330 ;
        RECT 224.755 43.950 225.060 45.090 ;
        RECT 225.230 44.260 225.485 45.140 ;
        RECT 226.120 45.680 226.805 46.320 ;
        RECT 226.975 45.680 227.145 46.500 ;
        RECT 227.315 45.850 227.645 46.315 ;
        RECT 227.815 46.030 227.985 46.500 ;
        RECT 228.245 46.110 229.430 46.280 ;
        RECT 229.600 45.940 229.930 46.330 ;
        RECT 228.630 45.850 229.015 45.940 ;
        RECT 227.315 45.680 229.015 45.850 ;
        RECT 229.420 45.760 229.930 45.940 ;
        RECT 230.265 45.950 230.520 46.240 ;
        RECT 230.690 46.120 231.020 46.500 ;
        RECT 230.265 45.780 231.015 45.950 ;
        RECT 226.120 44.710 226.370 45.680 ;
        RECT 226.540 45.300 226.875 45.510 ;
        RECT 227.045 45.300 227.495 45.510 ;
        RECT 227.685 45.480 228.170 45.510 ;
        RECT 227.685 45.310 228.190 45.480 ;
        RECT 227.685 45.300 228.170 45.310 ;
        RECT 226.705 45.130 226.875 45.300 ;
        RECT 226.705 44.960 227.625 45.130 ;
        RECT 226.120 44.120 226.785 44.710 ;
        RECT 226.955 43.950 227.285 44.790 ;
        RECT 227.455 44.710 227.625 44.960 ;
        RECT 227.795 44.880 228.170 45.300 ;
        RECT 228.360 45.260 228.740 45.510 ;
        RECT 228.920 45.300 229.250 45.510 ;
        RECT 228.360 44.880 228.680 45.260 ;
        RECT 229.420 45.130 229.590 45.760 ;
        RECT 229.760 45.300 230.090 45.590 ;
        RECT 228.850 44.960 229.935 45.130 ;
        RECT 230.265 44.960 230.615 45.610 ;
        RECT 228.850 44.710 229.020 44.960 ;
        RECT 227.455 44.540 229.020 44.710 ;
        RECT 227.795 44.120 228.600 44.540 ;
        RECT 229.190 43.950 229.440 44.790 ;
        RECT 229.635 44.120 229.935 44.960 ;
        RECT 230.785 44.790 231.015 45.780 ;
        RECT 230.265 44.620 231.015 44.790 ;
        RECT 230.265 44.120 230.520 44.620 ;
        RECT 230.690 43.950 231.020 44.450 ;
        RECT 231.190 44.120 231.360 46.240 ;
        RECT 231.720 46.140 232.050 46.500 ;
        RECT 232.220 46.110 232.715 46.280 ;
        RECT 232.920 46.110 233.775 46.280 ;
        RECT 231.590 44.920 232.050 45.970 ;
        RECT 231.530 44.135 231.855 44.920 ;
        RECT 232.220 44.750 232.390 46.110 ;
        RECT 232.560 45.200 232.910 45.820 ;
        RECT 233.080 45.600 233.435 45.820 ;
        RECT 233.080 45.010 233.250 45.600 ;
        RECT 233.605 45.400 233.775 46.110 ;
        RECT 234.650 46.040 234.980 46.500 ;
        RECT 235.190 46.140 235.540 46.310 ;
        RECT 233.980 45.570 234.770 45.820 ;
        RECT 235.190 45.750 235.450 46.140 ;
        RECT 235.760 46.050 236.710 46.330 ;
        RECT 236.880 46.060 237.070 46.500 ;
        RECT 237.240 46.120 238.310 46.290 ;
        RECT 234.940 45.400 235.110 45.580 ;
        RECT 232.220 44.580 232.615 44.750 ;
        RECT 232.785 44.620 233.250 45.010 ;
        RECT 233.420 45.230 235.110 45.400 ;
        RECT 232.445 44.450 232.615 44.580 ;
        RECT 233.420 44.450 233.590 45.230 ;
        RECT 235.280 45.060 235.450 45.750 ;
        RECT 233.950 44.890 235.450 45.060 ;
        RECT 235.640 45.090 235.850 45.880 ;
        RECT 236.020 45.260 236.370 45.880 ;
        RECT 236.540 45.270 236.710 46.050 ;
        RECT 237.240 45.890 237.410 46.120 ;
        RECT 236.880 45.720 237.410 45.890 ;
        RECT 236.880 45.440 237.100 45.720 ;
        RECT 237.580 45.550 237.820 45.950 ;
        RECT 236.540 45.100 236.945 45.270 ;
        RECT 237.280 45.180 237.820 45.550 ;
        RECT 237.990 45.765 238.310 46.120 ;
        RECT 238.555 46.040 238.860 46.500 ;
        RECT 239.030 45.790 239.285 46.320 ;
        RECT 237.990 45.590 238.315 45.765 ;
        RECT 237.990 45.290 238.905 45.590 ;
        RECT 238.165 45.260 238.905 45.290 ;
        RECT 235.640 44.930 236.315 45.090 ;
        RECT 236.775 45.010 236.945 45.100 ;
        RECT 235.640 44.920 236.605 44.930 ;
        RECT 235.280 44.750 235.450 44.890 ;
        RECT 232.025 43.950 232.275 44.410 ;
        RECT 232.445 44.120 232.695 44.450 ;
        RECT 232.910 44.120 233.590 44.450 ;
        RECT 233.760 44.550 234.835 44.720 ;
        RECT 235.280 44.580 235.840 44.750 ;
        RECT 236.145 44.630 236.605 44.920 ;
        RECT 236.775 44.840 237.995 45.010 ;
        RECT 233.760 44.210 233.930 44.550 ;
        RECT 234.165 43.950 234.495 44.380 ;
        RECT 234.665 44.210 234.835 44.550 ;
        RECT 235.130 43.950 235.500 44.410 ;
        RECT 235.670 44.120 235.840 44.580 ;
        RECT 236.775 44.460 236.945 44.840 ;
        RECT 238.165 44.670 238.335 45.260 ;
        RECT 239.075 45.140 239.285 45.790 ;
        RECT 239.460 45.775 239.750 46.500 ;
        RECT 240.080 45.940 240.410 46.330 ;
        RECT 240.580 46.110 241.765 46.280 ;
        RECT 242.025 46.030 242.195 46.500 ;
        RECT 240.080 45.760 240.590 45.940 ;
        RECT 239.920 45.300 240.250 45.590 ;
        RECT 236.075 44.120 236.945 44.460 ;
        RECT 237.535 44.500 238.335 44.670 ;
        RECT 237.115 43.950 237.365 44.410 ;
        RECT 237.535 44.210 237.705 44.500 ;
        RECT 237.885 43.950 238.215 44.330 ;
        RECT 238.555 43.950 238.860 45.090 ;
        RECT 239.030 44.260 239.285 45.140 ;
        RECT 240.420 45.130 240.590 45.760 ;
        RECT 240.995 45.850 241.380 45.940 ;
        RECT 242.365 45.850 242.695 46.315 ;
        RECT 240.995 45.680 242.695 45.850 ;
        RECT 242.865 45.680 243.035 46.500 ;
        RECT 243.205 45.680 243.890 46.320 ;
        RECT 240.760 45.300 241.090 45.510 ;
        RECT 241.270 45.260 241.650 45.510 ;
        RECT 239.460 43.950 239.750 45.115 ;
        RECT 240.075 44.960 241.160 45.130 ;
        RECT 240.075 44.120 240.375 44.960 ;
        RECT 240.570 43.950 240.820 44.790 ;
        RECT 240.990 44.710 241.160 44.960 ;
        RECT 241.330 44.880 241.650 45.260 ;
        RECT 241.840 45.300 242.325 45.510 ;
        RECT 242.515 45.300 242.965 45.510 ;
        RECT 243.135 45.300 243.470 45.510 ;
        RECT 241.840 45.140 242.215 45.300 ;
        RECT 241.820 44.970 242.215 45.140 ;
        RECT 243.135 45.130 243.305 45.300 ;
        RECT 241.840 44.880 242.215 44.970 ;
        RECT 242.385 44.960 243.305 45.130 ;
        RECT 242.385 44.710 242.555 44.960 ;
        RECT 240.990 44.540 242.555 44.710 ;
        RECT 241.410 44.120 242.215 44.540 ;
        RECT 242.725 43.950 243.055 44.790 ;
        RECT 243.640 44.710 243.890 45.680 ;
        RECT 243.225 44.120 243.890 44.710 ;
        RECT 244.060 45.760 244.445 46.330 ;
        RECT 244.615 46.040 244.940 46.500 ;
        RECT 245.460 45.870 245.740 46.330 ;
        RECT 244.060 45.090 244.340 45.760 ;
        RECT 244.615 45.700 245.740 45.870 ;
        RECT 244.615 45.590 245.065 45.700 ;
        RECT 244.510 45.260 245.065 45.590 ;
        RECT 245.930 45.530 246.330 46.330 ;
        RECT 246.730 46.040 247.000 46.500 ;
        RECT 247.170 45.870 247.455 46.330 ;
        RECT 244.060 44.120 244.445 45.090 ;
        RECT 244.615 44.800 245.065 45.260 ;
        RECT 245.235 44.970 246.330 45.530 ;
        RECT 244.615 44.580 245.740 44.800 ;
        RECT 244.615 43.950 244.940 44.410 ;
        RECT 245.460 44.120 245.740 44.580 ;
        RECT 245.930 44.120 246.330 44.970 ;
        RECT 246.500 45.700 247.455 45.870 ;
        RECT 248.205 45.950 248.460 46.240 ;
        RECT 248.630 46.120 248.960 46.500 ;
        RECT 248.205 45.780 248.955 45.950 ;
        RECT 246.500 44.800 246.710 45.700 ;
        RECT 246.880 44.970 247.570 45.530 ;
        RECT 248.205 44.960 248.555 45.610 ;
        RECT 246.500 44.580 247.455 44.800 ;
        RECT 248.725 44.790 248.955 45.780 ;
        RECT 246.730 43.950 247.000 44.410 ;
        RECT 247.170 44.120 247.455 44.580 ;
        RECT 248.205 44.620 248.955 44.790 ;
        RECT 248.205 44.120 248.460 44.620 ;
        RECT 248.630 43.950 248.960 44.450 ;
        RECT 249.130 44.120 249.300 46.240 ;
        RECT 249.660 46.140 249.990 46.500 ;
        RECT 250.160 46.110 250.655 46.280 ;
        RECT 250.860 46.110 251.715 46.280 ;
        RECT 249.530 44.920 249.990 45.970 ;
        RECT 249.470 44.135 249.795 44.920 ;
        RECT 250.160 44.750 250.330 46.110 ;
        RECT 250.500 45.200 250.850 45.820 ;
        RECT 251.020 45.600 251.375 45.820 ;
        RECT 251.020 45.010 251.190 45.600 ;
        RECT 251.545 45.400 251.715 46.110 ;
        RECT 252.590 46.040 252.920 46.500 ;
        RECT 253.130 46.140 253.480 46.310 ;
        RECT 251.920 45.570 252.710 45.820 ;
        RECT 253.130 45.750 253.390 46.140 ;
        RECT 253.700 46.050 254.650 46.330 ;
        RECT 254.820 46.060 255.010 46.500 ;
        RECT 255.180 46.120 256.250 46.290 ;
        RECT 252.880 45.400 253.050 45.580 ;
        RECT 250.160 44.580 250.555 44.750 ;
        RECT 250.725 44.620 251.190 45.010 ;
        RECT 251.360 45.230 253.050 45.400 ;
        RECT 250.385 44.450 250.555 44.580 ;
        RECT 251.360 44.450 251.530 45.230 ;
        RECT 253.220 45.060 253.390 45.750 ;
        RECT 251.890 44.890 253.390 45.060 ;
        RECT 253.580 45.090 253.790 45.880 ;
        RECT 253.960 45.260 254.310 45.880 ;
        RECT 254.480 45.270 254.650 46.050 ;
        RECT 255.180 45.890 255.350 46.120 ;
        RECT 254.820 45.720 255.350 45.890 ;
        RECT 254.820 45.440 255.040 45.720 ;
        RECT 255.520 45.550 255.760 45.950 ;
        RECT 254.480 45.100 254.885 45.270 ;
        RECT 255.220 45.180 255.760 45.550 ;
        RECT 255.930 45.765 256.250 46.120 ;
        RECT 256.495 46.040 256.800 46.500 ;
        RECT 256.970 45.790 257.225 46.320 ;
        RECT 255.930 45.590 256.255 45.765 ;
        RECT 255.930 45.290 256.845 45.590 ;
        RECT 256.105 45.260 256.845 45.290 ;
        RECT 253.580 44.930 254.255 45.090 ;
        RECT 254.715 45.010 254.885 45.100 ;
        RECT 253.580 44.920 254.545 44.930 ;
        RECT 253.220 44.750 253.390 44.890 ;
        RECT 249.965 43.950 250.215 44.410 ;
        RECT 250.385 44.120 250.635 44.450 ;
        RECT 250.850 44.120 251.530 44.450 ;
        RECT 251.700 44.550 252.775 44.720 ;
        RECT 253.220 44.580 253.780 44.750 ;
        RECT 254.085 44.630 254.545 44.920 ;
        RECT 254.715 44.840 255.935 45.010 ;
        RECT 251.700 44.210 251.870 44.550 ;
        RECT 252.105 43.950 252.435 44.380 ;
        RECT 252.605 44.210 252.775 44.550 ;
        RECT 253.070 43.950 253.440 44.410 ;
        RECT 253.610 44.120 253.780 44.580 ;
        RECT 254.715 44.460 254.885 44.840 ;
        RECT 256.105 44.670 256.275 45.260 ;
        RECT 257.015 45.140 257.225 45.790 ;
        RECT 254.015 44.120 254.885 44.460 ;
        RECT 255.475 44.500 256.275 44.670 ;
        RECT 255.055 43.950 255.305 44.410 ;
        RECT 255.475 44.210 255.645 44.500 ;
        RECT 255.825 43.950 256.155 44.330 ;
        RECT 256.495 43.950 256.800 45.090 ;
        RECT 256.970 44.260 257.225 45.140 ;
        RECT 257.400 45.760 257.785 46.330 ;
        RECT 257.955 46.040 258.280 46.500 ;
        RECT 258.800 45.870 259.080 46.330 ;
        RECT 257.400 45.090 257.680 45.760 ;
        RECT 257.955 45.700 259.080 45.870 ;
        RECT 257.955 45.590 258.405 45.700 ;
        RECT 257.850 45.260 258.405 45.590 ;
        RECT 259.270 45.530 259.670 46.330 ;
        RECT 260.070 46.040 260.340 46.500 ;
        RECT 260.510 45.870 260.795 46.330 ;
        RECT 257.400 44.120 257.785 45.090 ;
        RECT 257.955 44.800 258.405 45.260 ;
        RECT 258.575 44.970 259.670 45.530 ;
        RECT 257.955 44.580 259.080 44.800 ;
        RECT 257.955 43.950 258.280 44.410 ;
        RECT 258.800 44.120 259.080 44.580 ;
        RECT 259.270 44.120 259.670 44.970 ;
        RECT 259.840 45.700 260.795 45.870 ;
        RECT 261.080 46.000 261.340 46.330 ;
        RECT 261.510 46.140 261.840 46.500 ;
        RECT 262.095 46.120 263.395 46.330 ;
        RECT 259.840 44.800 260.050 45.700 ;
        RECT 260.220 44.970 260.910 45.530 ;
        RECT 261.080 44.800 261.250 46.000 ;
        RECT 262.095 45.970 262.265 46.120 ;
        RECT 261.510 45.845 262.265 45.970 ;
        RECT 261.420 45.800 262.265 45.845 ;
        RECT 261.420 45.680 261.690 45.800 ;
        RECT 261.420 45.105 261.590 45.680 ;
        RECT 261.820 45.240 262.230 45.545 ;
        RECT 262.520 45.510 262.730 45.910 ;
        RECT 262.400 45.300 262.730 45.510 ;
        RECT 262.975 45.510 263.195 45.910 ;
        RECT 263.670 45.735 264.125 46.500 ;
        RECT 265.220 45.775 265.510 46.500 ;
        RECT 265.680 46.120 266.570 46.290 ;
        RECT 265.680 45.565 266.230 45.950 ;
        RECT 262.975 45.300 263.450 45.510 ;
        RECT 263.640 45.310 264.130 45.510 ;
        RECT 266.400 45.395 266.570 46.120 ;
        RECT 265.680 45.325 266.570 45.395 ;
        RECT 266.740 45.795 266.960 46.280 ;
        RECT 267.130 45.960 267.380 46.500 ;
        RECT 267.550 45.850 267.810 46.330 ;
        RECT 268.005 46.100 268.335 46.500 ;
        RECT 268.505 45.930 268.675 46.200 ;
        RECT 268.845 45.990 269.160 46.500 ;
        RECT 269.390 45.990 269.680 46.330 ;
        RECT 269.850 45.990 270.090 46.500 ;
        RECT 270.390 46.120 271.560 46.330 ;
        RECT 270.390 46.100 270.720 46.120 ;
        RECT 266.740 45.370 267.070 45.795 ;
        RECT 265.680 45.300 266.575 45.325 ;
        RECT 265.680 45.285 266.585 45.300 ;
        RECT 265.680 45.270 266.590 45.285 ;
        RECT 265.680 45.265 266.600 45.270 ;
        RECT 265.680 45.255 266.605 45.265 ;
        RECT 265.680 45.245 266.610 45.255 ;
        RECT 265.680 45.240 266.620 45.245 ;
        RECT 265.680 45.230 266.630 45.240 ;
        RECT 265.680 45.225 266.640 45.230 ;
        RECT 261.420 45.070 261.620 45.105 ;
        RECT 262.950 45.070 264.125 45.130 ;
        RECT 261.420 44.960 264.125 45.070 ;
        RECT 261.480 44.900 263.280 44.960 ;
        RECT 262.950 44.870 263.280 44.900 ;
        RECT 259.840 44.580 260.795 44.800 ;
        RECT 260.070 43.950 260.340 44.410 ;
        RECT 260.510 44.120 260.795 44.580 ;
        RECT 261.080 44.120 261.340 44.800 ;
        RECT 261.510 43.950 261.760 44.730 ;
        RECT 262.010 44.700 262.845 44.710 ;
        RECT 263.435 44.700 263.620 44.790 ;
        RECT 262.010 44.500 263.620 44.700 ;
        RECT 262.010 44.120 262.260 44.500 ;
        RECT 263.390 44.460 263.620 44.500 ;
        RECT 263.870 44.340 264.125 44.960 ;
        RECT 262.430 43.950 262.785 44.330 ;
        RECT 263.790 44.120 264.125 44.340 ;
        RECT 265.220 43.950 265.510 45.115 ;
        RECT 265.680 44.775 265.940 45.225 ;
        RECT 266.305 45.220 266.640 45.225 ;
        RECT 266.305 45.215 266.655 45.220 ;
        RECT 266.305 45.205 266.670 45.215 ;
        RECT 266.305 45.200 266.695 45.205 ;
        RECT 267.240 45.200 267.470 45.595 ;
        RECT 266.305 45.195 267.470 45.200 ;
        RECT 266.335 45.160 267.470 45.195 ;
        RECT 266.370 45.135 267.470 45.160 ;
        RECT 266.400 45.105 267.470 45.135 ;
        RECT 266.420 45.075 267.470 45.105 ;
        RECT 266.440 45.045 267.470 45.075 ;
        RECT 266.510 45.035 267.470 45.045 ;
        RECT 266.535 45.025 267.470 45.035 ;
        RECT 266.555 45.010 267.470 45.025 ;
        RECT 266.575 44.995 267.470 45.010 ;
        RECT 266.580 44.985 267.365 44.995 ;
        RECT 266.595 44.950 267.365 44.985 ;
        RECT 266.110 44.630 266.440 44.875 ;
        RECT 266.610 44.700 267.365 44.950 ;
        RECT 267.640 44.820 267.810 45.850 ;
        RECT 266.110 44.605 266.295 44.630 ;
        RECT 265.680 44.505 266.295 44.605 ;
        RECT 265.680 43.950 266.285 44.505 ;
        RECT 266.460 44.120 266.940 44.460 ;
        RECT 267.110 43.950 267.365 44.495 ;
        RECT 267.535 44.120 267.810 44.820 ;
        RECT 267.980 45.760 268.675 45.930 ;
        RECT 267.980 44.750 268.410 45.760 ;
        RECT 268.580 45.090 268.750 45.590 ;
        RECT 268.920 45.260 269.330 45.820 ;
        RECT 269.500 45.090 269.680 45.990 ;
        RECT 269.850 45.480 270.045 45.820 ;
        RECT 270.280 45.680 271.140 45.930 ;
        RECT 271.310 45.870 271.560 46.120 ;
        RECT 271.730 46.040 271.900 46.500 ;
        RECT 272.070 45.870 272.410 46.330 ;
        RECT 272.580 45.955 277.925 46.500 ;
        RECT 271.310 45.700 272.410 45.870 ;
        RECT 269.850 45.310 270.050 45.480 ;
        RECT 269.850 45.260 270.045 45.310 ;
        RECT 270.280 45.090 270.560 45.680 ;
        RECT 270.730 45.260 271.480 45.510 ;
        RECT 271.650 45.260 272.410 45.510 ;
        RECT 274.165 45.125 274.505 45.955 ;
        RECT 278.835 45.690 279.080 46.295 ;
        RECT 279.300 45.965 279.810 46.500 ;
        RECT 268.580 44.920 270.040 45.090 ;
        RECT 270.280 44.920 271.980 45.090 ;
        RECT 267.980 44.580 268.755 44.750 ;
        RECT 268.085 43.950 268.255 44.410 ;
        RECT 268.425 44.120 268.755 44.580 ;
        RECT 268.925 43.950 269.095 44.750 ;
        RECT 269.680 44.745 270.040 44.920 ;
        RECT 270.385 43.950 270.640 44.750 ;
        RECT 270.810 44.120 271.140 44.920 ;
        RECT 271.310 43.950 271.480 44.750 ;
        RECT 271.650 44.120 271.980 44.920 ;
        RECT 272.150 43.950 272.410 45.090 ;
        RECT 275.985 44.385 276.335 45.635 ;
        RECT 278.560 45.520 279.790 45.690 ;
        RECT 278.560 44.710 278.900 45.520 ;
        RECT 279.070 44.955 279.820 45.145 ;
        RECT 272.580 43.950 277.925 44.385 ;
        RECT 278.560 44.300 279.075 44.710 ;
        RECT 279.310 43.950 279.480 44.710 ;
        RECT 279.650 44.290 279.820 44.955 ;
        RECT 279.990 44.970 280.180 46.330 ;
        RECT 280.350 46.160 280.625 46.330 ;
        RECT 280.350 45.990 280.630 46.160 ;
        RECT 280.350 45.170 280.625 45.990 ;
        RECT 280.815 45.965 281.345 46.330 ;
        RECT 281.770 46.100 282.100 46.500 ;
        RECT 281.170 45.930 281.345 45.965 ;
        RECT 280.830 44.970 281.000 45.770 ;
        RECT 279.990 44.800 281.000 44.970 ;
        RECT 281.170 45.760 282.100 45.930 ;
        RECT 282.270 45.760 282.525 46.330 ;
        RECT 281.170 44.630 281.340 45.760 ;
        RECT 281.930 45.590 282.100 45.760 ;
        RECT 280.215 44.460 281.340 44.630 ;
        RECT 281.510 45.260 281.705 45.590 ;
        RECT 281.930 45.260 282.185 45.590 ;
        RECT 281.510 44.290 281.680 45.260 ;
        RECT 282.355 45.090 282.525 45.760 ;
        RECT 282.815 45.870 283.100 46.330 ;
        RECT 283.270 46.040 283.540 46.500 ;
        RECT 282.815 45.700 283.770 45.870 ;
        RECT 279.650 44.120 281.680 44.290 ;
        RECT 281.850 43.950 282.020 45.090 ;
        RECT 282.190 44.120 282.525 45.090 ;
        RECT 282.700 44.970 283.390 45.530 ;
        RECT 283.560 44.800 283.770 45.700 ;
        RECT 282.815 44.580 283.770 44.800 ;
        RECT 283.940 45.530 284.340 46.330 ;
        RECT 284.530 45.870 284.810 46.330 ;
        RECT 285.330 46.040 285.655 46.500 ;
        RECT 284.530 45.700 285.655 45.870 ;
        RECT 285.825 45.760 286.210 46.330 ;
        RECT 285.205 45.590 285.655 45.700 ;
        RECT 283.940 44.970 285.035 45.530 ;
        RECT 285.205 45.260 285.760 45.590 ;
        RECT 282.815 44.120 283.100 44.580 ;
        RECT 283.270 43.950 283.540 44.410 ;
        RECT 283.940 44.120 284.340 44.970 ;
        RECT 285.205 44.800 285.655 45.260 ;
        RECT 285.930 45.090 286.210 45.760 ;
        RECT 286.380 45.730 289.890 46.500 ;
        RECT 290.980 45.775 291.270 46.500 ;
        RECT 291.445 45.790 291.700 46.320 ;
        RECT 291.870 46.040 292.175 46.500 ;
        RECT 292.420 46.120 293.490 46.290 ;
        RECT 286.380 45.210 288.030 45.730 ;
        RECT 284.530 44.580 285.655 44.800 ;
        RECT 284.530 44.120 284.810 44.580 ;
        RECT 285.330 43.950 285.655 44.410 ;
        RECT 285.825 44.120 286.210 45.090 ;
        RECT 288.200 45.040 289.890 45.560 ;
        RECT 291.445 45.140 291.655 45.790 ;
        RECT 292.420 45.765 292.740 46.120 ;
        RECT 292.415 45.590 292.740 45.765 ;
        RECT 291.825 45.290 292.740 45.590 ;
        RECT 292.910 45.550 293.150 45.950 ;
        RECT 293.320 45.890 293.490 46.120 ;
        RECT 293.660 46.060 293.850 46.500 ;
        RECT 294.020 46.050 294.970 46.330 ;
        RECT 295.190 46.140 295.540 46.310 ;
        RECT 293.320 45.720 293.850 45.890 ;
        RECT 291.825 45.260 292.565 45.290 ;
        RECT 286.380 43.950 289.890 45.040 ;
        RECT 290.980 43.950 291.270 45.115 ;
        RECT 291.445 44.260 291.700 45.140 ;
        RECT 291.870 43.950 292.175 45.090 ;
        RECT 292.395 44.670 292.565 45.260 ;
        RECT 292.910 45.180 293.450 45.550 ;
        RECT 293.630 45.440 293.850 45.720 ;
        RECT 294.020 45.270 294.190 46.050 ;
        RECT 293.785 45.100 294.190 45.270 ;
        RECT 294.360 45.260 294.710 45.880 ;
        RECT 293.785 45.010 293.955 45.100 ;
        RECT 294.880 45.090 295.090 45.880 ;
        RECT 292.735 44.840 293.955 45.010 ;
        RECT 294.415 44.930 295.090 45.090 ;
        RECT 292.395 44.500 293.195 44.670 ;
        RECT 292.515 43.950 292.845 44.330 ;
        RECT 293.025 44.210 293.195 44.500 ;
        RECT 293.785 44.460 293.955 44.840 ;
        RECT 294.125 44.920 295.090 44.930 ;
        RECT 295.280 45.750 295.540 46.140 ;
        RECT 295.750 46.040 296.080 46.500 ;
        RECT 296.955 46.110 297.810 46.280 ;
        RECT 298.015 46.110 298.510 46.280 ;
        RECT 298.680 46.140 299.010 46.500 ;
        RECT 295.280 45.060 295.450 45.750 ;
        RECT 295.620 45.400 295.790 45.580 ;
        RECT 295.960 45.570 296.750 45.820 ;
        RECT 296.955 45.400 297.125 46.110 ;
        RECT 297.295 45.600 297.650 45.820 ;
        RECT 295.620 45.230 297.310 45.400 ;
        RECT 294.125 44.630 294.585 44.920 ;
        RECT 295.280 44.890 296.780 45.060 ;
        RECT 295.280 44.750 295.450 44.890 ;
        RECT 294.890 44.580 295.450 44.750 ;
        RECT 293.365 43.950 293.615 44.410 ;
        RECT 293.785 44.120 294.655 44.460 ;
        RECT 294.890 44.120 295.060 44.580 ;
        RECT 295.895 44.550 296.970 44.720 ;
        RECT 295.230 43.950 295.600 44.410 ;
        RECT 295.895 44.210 296.065 44.550 ;
        RECT 296.235 43.950 296.565 44.380 ;
        RECT 296.800 44.210 296.970 44.550 ;
        RECT 297.140 44.450 297.310 45.230 ;
        RECT 297.480 45.010 297.650 45.600 ;
        RECT 297.820 45.200 298.170 45.820 ;
        RECT 297.480 44.620 297.945 45.010 ;
        RECT 298.340 44.750 298.510 46.110 ;
        RECT 298.680 44.920 299.140 45.970 ;
        RECT 298.115 44.580 298.510 44.750 ;
        RECT 298.115 44.450 298.285 44.580 ;
        RECT 297.140 44.120 297.820 44.450 ;
        RECT 298.035 44.120 298.285 44.450 ;
        RECT 298.455 43.950 298.705 44.410 ;
        RECT 298.875 44.135 299.200 44.920 ;
        RECT 299.370 44.120 299.540 46.240 ;
        RECT 299.710 46.120 300.040 46.500 ;
        RECT 300.210 45.950 300.465 46.240 ;
        RECT 300.640 45.955 305.985 46.500 ;
        RECT 299.715 45.780 300.465 45.950 ;
        RECT 299.715 44.790 299.945 45.780 ;
        RECT 300.115 44.960 300.465 45.610 ;
        RECT 302.225 45.125 302.565 45.955 ;
        RECT 306.160 45.730 309.670 46.500 ;
        RECT 309.840 45.750 311.050 46.500 ;
        RECT 299.715 44.620 300.465 44.790 ;
        RECT 299.710 43.950 300.040 44.450 ;
        RECT 300.210 44.120 300.465 44.620 ;
        RECT 304.045 44.385 304.395 45.635 ;
        RECT 306.160 45.210 307.810 45.730 ;
        RECT 307.980 45.040 309.670 45.560 ;
        RECT 300.640 43.950 305.985 44.385 ;
        RECT 306.160 43.950 309.670 45.040 ;
        RECT 309.840 45.040 310.360 45.580 ;
        RECT 310.530 45.210 311.050 45.750 ;
        RECT 309.840 43.950 311.050 45.040 ;
        RECT 162.095 43.780 311.135 43.950 ;
        RECT 162.180 42.690 163.390 43.780 ;
        RECT 163.560 42.690 165.230 43.780 ;
        RECT 165.865 43.110 166.120 43.610 ;
        RECT 166.290 43.280 166.620 43.780 ;
        RECT 165.865 42.940 166.615 43.110 ;
        RECT 162.180 41.980 162.700 42.520 ;
        RECT 162.870 42.150 163.390 42.690 ;
        RECT 163.560 42.000 164.310 42.520 ;
        RECT 164.480 42.170 165.230 42.690 ;
        RECT 165.865 42.120 166.215 42.770 ;
        RECT 162.180 41.230 163.390 41.980 ;
        RECT 163.560 41.230 165.230 42.000 ;
        RECT 166.385 41.950 166.615 42.940 ;
        RECT 165.865 41.780 166.615 41.950 ;
        RECT 165.865 41.490 166.120 41.780 ;
        RECT 166.290 41.230 166.620 41.610 ;
        RECT 166.790 41.490 166.960 43.610 ;
        RECT 167.130 42.810 167.455 43.595 ;
        RECT 167.625 43.320 167.875 43.780 ;
        RECT 168.045 43.280 168.295 43.610 ;
        RECT 168.510 43.280 169.190 43.610 ;
        RECT 168.045 43.150 168.215 43.280 ;
        RECT 167.820 42.980 168.215 43.150 ;
        RECT 167.190 41.760 167.650 42.810 ;
        RECT 167.820 41.620 167.990 42.980 ;
        RECT 168.385 42.720 168.850 43.110 ;
        RECT 168.160 41.910 168.510 42.530 ;
        RECT 168.680 42.130 168.850 42.720 ;
        RECT 169.020 42.500 169.190 43.280 ;
        RECT 169.360 43.180 169.530 43.520 ;
        RECT 169.765 43.350 170.095 43.780 ;
        RECT 170.265 43.180 170.435 43.520 ;
        RECT 170.730 43.320 171.100 43.780 ;
        RECT 169.360 43.010 170.435 43.180 ;
        RECT 171.270 43.150 171.440 43.610 ;
        RECT 171.675 43.270 172.545 43.610 ;
        RECT 172.715 43.320 172.965 43.780 ;
        RECT 170.880 42.980 171.440 43.150 ;
        RECT 170.880 42.840 171.050 42.980 ;
        RECT 169.550 42.670 171.050 42.840 ;
        RECT 171.745 42.810 172.205 43.100 ;
        RECT 169.020 42.330 170.710 42.500 ;
        RECT 168.680 41.910 169.035 42.130 ;
        RECT 169.205 41.620 169.375 42.330 ;
        RECT 169.580 41.910 170.370 42.160 ;
        RECT 170.540 42.150 170.710 42.330 ;
        RECT 170.880 41.980 171.050 42.670 ;
        RECT 167.320 41.230 167.650 41.590 ;
        RECT 167.820 41.450 168.315 41.620 ;
        RECT 168.520 41.450 169.375 41.620 ;
        RECT 170.250 41.230 170.580 41.690 ;
        RECT 170.790 41.590 171.050 41.980 ;
        RECT 171.240 42.800 172.205 42.810 ;
        RECT 172.375 42.890 172.545 43.270 ;
        RECT 173.135 43.230 173.305 43.520 ;
        RECT 173.485 43.400 173.815 43.780 ;
        RECT 173.135 43.060 173.935 43.230 ;
        RECT 171.240 42.640 171.915 42.800 ;
        RECT 172.375 42.720 173.595 42.890 ;
        RECT 171.240 41.850 171.450 42.640 ;
        RECT 172.375 42.630 172.545 42.720 ;
        RECT 171.620 41.850 171.970 42.470 ;
        RECT 172.140 42.460 172.545 42.630 ;
        RECT 172.140 41.680 172.310 42.460 ;
        RECT 172.480 42.010 172.700 42.290 ;
        RECT 172.880 42.180 173.420 42.550 ;
        RECT 173.765 42.470 173.935 43.060 ;
        RECT 174.155 42.640 174.460 43.780 ;
        RECT 174.630 42.590 174.885 43.470 ;
        RECT 175.060 42.615 175.350 43.780 ;
        RECT 175.525 43.110 175.780 43.610 ;
        RECT 175.950 43.280 176.280 43.780 ;
        RECT 175.525 42.940 176.275 43.110 ;
        RECT 173.765 42.440 174.505 42.470 ;
        RECT 172.480 41.840 173.010 42.010 ;
        RECT 170.790 41.420 171.140 41.590 ;
        RECT 171.360 41.400 172.310 41.680 ;
        RECT 172.480 41.230 172.670 41.670 ;
        RECT 172.840 41.610 173.010 41.840 ;
        RECT 173.180 41.780 173.420 42.180 ;
        RECT 173.590 42.140 174.505 42.440 ;
        RECT 173.590 41.965 173.915 42.140 ;
        RECT 173.590 41.610 173.910 41.965 ;
        RECT 174.675 41.940 174.885 42.590 ;
        RECT 175.525 42.120 175.875 42.770 ;
        RECT 172.840 41.440 173.910 41.610 ;
        RECT 174.155 41.230 174.460 41.690 ;
        RECT 174.630 41.410 174.885 41.940 ;
        RECT 175.060 41.230 175.350 41.955 ;
        RECT 176.045 41.950 176.275 42.940 ;
        RECT 175.525 41.780 176.275 41.950 ;
        RECT 175.525 41.490 175.780 41.780 ;
        RECT 175.950 41.230 176.280 41.610 ;
        RECT 176.450 41.490 176.620 43.610 ;
        RECT 176.790 42.810 177.115 43.595 ;
        RECT 177.285 43.320 177.535 43.780 ;
        RECT 177.705 43.280 177.955 43.610 ;
        RECT 178.170 43.280 178.850 43.610 ;
        RECT 177.705 43.150 177.875 43.280 ;
        RECT 177.480 42.980 177.875 43.150 ;
        RECT 176.850 41.760 177.310 42.810 ;
        RECT 177.480 41.620 177.650 42.980 ;
        RECT 178.045 42.720 178.510 43.110 ;
        RECT 177.820 41.910 178.170 42.530 ;
        RECT 178.340 42.130 178.510 42.720 ;
        RECT 178.680 42.500 178.850 43.280 ;
        RECT 179.020 43.180 179.190 43.520 ;
        RECT 179.425 43.350 179.755 43.780 ;
        RECT 179.925 43.180 180.095 43.520 ;
        RECT 180.390 43.320 180.760 43.780 ;
        RECT 179.020 43.010 180.095 43.180 ;
        RECT 180.930 43.150 181.100 43.610 ;
        RECT 181.335 43.270 182.205 43.610 ;
        RECT 182.375 43.320 182.625 43.780 ;
        RECT 180.540 42.980 181.100 43.150 ;
        RECT 180.540 42.840 180.710 42.980 ;
        RECT 179.210 42.670 180.710 42.840 ;
        RECT 181.405 42.810 181.865 43.100 ;
        RECT 178.680 42.330 180.370 42.500 ;
        RECT 178.340 41.910 178.695 42.130 ;
        RECT 178.865 41.620 179.035 42.330 ;
        RECT 179.240 41.910 180.030 42.160 ;
        RECT 180.200 42.150 180.370 42.330 ;
        RECT 180.540 41.980 180.710 42.670 ;
        RECT 176.980 41.230 177.310 41.590 ;
        RECT 177.480 41.450 177.975 41.620 ;
        RECT 178.180 41.450 179.035 41.620 ;
        RECT 179.910 41.230 180.240 41.690 ;
        RECT 180.450 41.590 180.710 41.980 ;
        RECT 180.900 42.800 181.865 42.810 ;
        RECT 182.035 42.890 182.205 43.270 ;
        RECT 182.795 43.230 182.965 43.520 ;
        RECT 183.145 43.400 183.475 43.780 ;
        RECT 182.795 43.060 183.595 43.230 ;
        RECT 180.900 42.640 181.575 42.800 ;
        RECT 182.035 42.720 183.255 42.890 ;
        RECT 180.900 41.850 181.110 42.640 ;
        RECT 182.035 42.630 182.205 42.720 ;
        RECT 181.280 41.850 181.630 42.470 ;
        RECT 181.800 42.460 182.205 42.630 ;
        RECT 181.800 41.680 181.970 42.460 ;
        RECT 182.140 42.010 182.360 42.290 ;
        RECT 182.540 42.180 183.080 42.550 ;
        RECT 183.425 42.470 183.595 43.060 ;
        RECT 183.815 42.640 184.120 43.780 ;
        RECT 184.290 42.590 184.545 43.470 ;
        RECT 184.725 43.110 184.980 43.610 ;
        RECT 185.150 43.280 185.480 43.780 ;
        RECT 184.725 42.940 185.475 43.110 ;
        RECT 183.425 42.440 184.165 42.470 ;
        RECT 182.140 41.840 182.670 42.010 ;
        RECT 180.450 41.420 180.800 41.590 ;
        RECT 181.020 41.400 181.970 41.680 ;
        RECT 182.140 41.230 182.330 41.670 ;
        RECT 182.500 41.610 182.670 41.840 ;
        RECT 182.840 41.780 183.080 42.180 ;
        RECT 183.250 42.140 184.165 42.440 ;
        RECT 183.250 41.965 183.575 42.140 ;
        RECT 183.250 41.610 183.570 41.965 ;
        RECT 184.335 41.940 184.545 42.590 ;
        RECT 184.725 42.120 185.075 42.770 ;
        RECT 185.245 41.950 185.475 42.940 ;
        RECT 182.500 41.440 183.570 41.610 ;
        RECT 183.815 41.230 184.120 41.690 ;
        RECT 184.290 41.410 184.545 41.940 ;
        RECT 184.725 41.780 185.475 41.950 ;
        RECT 184.725 41.490 184.980 41.780 ;
        RECT 185.150 41.230 185.480 41.610 ;
        RECT 185.650 41.490 185.820 43.610 ;
        RECT 185.990 42.810 186.315 43.595 ;
        RECT 186.485 43.320 186.735 43.780 ;
        RECT 186.905 43.280 187.155 43.610 ;
        RECT 187.370 43.280 188.050 43.610 ;
        RECT 186.905 43.150 187.075 43.280 ;
        RECT 186.680 42.980 187.075 43.150 ;
        RECT 186.050 41.760 186.510 42.810 ;
        RECT 186.680 41.620 186.850 42.980 ;
        RECT 187.245 42.720 187.710 43.110 ;
        RECT 187.020 41.910 187.370 42.530 ;
        RECT 187.540 42.130 187.710 42.720 ;
        RECT 187.880 42.500 188.050 43.280 ;
        RECT 188.220 43.180 188.390 43.520 ;
        RECT 188.625 43.350 188.955 43.780 ;
        RECT 189.125 43.180 189.295 43.520 ;
        RECT 189.590 43.320 189.960 43.780 ;
        RECT 188.220 43.010 189.295 43.180 ;
        RECT 190.130 43.150 190.300 43.610 ;
        RECT 190.535 43.270 191.405 43.610 ;
        RECT 191.575 43.320 191.825 43.780 ;
        RECT 189.740 42.980 190.300 43.150 ;
        RECT 189.740 42.840 189.910 42.980 ;
        RECT 188.410 42.670 189.910 42.840 ;
        RECT 190.605 42.810 191.065 43.100 ;
        RECT 187.880 42.330 189.570 42.500 ;
        RECT 187.540 41.910 187.895 42.130 ;
        RECT 188.065 41.620 188.235 42.330 ;
        RECT 188.440 41.910 189.230 42.160 ;
        RECT 189.400 42.150 189.570 42.330 ;
        RECT 189.740 41.980 189.910 42.670 ;
        RECT 186.180 41.230 186.510 41.590 ;
        RECT 186.680 41.450 187.175 41.620 ;
        RECT 187.380 41.450 188.235 41.620 ;
        RECT 189.110 41.230 189.440 41.690 ;
        RECT 189.650 41.590 189.910 41.980 ;
        RECT 190.100 42.800 191.065 42.810 ;
        RECT 191.235 42.890 191.405 43.270 ;
        RECT 191.995 43.230 192.165 43.520 ;
        RECT 192.345 43.400 192.675 43.780 ;
        RECT 191.995 43.060 192.795 43.230 ;
        RECT 190.100 42.640 190.775 42.800 ;
        RECT 191.235 42.720 192.455 42.890 ;
        RECT 190.100 41.850 190.310 42.640 ;
        RECT 191.235 42.630 191.405 42.720 ;
        RECT 190.480 41.850 190.830 42.470 ;
        RECT 191.000 42.460 191.405 42.630 ;
        RECT 191.000 41.680 191.170 42.460 ;
        RECT 191.340 42.010 191.560 42.290 ;
        RECT 191.740 42.180 192.280 42.550 ;
        RECT 192.625 42.470 192.795 43.060 ;
        RECT 193.015 42.640 193.320 43.780 ;
        RECT 193.490 42.590 193.740 43.470 ;
        RECT 193.910 42.640 194.160 43.780 ;
        RECT 194.385 42.640 194.720 43.610 ;
        RECT 194.890 42.640 195.060 43.780 ;
        RECT 195.230 43.440 197.260 43.610 ;
        RECT 192.625 42.440 193.365 42.470 ;
        RECT 191.340 41.840 191.870 42.010 ;
        RECT 189.650 41.420 190.000 41.590 ;
        RECT 190.220 41.400 191.170 41.680 ;
        RECT 191.340 41.230 191.530 41.670 ;
        RECT 191.700 41.610 191.870 41.840 ;
        RECT 192.040 41.780 192.280 42.180 ;
        RECT 192.450 42.140 193.365 42.440 ;
        RECT 192.450 41.965 192.775 42.140 ;
        RECT 192.450 41.610 192.770 41.965 ;
        RECT 193.535 41.940 193.740 42.590 ;
        RECT 191.700 41.440 192.770 41.610 ;
        RECT 193.015 41.230 193.320 41.690 ;
        RECT 193.490 41.410 193.740 41.940 ;
        RECT 193.910 41.230 194.160 41.985 ;
        RECT 194.385 41.970 194.555 42.640 ;
        RECT 195.230 42.470 195.400 43.440 ;
        RECT 194.725 42.140 194.980 42.470 ;
        RECT 195.205 42.140 195.400 42.470 ;
        RECT 195.570 43.100 196.695 43.270 ;
        RECT 194.810 41.970 194.980 42.140 ;
        RECT 195.570 41.970 195.740 43.100 ;
        RECT 194.385 41.400 194.640 41.970 ;
        RECT 194.810 41.800 195.740 41.970 ;
        RECT 195.910 42.760 196.920 42.930 ;
        RECT 195.910 41.960 196.080 42.760 ;
        RECT 195.565 41.765 195.740 41.800 ;
        RECT 194.810 41.230 195.140 41.630 ;
        RECT 195.565 41.400 196.095 41.765 ;
        RECT 196.285 41.740 196.560 42.560 ;
        RECT 196.280 41.570 196.560 41.740 ;
        RECT 196.285 41.400 196.560 41.570 ;
        RECT 196.730 41.400 196.920 42.760 ;
        RECT 197.090 42.775 197.260 43.440 ;
        RECT 197.430 43.020 197.600 43.780 ;
        RECT 197.835 43.020 198.350 43.430 ;
        RECT 197.090 42.585 197.840 42.775 ;
        RECT 198.010 42.210 198.350 43.020 ;
        RECT 198.520 42.690 200.190 43.780 ;
        RECT 197.120 42.040 198.350 42.210 ;
        RECT 197.100 41.230 197.610 41.765 ;
        RECT 197.830 41.435 198.075 42.040 ;
        RECT 198.520 42.000 199.270 42.520 ;
        RECT 199.440 42.170 200.190 42.690 ;
        RECT 200.820 42.615 201.110 43.780 ;
        RECT 201.285 43.110 201.540 43.610 ;
        RECT 201.710 43.280 202.040 43.780 ;
        RECT 201.285 42.940 202.035 43.110 ;
        RECT 201.285 42.120 201.635 42.770 ;
        RECT 198.520 41.230 200.190 42.000 ;
        RECT 200.820 41.230 201.110 41.955 ;
        RECT 201.805 41.950 202.035 42.940 ;
        RECT 201.285 41.780 202.035 41.950 ;
        RECT 201.285 41.490 201.540 41.780 ;
        RECT 201.710 41.230 202.040 41.610 ;
        RECT 202.210 41.490 202.380 43.610 ;
        RECT 202.550 42.810 202.875 43.595 ;
        RECT 203.045 43.320 203.295 43.780 ;
        RECT 203.465 43.280 203.715 43.610 ;
        RECT 203.930 43.280 204.610 43.610 ;
        RECT 203.465 43.150 203.635 43.280 ;
        RECT 203.240 42.980 203.635 43.150 ;
        RECT 202.610 41.760 203.070 42.810 ;
        RECT 203.240 41.620 203.410 42.980 ;
        RECT 203.805 42.720 204.270 43.110 ;
        RECT 203.580 41.910 203.930 42.530 ;
        RECT 204.100 42.130 204.270 42.720 ;
        RECT 204.440 42.500 204.610 43.280 ;
        RECT 204.780 43.180 204.950 43.520 ;
        RECT 205.185 43.350 205.515 43.780 ;
        RECT 205.685 43.180 205.855 43.520 ;
        RECT 206.150 43.320 206.520 43.780 ;
        RECT 204.780 43.010 205.855 43.180 ;
        RECT 206.690 43.150 206.860 43.610 ;
        RECT 207.095 43.270 207.965 43.610 ;
        RECT 208.135 43.320 208.385 43.780 ;
        RECT 206.300 42.980 206.860 43.150 ;
        RECT 206.300 42.840 206.470 42.980 ;
        RECT 204.970 42.670 206.470 42.840 ;
        RECT 207.165 42.810 207.625 43.100 ;
        RECT 204.440 42.330 206.130 42.500 ;
        RECT 204.100 41.910 204.455 42.130 ;
        RECT 204.625 41.620 204.795 42.330 ;
        RECT 205.000 41.910 205.790 42.160 ;
        RECT 205.960 42.150 206.130 42.330 ;
        RECT 206.300 41.980 206.470 42.670 ;
        RECT 202.740 41.230 203.070 41.590 ;
        RECT 203.240 41.450 203.735 41.620 ;
        RECT 203.940 41.450 204.795 41.620 ;
        RECT 205.670 41.230 206.000 41.690 ;
        RECT 206.210 41.590 206.470 41.980 ;
        RECT 206.660 42.800 207.625 42.810 ;
        RECT 207.795 42.890 207.965 43.270 ;
        RECT 208.555 43.230 208.725 43.520 ;
        RECT 208.905 43.400 209.235 43.780 ;
        RECT 208.555 43.060 209.355 43.230 ;
        RECT 206.660 42.640 207.335 42.800 ;
        RECT 207.795 42.720 209.015 42.890 ;
        RECT 206.660 41.850 206.870 42.640 ;
        RECT 207.795 42.630 207.965 42.720 ;
        RECT 207.040 41.850 207.390 42.470 ;
        RECT 207.560 42.460 207.965 42.630 ;
        RECT 207.560 41.680 207.730 42.460 ;
        RECT 207.900 42.010 208.120 42.290 ;
        RECT 208.300 42.180 208.840 42.550 ;
        RECT 209.185 42.470 209.355 43.060 ;
        RECT 209.575 42.640 209.880 43.780 ;
        RECT 210.050 42.590 210.305 43.470 ;
        RECT 210.570 43.160 210.740 43.590 ;
        RECT 210.910 43.330 211.240 43.780 ;
        RECT 210.570 42.930 211.250 43.160 ;
        RECT 209.185 42.440 209.925 42.470 ;
        RECT 207.900 41.840 208.430 42.010 ;
        RECT 206.210 41.420 206.560 41.590 ;
        RECT 206.780 41.400 207.730 41.680 ;
        RECT 207.900 41.230 208.090 41.670 ;
        RECT 208.260 41.610 208.430 41.840 ;
        RECT 208.600 41.780 208.840 42.180 ;
        RECT 209.010 42.140 209.925 42.440 ;
        RECT 209.010 41.965 209.335 42.140 ;
        RECT 209.010 41.610 209.330 41.965 ;
        RECT 210.095 41.940 210.305 42.590 ;
        RECT 210.545 42.080 210.845 42.760 ;
        RECT 208.260 41.440 209.330 41.610 ;
        RECT 209.575 41.230 209.880 41.690 ;
        RECT 210.050 41.410 210.305 41.940 ;
        RECT 210.540 41.910 210.845 42.080 ;
        RECT 211.015 42.280 211.250 42.930 ;
        RECT 211.440 42.620 211.725 43.565 ;
        RECT 211.905 43.310 212.590 43.780 ;
        RECT 211.900 42.790 212.595 43.100 ;
        RECT 212.770 42.725 213.075 43.510 ;
        RECT 213.260 42.825 213.530 43.780 ;
        RECT 213.705 43.110 213.960 43.610 ;
        RECT 214.130 43.280 214.460 43.780 ;
        RECT 213.705 42.940 214.455 43.110 ;
        RECT 211.440 42.470 212.300 42.620 ;
        RECT 211.440 42.450 212.730 42.470 ;
        RECT 211.015 41.950 211.570 42.280 ;
        RECT 211.740 42.090 212.730 42.450 ;
        RECT 211.015 41.800 211.230 41.950 ;
        RECT 210.490 41.230 210.820 41.735 ;
        RECT 210.990 41.425 211.230 41.800 ;
        RECT 211.740 41.755 211.910 42.090 ;
        RECT 212.900 41.920 213.075 42.725 ;
        RECT 213.705 42.120 214.055 42.770 ;
        RECT 214.225 41.950 214.455 42.940 ;
        RECT 211.510 41.560 211.910 41.755 ;
        RECT 211.510 41.415 211.680 41.560 ;
        RECT 212.270 41.230 212.670 41.725 ;
        RECT 212.840 41.400 213.075 41.920 ;
        RECT 213.260 41.230 213.530 41.865 ;
        RECT 213.705 41.780 214.455 41.950 ;
        RECT 213.705 41.490 213.960 41.780 ;
        RECT 214.130 41.230 214.460 41.610 ;
        RECT 214.630 41.490 214.800 43.610 ;
        RECT 214.970 42.810 215.295 43.595 ;
        RECT 215.465 43.320 215.715 43.780 ;
        RECT 215.885 43.280 216.135 43.610 ;
        RECT 216.350 43.280 217.030 43.610 ;
        RECT 215.885 43.150 216.055 43.280 ;
        RECT 215.660 42.980 216.055 43.150 ;
        RECT 215.030 41.760 215.490 42.810 ;
        RECT 215.660 41.620 215.830 42.980 ;
        RECT 216.225 42.720 216.690 43.110 ;
        RECT 216.000 41.910 216.350 42.530 ;
        RECT 216.520 42.130 216.690 42.720 ;
        RECT 216.860 42.500 217.030 43.280 ;
        RECT 217.200 43.180 217.370 43.520 ;
        RECT 217.605 43.350 217.935 43.780 ;
        RECT 218.105 43.180 218.275 43.520 ;
        RECT 218.570 43.320 218.940 43.780 ;
        RECT 217.200 43.010 218.275 43.180 ;
        RECT 219.110 43.150 219.280 43.610 ;
        RECT 219.515 43.270 220.385 43.610 ;
        RECT 220.555 43.320 220.805 43.780 ;
        RECT 218.720 42.980 219.280 43.150 ;
        RECT 218.720 42.840 218.890 42.980 ;
        RECT 217.390 42.670 218.890 42.840 ;
        RECT 219.585 42.810 220.045 43.100 ;
        RECT 216.860 42.330 218.550 42.500 ;
        RECT 216.520 41.910 216.875 42.130 ;
        RECT 217.045 41.620 217.215 42.330 ;
        RECT 217.420 41.910 218.210 42.160 ;
        RECT 218.380 42.150 218.550 42.330 ;
        RECT 218.720 41.980 218.890 42.670 ;
        RECT 215.160 41.230 215.490 41.590 ;
        RECT 215.660 41.450 216.155 41.620 ;
        RECT 216.360 41.450 217.215 41.620 ;
        RECT 218.090 41.230 218.420 41.690 ;
        RECT 218.630 41.590 218.890 41.980 ;
        RECT 219.080 42.800 220.045 42.810 ;
        RECT 220.215 42.890 220.385 43.270 ;
        RECT 220.975 43.230 221.145 43.520 ;
        RECT 221.325 43.400 221.655 43.780 ;
        RECT 220.975 43.060 221.775 43.230 ;
        RECT 219.080 42.640 219.755 42.800 ;
        RECT 220.215 42.720 221.435 42.890 ;
        RECT 219.080 41.850 219.290 42.640 ;
        RECT 220.215 42.630 220.385 42.720 ;
        RECT 219.460 41.850 219.810 42.470 ;
        RECT 219.980 42.460 220.385 42.630 ;
        RECT 219.980 41.680 220.150 42.460 ;
        RECT 220.320 42.010 220.540 42.290 ;
        RECT 220.720 42.180 221.260 42.550 ;
        RECT 221.605 42.470 221.775 43.060 ;
        RECT 221.995 42.640 222.300 43.780 ;
        RECT 222.470 42.590 222.725 43.470 ;
        RECT 223.015 43.150 223.300 43.610 ;
        RECT 223.470 43.320 223.740 43.780 ;
        RECT 223.015 42.930 223.970 43.150 ;
        RECT 221.605 42.440 222.345 42.470 ;
        RECT 220.320 41.840 220.850 42.010 ;
        RECT 218.630 41.420 218.980 41.590 ;
        RECT 219.200 41.400 220.150 41.680 ;
        RECT 220.320 41.230 220.510 41.670 ;
        RECT 220.680 41.610 220.850 41.840 ;
        RECT 221.020 41.780 221.260 42.180 ;
        RECT 221.430 42.140 222.345 42.440 ;
        RECT 221.430 41.965 221.755 42.140 ;
        RECT 221.430 41.610 221.750 41.965 ;
        RECT 222.515 41.940 222.725 42.590 ;
        RECT 222.900 42.200 223.590 42.760 ;
        RECT 223.760 42.030 223.970 42.930 ;
        RECT 220.680 41.440 221.750 41.610 ;
        RECT 221.995 41.230 222.300 41.690 ;
        RECT 222.470 41.410 222.725 41.940 ;
        RECT 223.015 41.860 223.970 42.030 ;
        RECT 224.140 42.760 224.540 43.610 ;
        RECT 224.730 43.150 225.010 43.610 ;
        RECT 225.530 43.320 225.855 43.780 ;
        RECT 224.730 42.930 225.855 43.150 ;
        RECT 224.140 42.200 225.235 42.760 ;
        RECT 225.405 42.470 225.855 42.930 ;
        RECT 226.025 42.640 226.410 43.610 ;
        RECT 223.015 41.400 223.300 41.860 ;
        RECT 223.470 41.230 223.740 41.690 ;
        RECT 224.140 41.400 224.540 42.200 ;
        RECT 225.405 42.140 225.960 42.470 ;
        RECT 225.405 42.030 225.855 42.140 ;
        RECT 224.730 41.860 225.855 42.030 ;
        RECT 226.130 41.970 226.410 42.640 ;
        RECT 226.580 42.615 226.870 43.780 ;
        RECT 227.095 42.910 227.380 43.780 ;
        RECT 227.550 43.150 227.810 43.610 ;
        RECT 227.985 43.320 228.240 43.780 ;
        RECT 228.410 43.150 228.670 43.610 ;
        RECT 227.550 42.980 228.670 43.150 ;
        RECT 228.840 42.980 229.150 43.780 ;
        RECT 227.550 42.730 227.810 42.980 ;
        RECT 229.320 42.810 229.630 43.610 ;
        RECT 230.265 43.110 230.520 43.610 ;
        RECT 230.690 43.280 231.020 43.780 ;
        RECT 230.265 42.940 231.015 43.110 ;
        RECT 224.730 41.400 225.010 41.860 ;
        RECT 225.530 41.230 225.855 41.690 ;
        RECT 226.025 41.400 226.410 41.970 ;
        RECT 227.055 42.560 227.810 42.730 ;
        RECT 228.600 42.640 229.630 42.810 ;
        RECT 227.055 42.050 227.460 42.560 ;
        RECT 228.600 42.390 228.770 42.640 ;
        RECT 227.630 42.220 228.770 42.390 ;
        RECT 226.580 41.230 226.870 41.955 ;
        RECT 227.055 41.880 228.705 42.050 ;
        RECT 228.940 41.900 229.290 42.470 ;
        RECT 227.100 41.230 227.380 41.710 ;
        RECT 227.550 41.490 227.810 41.880 ;
        RECT 227.985 41.230 228.240 41.710 ;
        RECT 228.410 41.490 228.705 41.880 ;
        RECT 229.460 41.730 229.630 42.640 ;
        RECT 230.265 42.120 230.615 42.770 ;
        RECT 230.785 41.950 231.015 42.940 ;
        RECT 228.885 41.230 229.160 41.710 ;
        RECT 229.330 41.400 229.630 41.730 ;
        RECT 230.265 41.780 231.015 41.950 ;
        RECT 230.265 41.490 230.520 41.780 ;
        RECT 230.690 41.230 231.020 41.610 ;
        RECT 231.190 41.490 231.360 43.610 ;
        RECT 231.530 42.810 231.855 43.595 ;
        RECT 232.025 43.320 232.275 43.780 ;
        RECT 232.445 43.280 232.695 43.610 ;
        RECT 232.910 43.280 233.590 43.610 ;
        RECT 232.445 43.150 232.615 43.280 ;
        RECT 232.220 42.980 232.615 43.150 ;
        RECT 231.590 41.760 232.050 42.810 ;
        RECT 232.220 41.620 232.390 42.980 ;
        RECT 232.785 42.720 233.250 43.110 ;
        RECT 232.560 41.910 232.910 42.530 ;
        RECT 233.080 42.130 233.250 42.720 ;
        RECT 233.420 42.500 233.590 43.280 ;
        RECT 233.760 43.180 233.930 43.520 ;
        RECT 234.165 43.350 234.495 43.780 ;
        RECT 234.665 43.180 234.835 43.520 ;
        RECT 235.130 43.320 235.500 43.780 ;
        RECT 233.760 43.010 234.835 43.180 ;
        RECT 235.670 43.150 235.840 43.610 ;
        RECT 236.075 43.270 236.945 43.610 ;
        RECT 237.115 43.320 237.365 43.780 ;
        RECT 235.280 42.980 235.840 43.150 ;
        RECT 235.280 42.840 235.450 42.980 ;
        RECT 233.950 42.670 235.450 42.840 ;
        RECT 236.145 42.810 236.605 43.100 ;
        RECT 233.420 42.330 235.110 42.500 ;
        RECT 233.080 41.910 233.435 42.130 ;
        RECT 233.605 41.620 233.775 42.330 ;
        RECT 233.980 41.910 234.770 42.160 ;
        RECT 234.940 42.150 235.110 42.330 ;
        RECT 235.280 41.980 235.450 42.670 ;
        RECT 231.720 41.230 232.050 41.590 ;
        RECT 232.220 41.450 232.715 41.620 ;
        RECT 232.920 41.450 233.775 41.620 ;
        RECT 234.650 41.230 234.980 41.690 ;
        RECT 235.190 41.590 235.450 41.980 ;
        RECT 235.640 42.800 236.605 42.810 ;
        RECT 236.775 42.890 236.945 43.270 ;
        RECT 237.535 43.230 237.705 43.520 ;
        RECT 237.885 43.400 238.215 43.780 ;
        RECT 237.535 43.060 238.335 43.230 ;
        RECT 235.640 42.640 236.315 42.800 ;
        RECT 236.775 42.720 237.995 42.890 ;
        RECT 235.640 41.850 235.850 42.640 ;
        RECT 236.775 42.630 236.945 42.720 ;
        RECT 236.020 41.850 236.370 42.470 ;
        RECT 236.540 42.460 236.945 42.630 ;
        RECT 236.540 41.680 236.710 42.460 ;
        RECT 236.880 42.010 237.100 42.290 ;
        RECT 237.280 42.180 237.820 42.550 ;
        RECT 238.165 42.470 238.335 43.060 ;
        RECT 238.555 42.640 238.860 43.780 ;
        RECT 239.030 42.590 239.285 43.470 ;
        RECT 238.165 42.440 238.905 42.470 ;
        RECT 236.880 41.840 237.410 42.010 ;
        RECT 235.190 41.420 235.540 41.590 ;
        RECT 235.760 41.400 236.710 41.680 ;
        RECT 236.880 41.230 237.070 41.670 ;
        RECT 237.240 41.610 237.410 41.840 ;
        RECT 237.580 41.780 237.820 42.180 ;
        RECT 237.990 42.140 238.905 42.440 ;
        RECT 237.990 41.965 238.315 42.140 ;
        RECT 237.990 41.610 238.310 41.965 ;
        RECT 239.075 41.940 239.285 42.590 ;
        RECT 237.240 41.440 238.310 41.610 ;
        RECT 238.555 41.230 238.860 41.690 ;
        RECT 239.030 41.410 239.285 41.940 ;
        RECT 239.460 43.020 240.125 43.610 ;
        RECT 239.460 42.050 239.710 43.020 ;
        RECT 240.295 42.940 240.625 43.780 ;
        RECT 241.135 43.190 241.940 43.610 ;
        RECT 240.795 43.020 242.360 43.190 ;
        RECT 240.795 42.770 240.965 43.020 ;
        RECT 240.045 42.600 240.965 42.770 ;
        RECT 241.135 42.760 241.510 42.850 ;
        RECT 240.045 42.430 240.215 42.600 ;
        RECT 241.135 42.590 241.530 42.760 ;
        RECT 241.135 42.430 241.510 42.590 ;
        RECT 239.880 42.220 240.215 42.430 ;
        RECT 240.385 42.220 240.835 42.430 ;
        RECT 241.025 42.220 241.510 42.430 ;
        RECT 241.700 42.470 242.020 42.850 ;
        RECT 242.190 42.770 242.360 43.020 ;
        RECT 242.530 42.940 242.780 43.780 ;
        RECT 242.975 42.770 243.275 43.610 ;
        RECT 242.190 42.600 243.275 42.770 ;
        RECT 243.600 42.640 243.985 43.610 ;
        RECT 244.155 43.320 244.480 43.780 ;
        RECT 245.000 43.150 245.280 43.610 ;
        RECT 244.155 42.930 245.280 43.150 ;
        RECT 241.700 42.220 242.080 42.470 ;
        RECT 242.260 42.220 242.590 42.430 ;
        RECT 239.460 41.410 240.145 42.050 ;
        RECT 240.315 41.230 240.485 42.050 ;
        RECT 240.655 41.880 242.355 42.050 ;
        RECT 240.655 41.415 240.985 41.880 ;
        RECT 241.970 41.790 242.355 41.880 ;
        RECT 242.760 41.970 242.930 42.600 ;
        RECT 243.100 42.140 243.430 42.430 ;
        RECT 243.600 41.970 243.880 42.640 ;
        RECT 244.155 42.470 244.605 42.930 ;
        RECT 245.470 42.760 245.870 43.610 ;
        RECT 246.270 43.320 246.540 43.780 ;
        RECT 246.710 43.150 246.995 43.610 ;
        RECT 244.050 42.140 244.605 42.470 ;
        RECT 244.775 42.200 245.870 42.760 ;
        RECT 244.155 42.030 244.605 42.140 ;
        RECT 242.760 41.790 243.270 41.970 ;
        RECT 241.155 41.230 241.325 41.700 ;
        RECT 241.585 41.450 242.770 41.620 ;
        RECT 242.940 41.400 243.270 41.790 ;
        RECT 243.600 41.400 243.985 41.970 ;
        RECT 244.155 41.860 245.280 42.030 ;
        RECT 244.155 41.230 244.480 41.690 ;
        RECT 245.000 41.400 245.280 41.860 ;
        RECT 245.470 41.400 245.870 42.200 ;
        RECT 246.040 42.930 246.995 43.150 ;
        RECT 246.040 42.030 246.250 42.930 ;
        RECT 246.420 42.200 247.110 42.760 ;
        RECT 247.280 42.690 248.490 43.780 ;
        RECT 248.775 43.150 249.060 43.610 ;
        RECT 249.230 43.320 249.500 43.780 ;
        RECT 248.775 42.930 249.730 43.150 ;
        RECT 246.040 41.860 246.995 42.030 ;
        RECT 246.270 41.230 246.540 41.690 ;
        RECT 246.710 41.400 246.995 41.860 ;
        RECT 247.280 41.980 247.800 42.520 ;
        RECT 247.970 42.150 248.490 42.690 ;
        RECT 248.660 42.200 249.350 42.760 ;
        RECT 249.520 42.030 249.730 42.930 ;
        RECT 247.280 41.230 248.490 41.980 ;
        RECT 248.775 41.860 249.730 42.030 ;
        RECT 249.900 42.760 250.300 43.610 ;
        RECT 250.490 43.150 250.770 43.610 ;
        RECT 251.290 43.320 251.615 43.780 ;
        RECT 250.490 42.930 251.615 43.150 ;
        RECT 249.900 42.200 250.995 42.760 ;
        RECT 251.165 42.470 251.615 42.930 ;
        RECT 251.785 42.640 252.170 43.610 ;
        RECT 248.775 41.400 249.060 41.860 ;
        RECT 249.230 41.230 249.500 41.690 ;
        RECT 249.900 41.400 250.300 42.200 ;
        RECT 251.165 42.140 251.720 42.470 ;
        RECT 251.165 42.030 251.615 42.140 ;
        RECT 250.490 41.860 251.615 42.030 ;
        RECT 251.890 41.970 252.170 42.640 ;
        RECT 252.340 42.615 252.630 43.780 ;
        RECT 252.800 42.810 253.110 43.610 ;
        RECT 253.280 42.980 253.590 43.780 ;
        RECT 253.760 43.150 254.020 43.610 ;
        RECT 254.190 43.320 254.445 43.780 ;
        RECT 254.620 43.150 254.880 43.610 ;
        RECT 253.760 42.980 254.880 43.150 ;
        RECT 252.800 42.640 253.830 42.810 ;
        RECT 250.490 41.400 250.770 41.860 ;
        RECT 251.290 41.230 251.615 41.690 ;
        RECT 251.785 41.400 252.170 41.970 ;
        RECT 252.340 41.230 252.630 41.955 ;
        RECT 252.800 41.730 252.970 42.640 ;
        RECT 253.140 41.900 253.490 42.470 ;
        RECT 253.660 42.390 253.830 42.640 ;
        RECT 254.620 42.730 254.880 42.980 ;
        RECT 255.050 42.910 255.335 43.780 ;
        RECT 254.620 42.560 255.375 42.730 ;
        RECT 255.560 42.690 257.230 43.780 ;
        RECT 253.660 42.220 254.800 42.390 ;
        RECT 254.970 42.050 255.375 42.560 ;
        RECT 253.725 41.880 255.375 42.050 ;
        RECT 255.560 42.000 256.310 42.520 ;
        RECT 256.480 42.170 257.230 42.690 ;
        RECT 257.895 42.990 258.430 43.610 ;
        RECT 252.800 41.400 253.100 41.730 ;
        RECT 253.270 41.230 253.545 41.710 ;
        RECT 253.725 41.490 254.020 41.880 ;
        RECT 254.190 41.230 254.445 41.710 ;
        RECT 254.620 41.490 254.880 41.880 ;
        RECT 255.050 41.230 255.330 41.710 ;
        RECT 255.560 41.230 257.230 42.000 ;
        RECT 257.895 41.970 258.210 42.990 ;
        RECT 258.600 42.980 258.930 43.780 ;
        RECT 259.415 42.810 259.805 42.985 ;
        RECT 258.380 42.640 259.805 42.810 ;
        RECT 260.345 42.810 260.735 42.985 ;
        RECT 261.220 42.980 261.550 43.780 ;
        RECT 261.720 42.990 262.255 43.610 ;
        RECT 260.345 42.640 261.770 42.810 ;
        RECT 258.380 42.140 258.550 42.640 ;
        RECT 257.895 41.400 258.510 41.970 ;
        RECT 258.800 41.910 259.065 42.470 ;
        RECT 259.235 41.740 259.405 42.640 ;
        RECT 259.575 41.910 259.930 42.470 ;
        RECT 260.220 41.910 260.575 42.470 ;
        RECT 260.745 41.740 260.915 42.640 ;
        RECT 261.085 41.910 261.350 42.470 ;
        RECT 261.600 42.140 261.770 42.640 ;
        RECT 261.940 41.970 262.255 42.990 ;
        RECT 262.460 42.690 264.130 43.780 ;
        RECT 258.680 41.230 258.895 41.740 ;
        RECT 259.125 41.410 259.405 41.740 ;
        RECT 259.585 41.230 259.825 41.740 ;
        RECT 260.325 41.230 260.565 41.740 ;
        RECT 260.745 41.410 261.025 41.740 ;
        RECT 261.255 41.230 261.470 41.740 ;
        RECT 261.640 41.400 262.255 41.970 ;
        RECT 262.460 42.000 263.210 42.520 ;
        RECT 263.380 42.170 264.130 42.690 ;
        RECT 264.340 42.640 264.570 43.780 ;
        RECT 264.740 42.630 265.070 43.610 ;
        RECT 265.240 42.640 265.450 43.780 ;
        RECT 265.680 42.690 266.890 43.780 ;
        RECT 267.065 43.110 267.320 43.610 ;
        RECT 267.490 43.280 267.820 43.780 ;
        RECT 267.065 42.940 267.815 43.110 ;
        RECT 264.320 42.220 264.650 42.470 ;
        RECT 262.460 41.230 264.130 42.000 ;
        RECT 264.340 41.230 264.570 42.050 ;
        RECT 264.820 42.030 265.070 42.630 ;
        RECT 264.740 41.400 265.070 42.030 ;
        RECT 265.240 41.230 265.450 42.050 ;
        RECT 265.680 41.980 266.200 42.520 ;
        RECT 266.370 42.150 266.890 42.690 ;
        RECT 267.065 42.120 267.415 42.770 ;
        RECT 265.680 41.230 266.890 41.980 ;
        RECT 267.585 41.950 267.815 42.940 ;
        RECT 267.065 41.780 267.815 41.950 ;
        RECT 267.065 41.490 267.320 41.780 ;
        RECT 267.490 41.230 267.820 41.610 ;
        RECT 267.990 41.490 268.160 43.610 ;
        RECT 268.330 42.810 268.655 43.595 ;
        RECT 268.825 43.320 269.075 43.780 ;
        RECT 269.245 43.280 269.495 43.610 ;
        RECT 269.710 43.280 270.390 43.610 ;
        RECT 269.245 43.150 269.415 43.280 ;
        RECT 269.020 42.980 269.415 43.150 ;
        RECT 268.390 41.760 268.850 42.810 ;
        RECT 269.020 41.620 269.190 42.980 ;
        RECT 269.585 42.720 270.050 43.110 ;
        RECT 269.360 41.910 269.710 42.530 ;
        RECT 269.880 42.130 270.050 42.720 ;
        RECT 270.220 42.500 270.390 43.280 ;
        RECT 270.560 43.180 270.730 43.520 ;
        RECT 270.965 43.350 271.295 43.780 ;
        RECT 271.465 43.180 271.635 43.520 ;
        RECT 271.930 43.320 272.300 43.780 ;
        RECT 270.560 43.010 271.635 43.180 ;
        RECT 272.470 43.150 272.640 43.610 ;
        RECT 272.875 43.270 273.745 43.610 ;
        RECT 273.915 43.320 274.165 43.780 ;
        RECT 272.080 42.980 272.640 43.150 ;
        RECT 272.080 42.840 272.250 42.980 ;
        RECT 270.750 42.670 272.250 42.840 ;
        RECT 272.945 42.810 273.405 43.100 ;
        RECT 270.220 42.330 271.910 42.500 ;
        RECT 269.880 41.910 270.235 42.130 ;
        RECT 270.405 41.620 270.575 42.330 ;
        RECT 270.780 41.910 271.570 42.160 ;
        RECT 271.740 42.150 271.910 42.330 ;
        RECT 272.080 41.980 272.250 42.670 ;
        RECT 268.520 41.230 268.850 41.590 ;
        RECT 269.020 41.450 269.515 41.620 ;
        RECT 269.720 41.450 270.575 41.620 ;
        RECT 271.450 41.230 271.780 41.690 ;
        RECT 271.990 41.590 272.250 41.980 ;
        RECT 272.440 42.800 273.405 42.810 ;
        RECT 273.575 42.890 273.745 43.270 ;
        RECT 274.335 43.230 274.505 43.520 ;
        RECT 274.685 43.400 275.015 43.780 ;
        RECT 274.335 43.060 275.135 43.230 ;
        RECT 272.440 42.640 273.115 42.800 ;
        RECT 273.575 42.720 274.795 42.890 ;
        RECT 272.440 41.850 272.650 42.640 ;
        RECT 273.575 42.630 273.745 42.720 ;
        RECT 272.820 41.850 273.170 42.470 ;
        RECT 273.340 42.460 273.745 42.630 ;
        RECT 273.340 41.680 273.510 42.460 ;
        RECT 273.680 42.010 273.900 42.290 ;
        RECT 274.080 42.180 274.620 42.550 ;
        RECT 274.965 42.470 275.135 43.060 ;
        RECT 275.355 42.640 275.660 43.780 ;
        RECT 275.830 42.590 276.085 43.470 ;
        RECT 276.265 42.980 276.520 43.780 ;
        RECT 276.720 42.930 277.050 43.610 ;
        RECT 274.965 42.440 275.705 42.470 ;
        RECT 273.680 41.840 274.210 42.010 ;
        RECT 271.990 41.420 272.340 41.590 ;
        RECT 272.560 41.400 273.510 41.680 ;
        RECT 273.680 41.230 273.870 41.670 ;
        RECT 274.040 41.610 274.210 41.840 ;
        RECT 274.380 41.780 274.620 42.180 ;
        RECT 274.790 42.140 275.705 42.440 ;
        RECT 274.790 41.965 275.115 42.140 ;
        RECT 274.790 41.610 275.110 41.965 ;
        RECT 275.875 41.940 276.085 42.590 ;
        RECT 276.265 42.440 276.510 42.800 ;
        RECT 276.700 42.650 277.050 42.930 ;
        RECT 276.700 42.270 276.870 42.650 ;
        RECT 277.230 42.470 277.425 43.520 ;
        RECT 277.605 42.640 277.925 43.780 ;
        RECT 278.100 42.615 278.390 43.780 ;
        RECT 278.570 43.170 278.900 43.600 ;
        RECT 279.080 43.340 279.275 43.780 ;
        RECT 279.445 43.170 279.775 43.600 ;
        RECT 278.570 43.000 279.775 43.170 ;
        RECT 278.570 42.670 279.465 43.000 ;
        RECT 279.945 42.830 280.220 43.600 ;
        RECT 279.635 42.640 280.220 42.830 ;
        RECT 280.860 42.640 281.245 43.610 ;
        RECT 281.415 43.320 281.740 43.780 ;
        RECT 282.260 43.150 282.540 43.610 ;
        RECT 281.415 42.930 282.540 43.150 ;
        RECT 274.040 41.440 275.110 41.610 ;
        RECT 275.355 41.230 275.660 41.690 ;
        RECT 275.830 41.410 276.085 41.940 ;
        RECT 276.350 42.100 276.870 42.270 ;
        RECT 277.040 42.140 277.425 42.470 ;
        RECT 277.605 42.140 277.865 42.470 ;
        RECT 278.575 42.140 278.870 42.470 ;
        RECT 279.050 42.140 279.465 42.470 ;
        RECT 276.350 41.535 276.520 42.100 ;
        RECT 276.710 41.760 277.925 41.930 ;
        RECT 276.710 41.455 276.940 41.760 ;
        RECT 277.110 41.230 277.440 41.590 ;
        RECT 277.635 41.410 277.925 41.760 ;
        RECT 278.100 41.230 278.390 41.955 ;
        RECT 278.570 41.230 278.870 41.960 ;
        RECT 279.050 41.520 279.280 42.140 ;
        RECT 279.635 41.970 279.810 42.640 ;
        RECT 279.480 41.790 279.810 41.970 ;
        RECT 279.980 41.820 280.220 42.470 ;
        RECT 280.860 41.970 281.140 42.640 ;
        RECT 281.415 42.470 281.865 42.930 ;
        RECT 282.730 42.760 283.130 43.610 ;
        RECT 283.530 43.320 283.800 43.780 ;
        RECT 283.970 43.150 284.255 43.610 ;
        RECT 281.310 42.140 281.865 42.470 ;
        RECT 282.035 42.200 283.130 42.760 ;
        RECT 281.415 42.030 281.865 42.140 ;
        RECT 279.480 41.410 279.705 41.790 ;
        RECT 279.875 41.230 280.205 41.620 ;
        RECT 280.860 41.400 281.245 41.970 ;
        RECT 281.415 41.860 282.540 42.030 ;
        RECT 281.415 41.230 281.740 41.690 ;
        RECT 282.260 41.400 282.540 41.860 ;
        RECT 282.730 41.400 283.130 42.200 ;
        RECT 283.300 42.930 284.255 43.150 ;
        RECT 283.300 42.030 283.510 42.930 ;
        RECT 283.680 42.200 284.370 42.760 ;
        RECT 284.580 42.640 284.810 43.780 ;
        RECT 284.980 42.630 285.310 43.610 ;
        RECT 285.480 42.640 285.690 43.780 ;
        RECT 285.920 42.640 286.305 43.610 ;
        RECT 286.475 43.320 286.800 43.780 ;
        RECT 287.320 43.150 287.600 43.610 ;
        RECT 286.475 42.930 287.600 43.150 ;
        RECT 284.560 42.220 284.890 42.470 ;
        RECT 283.300 41.860 284.255 42.030 ;
        RECT 283.530 41.230 283.800 41.690 ;
        RECT 283.970 41.400 284.255 41.860 ;
        RECT 284.580 41.230 284.810 42.050 ;
        RECT 285.060 42.030 285.310 42.630 ;
        RECT 284.980 41.400 285.310 42.030 ;
        RECT 285.480 41.230 285.690 42.050 ;
        RECT 285.920 41.970 286.200 42.640 ;
        RECT 286.475 42.470 286.925 42.930 ;
        RECT 287.790 42.760 288.190 43.610 ;
        RECT 288.590 43.320 288.860 43.780 ;
        RECT 289.030 43.150 289.315 43.610 ;
        RECT 289.600 43.345 294.945 43.780 ;
        RECT 295.120 43.345 300.465 43.780 ;
        RECT 286.370 42.140 286.925 42.470 ;
        RECT 287.095 42.200 288.190 42.760 ;
        RECT 286.475 42.030 286.925 42.140 ;
        RECT 285.920 41.400 286.305 41.970 ;
        RECT 286.475 41.860 287.600 42.030 ;
        RECT 286.475 41.230 286.800 41.690 ;
        RECT 287.320 41.400 287.600 41.860 ;
        RECT 287.790 41.400 288.190 42.200 ;
        RECT 288.360 42.930 289.315 43.150 ;
        RECT 288.360 42.030 288.570 42.930 ;
        RECT 288.740 42.200 289.430 42.760 ;
        RECT 288.360 41.860 289.315 42.030 ;
        RECT 288.590 41.230 288.860 41.690 ;
        RECT 289.030 41.400 289.315 41.860 ;
        RECT 291.185 41.775 291.525 42.605 ;
        RECT 293.005 42.095 293.355 43.345 ;
        RECT 296.705 41.775 297.045 42.605 ;
        RECT 298.525 42.095 298.875 43.345 ;
        RECT 300.640 42.690 303.230 43.780 ;
        RECT 300.640 42.000 301.850 42.520 ;
        RECT 302.020 42.170 303.230 42.690 ;
        RECT 303.860 42.615 304.150 43.780 ;
        RECT 304.320 42.690 305.990 43.780 ;
        RECT 304.320 42.000 305.070 42.520 ;
        RECT 305.240 42.170 305.990 42.690 ;
        RECT 306.250 42.850 306.420 43.610 ;
        RECT 306.635 43.020 306.965 43.780 ;
        RECT 306.250 42.680 306.965 42.850 ;
        RECT 307.135 42.705 307.390 43.610 ;
        RECT 306.160 42.130 306.515 42.500 ;
        RECT 306.795 42.470 306.965 42.680 ;
        RECT 306.795 42.140 307.050 42.470 ;
        RECT 289.600 41.230 294.945 41.775 ;
        RECT 295.120 41.230 300.465 41.775 ;
        RECT 300.640 41.230 303.230 42.000 ;
        RECT 303.860 41.230 304.150 41.955 ;
        RECT 304.320 41.230 305.990 42.000 ;
        RECT 306.795 41.950 306.965 42.140 ;
        RECT 307.220 41.975 307.390 42.705 ;
        RECT 307.565 42.630 307.825 43.780 ;
        RECT 308.000 42.690 309.670 43.780 ;
        RECT 306.250 41.780 306.965 41.950 ;
        RECT 306.250 41.400 306.420 41.780 ;
        RECT 306.635 41.230 306.965 41.610 ;
        RECT 307.135 41.400 307.390 41.975 ;
        RECT 307.565 41.230 307.825 42.070 ;
        RECT 308.000 42.000 308.750 42.520 ;
        RECT 308.920 42.170 309.670 42.690 ;
        RECT 309.840 42.690 311.050 43.780 ;
        RECT 309.840 42.150 310.360 42.690 ;
        RECT 308.000 41.230 309.670 42.000 ;
        RECT 310.530 41.980 311.050 42.520 ;
        RECT 309.840 41.230 311.050 41.980 ;
        RECT 162.095 41.060 311.135 41.230 ;
        RECT 162.180 40.310 163.390 41.060 ;
        RECT 164.135 40.430 164.420 40.890 ;
        RECT 164.590 40.600 164.860 41.060 ;
        RECT 162.180 39.770 162.700 40.310 ;
        RECT 164.135 40.260 165.090 40.430 ;
        RECT 162.870 39.600 163.390 40.140 ;
        RECT 162.180 38.510 163.390 39.600 ;
        RECT 164.020 39.530 164.710 40.090 ;
        RECT 164.880 39.360 165.090 40.260 ;
        RECT 164.135 39.140 165.090 39.360 ;
        RECT 165.260 40.090 165.660 40.890 ;
        RECT 165.850 40.430 166.130 40.890 ;
        RECT 166.650 40.600 166.975 41.060 ;
        RECT 165.850 40.260 166.975 40.430 ;
        RECT 167.145 40.320 167.530 40.890 ;
        RECT 166.525 40.150 166.975 40.260 ;
        RECT 165.260 39.530 166.355 40.090 ;
        RECT 166.525 39.820 167.080 40.150 ;
        RECT 164.135 38.680 164.420 39.140 ;
        RECT 164.590 38.510 164.860 38.970 ;
        RECT 165.260 38.680 165.660 39.530 ;
        RECT 166.525 39.360 166.975 39.820 ;
        RECT 167.250 39.650 167.530 40.320 ;
        RECT 165.850 39.140 166.975 39.360 ;
        RECT 165.850 38.680 166.130 39.140 ;
        RECT 166.650 38.510 166.975 38.970 ;
        RECT 167.145 38.680 167.530 39.650 ;
        RECT 167.705 40.350 167.960 40.880 ;
        RECT 168.130 40.600 168.435 41.060 ;
        RECT 168.680 40.680 169.750 40.850 ;
        RECT 167.705 39.700 167.915 40.350 ;
        RECT 168.680 40.325 169.000 40.680 ;
        RECT 168.675 40.150 169.000 40.325 ;
        RECT 168.085 39.850 169.000 40.150 ;
        RECT 169.170 40.110 169.410 40.510 ;
        RECT 169.580 40.450 169.750 40.680 ;
        RECT 169.920 40.620 170.110 41.060 ;
        RECT 170.280 40.610 171.230 40.890 ;
        RECT 171.450 40.700 171.800 40.870 ;
        RECT 169.580 40.280 170.110 40.450 ;
        RECT 168.085 39.820 168.825 39.850 ;
        RECT 167.705 38.820 167.960 39.700 ;
        RECT 168.130 38.510 168.435 39.650 ;
        RECT 168.655 39.230 168.825 39.820 ;
        RECT 169.170 39.740 169.710 40.110 ;
        RECT 169.890 40.000 170.110 40.280 ;
        RECT 170.280 39.830 170.450 40.610 ;
        RECT 170.045 39.660 170.450 39.830 ;
        RECT 170.620 39.820 170.970 40.440 ;
        RECT 170.045 39.570 170.215 39.660 ;
        RECT 171.140 39.650 171.350 40.440 ;
        RECT 168.995 39.400 170.215 39.570 ;
        RECT 170.675 39.490 171.350 39.650 ;
        RECT 168.655 39.060 169.455 39.230 ;
        RECT 168.775 38.510 169.105 38.890 ;
        RECT 169.285 38.770 169.455 39.060 ;
        RECT 170.045 39.020 170.215 39.400 ;
        RECT 170.385 39.480 171.350 39.490 ;
        RECT 171.540 40.310 171.800 40.700 ;
        RECT 172.010 40.600 172.340 41.060 ;
        RECT 173.215 40.670 174.070 40.840 ;
        RECT 174.275 40.670 174.770 40.840 ;
        RECT 174.940 40.700 175.270 41.060 ;
        RECT 171.540 39.620 171.710 40.310 ;
        RECT 171.880 39.960 172.050 40.140 ;
        RECT 172.220 40.130 173.010 40.380 ;
        RECT 173.215 39.960 173.385 40.670 ;
        RECT 173.555 40.160 173.910 40.380 ;
        RECT 171.880 39.790 173.570 39.960 ;
        RECT 170.385 39.190 170.845 39.480 ;
        RECT 171.540 39.450 173.040 39.620 ;
        RECT 171.540 39.310 171.710 39.450 ;
        RECT 171.150 39.140 171.710 39.310 ;
        RECT 169.625 38.510 169.875 38.970 ;
        RECT 170.045 38.680 170.915 39.020 ;
        RECT 171.150 38.680 171.320 39.140 ;
        RECT 172.155 39.110 173.230 39.280 ;
        RECT 171.490 38.510 171.860 38.970 ;
        RECT 172.155 38.770 172.325 39.110 ;
        RECT 172.495 38.510 172.825 38.940 ;
        RECT 173.060 38.770 173.230 39.110 ;
        RECT 173.400 39.010 173.570 39.790 ;
        RECT 173.740 39.570 173.910 40.160 ;
        RECT 174.080 39.760 174.430 40.380 ;
        RECT 173.740 39.180 174.205 39.570 ;
        RECT 174.600 39.310 174.770 40.670 ;
        RECT 174.940 39.480 175.400 40.530 ;
        RECT 174.375 39.140 174.770 39.310 ;
        RECT 174.375 39.010 174.545 39.140 ;
        RECT 173.400 38.680 174.080 39.010 ;
        RECT 174.295 38.680 174.545 39.010 ;
        RECT 174.715 38.510 174.965 38.970 ;
        RECT 175.135 38.695 175.460 39.480 ;
        RECT 175.630 38.680 175.800 40.800 ;
        RECT 175.970 40.680 176.300 41.060 ;
        RECT 176.470 40.510 176.725 40.800 ;
        RECT 175.975 40.340 176.725 40.510 ;
        RECT 175.975 39.350 176.205 40.340 ;
        RECT 176.905 40.320 177.160 40.890 ;
        RECT 177.330 40.660 177.660 41.060 ;
        RECT 178.085 40.525 178.615 40.890 ;
        RECT 178.805 40.720 179.080 40.890 ;
        RECT 178.800 40.550 179.080 40.720 ;
        RECT 178.085 40.490 178.260 40.525 ;
        RECT 177.330 40.320 178.260 40.490 ;
        RECT 176.375 39.520 176.725 40.170 ;
        RECT 176.905 39.650 177.075 40.320 ;
        RECT 177.330 40.150 177.500 40.320 ;
        RECT 177.245 39.820 177.500 40.150 ;
        RECT 177.725 39.820 177.920 40.150 ;
        RECT 175.975 39.180 176.725 39.350 ;
        RECT 175.970 38.510 176.300 39.010 ;
        RECT 176.470 38.680 176.725 39.180 ;
        RECT 176.905 38.680 177.240 39.650 ;
        RECT 177.410 38.510 177.580 39.650 ;
        RECT 177.750 38.850 177.920 39.820 ;
        RECT 178.090 39.190 178.260 40.320 ;
        RECT 178.430 39.530 178.600 40.330 ;
        RECT 178.805 39.730 179.080 40.550 ;
        RECT 179.250 39.530 179.440 40.890 ;
        RECT 179.620 40.525 180.130 41.060 ;
        RECT 180.350 40.250 180.595 40.855 ;
        RECT 181.040 40.290 183.630 41.060 ;
        RECT 184.260 40.320 184.645 40.890 ;
        RECT 184.815 40.600 185.140 41.060 ;
        RECT 185.660 40.430 185.940 40.890 ;
        RECT 179.640 40.080 180.870 40.250 ;
        RECT 178.430 39.360 179.440 39.530 ;
        RECT 179.610 39.515 180.360 39.705 ;
        RECT 178.090 39.020 179.215 39.190 ;
        RECT 179.610 38.850 179.780 39.515 ;
        RECT 180.530 39.270 180.870 40.080 ;
        RECT 181.040 39.770 182.250 40.290 ;
        RECT 182.420 39.600 183.630 40.120 ;
        RECT 177.750 38.680 179.780 38.850 ;
        RECT 179.950 38.510 180.120 39.270 ;
        RECT 180.355 38.860 180.870 39.270 ;
        RECT 181.040 38.510 183.630 39.600 ;
        RECT 184.260 39.650 184.540 40.320 ;
        RECT 184.815 40.260 185.940 40.430 ;
        RECT 184.815 40.150 185.265 40.260 ;
        RECT 184.710 39.820 185.265 40.150 ;
        RECT 186.130 40.090 186.530 40.890 ;
        RECT 186.930 40.600 187.200 41.060 ;
        RECT 187.370 40.430 187.655 40.890 ;
        RECT 184.260 38.680 184.645 39.650 ;
        RECT 184.815 39.360 185.265 39.820 ;
        RECT 185.435 39.530 186.530 40.090 ;
        RECT 184.815 39.140 185.940 39.360 ;
        RECT 184.815 38.510 185.140 38.970 ;
        RECT 185.660 38.680 185.940 39.140 ;
        RECT 186.130 38.680 186.530 39.530 ;
        RECT 186.700 40.260 187.655 40.430 ;
        RECT 187.940 40.335 188.230 41.060 ;
        RECT 188.405 40.320 188.660 40.890 ;
        RECT 188.830 40.660 189.160 41.060 ;
        RECT 189.585 40.525 190.115 40.890 ;
        RECT 190.305 40.720 190.580 40.890 ;
        RECT 190.300 40.550 190.580 40.720 ;
        RECT 189.585 40.490 189.760 40.525 ;
        RECT 188.830 40.320 189.760 40.490 ;
        RECT 186.700 39.360 186.910 40.260 ;
        RECT 187.080 39.530 187.770 40.090 ;
        RECT 186.700 39.140 187.655 39.360 ;
        RECT 186.930 38.510 187.200 38.970 ;
        RECT 187.370 38.680 187.655 39.140 ;
        RECT 187.940 38.510 188.230 39.675 ;
        RECT 188.405 39.650 188.575 40.320 ;
        RECT 188.830 40.150 189.000 40.320 ;
        RECT 188.745 39.820 189.000 40.150 ;
        RECT 189.225 39.820 189.420 40.150 ;
        RECT 188.405 38.680 188.740 39.650 ;
        RECT 188.910 38.510 189.080 39.650 ;
        RECT 189.250 38.850 189.420 39.820 ;
        RECT 189.590 39.190 189.760 40.320 ;
        RECT 189.930 39.530 190.100 40.330 ;
        RECT 190.305 39.730 190.580 40.550 ;
        RECT 190.750 39.530 190.940 40.890 ;
        RECT 191.120 40.525 191.630 41.060 ;
        RECT 191.850 40.250 192.095 40.855 ;
        RECT 192.545 40.660 192.880 41.060 ;
        RECT 193.050 40.490 193.255 40.890 ;
        RECT 193.465 40.580 193.740 41.060 ;
        RECT 193.950 40.560 194.210 40.890 ;
        RECT 192.570 40.320 193.255 40.490 ;
        RECT 191.140 40.080 192.370 40.250 ;
        RECT 189.930 39.360 190.940 39.530 ;
        RECT 191.110 39.515 191.860 39.705 ;
        RECT 189.590 39.020 190.715 39.190 ;
        RECT 191.110 38.850 191.280 39.515 ;
        RECT 192.030 39.270 192.370 40.080 ;
        RECT 189.250 38.680 191.280 38.850 ;
        RECT 191.450 38.510 191.620 39.270 ;
        RECT 191.855 38.860 192.370 39.270 ;
        RECT 192.570 39.290 192.910 40.320 ;
        RECT 193.080 39.650 193.330 40.150 ;
        RECT 193.510 39.820 193.870 40.400 ;
        RECT 194.040 39.650 194.210 40.560 ;
        RECT 194.380 40.310 195.590 41.060 ;
        RECT 195.765 40.510 196.020 40.800 ;
        RECT 196.190 40.680 196.520 41.060 ;
        RECT 195.765 40.340 196.515 40.510 ;
        RECT 194.380 39.770 194.900 40.310 ;
        RECT 193.080 39.480 194.210 39.650 ;
        RECT 195.070 39.600 195.590 40.140 ;
        RECT 192.570 39.115 193.235 39.290 ;
        RECT 192.545 38.510 192.880 38.935 ;
        RECT 193.050 38.710 193.235 39.115 ;
        RECT 193.440 38.510 193.770 39.290 ;
        RECT 193.940 38.710 194.210 39.480 ;
        RECT 194.380 38.510 195.590 39.600 ;
        RECT 195.765 39.520 196.115 40.170 ;
        RECT 196.285 39.350 196.515 40.340 ;
        RECT 195.765 39.180 196.515 39.350 ;
        RECT 195.765 38.680 196.020 39.180 ;
        RECT 196.190 38.510 196.520 39.010 ;
        RECT 196.690 38.680 196.860 40.800 ;
        RECT 197.220 40.700 197.550 41.060 ;
        RECT 197.720 40.670 198.215 40.840 ;
        RECT 198.420 40.670 199.275 40.840 ;
        RECT 197.090 39.480 197.550 40.530 ;
        RECT 197.030 38.695 197.355 39.480 ;
        RECT 197.720 39.310 197.890 40.670 ;
        RECT 198.060 39.760 198.410 40.380 ;
        RECT 198.580 40.160 198.935 40.380 ;
        RECT 198.580 39.570 198.750 40.160 ;
        RECT 199.105 39.960 199.275 40.670 ;
        RECT 200.150 40.600 200.480 41.060 ;
        RECT 200.690 40.700 201.040 40.870 ;
        RECT 199.480 40.130 200.270 40.380 ;
        RECT 200.690 40.310 200.950 40.700 ;
        RECT 201.260 40.610 202.210 40.890 ;
        RECT 202.380 40.620 202.570 41.060 ;
        RECT 202.740 40.680 203.810 40.850 ;
        RECT 200.440 39.960 200.610 40.140 ;
        RECT 197.720 39.140 198.115 39.310 ;
        RECT 198.285 39.180 198.750 39.570 ;
        RECT 198.920 39.790 200.610 39.960 ;
        RECT 197.945 39.010 198.115 39.140 ;
        RECT 198.920 39.010 199.090 39.790 ;
        RECT 200.780 39.620 200.950 40.310 ;
        RECT 199.450 39.450 200.950 39.620 ;
        RECT 201.140 39.650 201.350 40.440 ;
        RECT 201.520 39.820 201.870 40.440 ;
        RECT 202.040 39.830 202.210 40.610 ;
        RECT 202.740 40.450 202.910 40.680 ;
        RECT 202.380 40.280 202.910 40.450 ;
        RECT 202.380 40.000 202.600 40.280 ;
        RECT 203.080 40.110 203.320 40.510 ;
        RECT 202.040 39.660 202.445 39.830 ;
        RECT 202.780 39.740 203.320 40.110 ;
        RECT 203.490 40.325 203.810 40.680 ;
        RECT 204.055 40.600 204.360 41.060 ;
        RECT 204.530 40.350 204.785 40.880 ;
        RECT 203.490 40.150 203.815 40.325 ;
        RECT 203.490 39.850 204.405 40.150 ;
        RECT 203.665 39.820 204.405 39.850 ;
        RECT 201.140 39.490 201.815 39.650 ;
        RECT 202.275 39.570 202.445 39.660 ;
        RECT 201.140 39.480 202.105 39.490 ;
        RECT 200.780 39.310 200.950 39.450 ;
        RECT 197.525 38.510 197.775 38.970 ;
        RECT 197.945 38.680 198.195 39.010 ;
        RECT 198.410 38.680 199.090 39.010 ;
        RECT 199.260 39.110 200.335 39.280 ;
        RECT 200.780 39.140 201.340 39.310 ;
        RECT 201.645 39.190 202.105 39.480 ;
        RECT 202.275 39.400 203.495 39.570 ;
        RECT 199.260 38.770 199.430 39.110 ;
        RECT 199.665 38.510 199.995 38.940 ;
        RECT 200.165 38.770 200.335 39.110 ;
        RECT 200.630 38.510 201.000 38.970 ;
        RECT 201.170 38.680 201.340 39.140 ;
        RECT 202.275 39.020 202.445 39.400 ;
        RECT 203.665 39.230 203.835 39.820 ;
        RECT 204.575 39.700 204.785 40.350 ;
        RECT 201.575 38.680 202.445 39.020 ;
        RECT 203.035 39.060 203.835 39.230 ;
        RECT 202.615 38.510 202.865 38.970 ;
        RECT 203.035 38.770 203.205 39.060 ;
        RECT 203.385 38.510 203.715 38.890 ;
        RECT 204.055 38.510 204.360 39.650 ;
        RECT 204.530 38.820 204.785 39.700 ;
        RECT 204.960 40.320 205.345 40.890 ;
        RECT 205.515 40.600 205.840 41.060 ;
        RECT 206.360 40.430 206.640 40.890 ;
        RECT 204.960 39.650 205.240 40.320 ;
        RECT 205.515 40.260 206.640 40.430 ;
        RECT 205.515 40.150 205.965 40.260 ;
        RECT 205.410 39.820 205.965 40.150 ;
        RECT 206.830 40.090 207.230 40.890 ;
        RECT 207.630 40.600 207.900 41.060 ;
        RECT 208.070 40.430 208.355 40.890 ;
        RECT 204.960 38.680 205.345 39.650 ;
        RECT 205.515 39.360 205.965 39.820 ;
        RECT 206.135 39.530 207.230 40.090 ;
        RECT 205.515 39.140 206.640 39.360 ;
        RECT 205.515 38.510 205.840 38.970 ;
        RECT 206.360 38.680 206.640 39.140 ;
        RECT 206.830 38.680 207.230 39.530 ;
        RECT 207.400 40.260 208.355 40.430 ;
        RECT 208.640 40.310 209.850 41.060 ;
        RECT 210.020 40.320 210.405 40.890 ;
        RECT 210.575 40.600 210.900 41.060 ;
        RECT 211.420 40.430 211.700 40.890 ;
        RECT 207.400 39.360 207.610 40.260 ;
        RECT 207.780 39.530 208.470 40.090 ;
        RECT 208.640 39.770 209.160 40.310 ;
        RECT 209.330 39.600 209.850 40.140 ;
        RECT 207.400 39.140 208.355 39.360 ;
        RECT 207.630 38.510 207.900 38.970 ;
        RECT 208.070 38.680 208.355 39.140 ;
        RECT 208.640 38.510 209.850 39.600 ;
        RECT 210.020 39.650 210.300 40.320 ;
        RECT 210.575 40.260 211.700 40.430 ;
        RECT 210.575 40.150 211.025 40.260 ;
        RECT 210.470 39.820 211.025 40.150 ;
        RECT 211.890 40.090 212.290 40.890 ;
        RECT 212.690 40.600 212.960 41.060 ;
        RECT 213.130 40.430 213.415 40.890 ;
        RECT 210.020 38.680 210.405 39.650 ;
        RECT 210.575 39.360 211.025 39.820 ;
        RECT 211.195 39.530 212.290 40.090 ;
        RECT 210.575 39.140 211.700 39.360 ;
        RECT 210.575 38.510 210.900 38.970 ;
        RECT 211.420 38.680 211.700 39.140 ;
        RECT 211.890 38.680 212.290 39.530 ;
        RECT 212.460 40.260 213.415 40.430 ;
        RECT 213.700 40.335 213.990 41.060 ;
        RECT 214.165 40.350 214.420 40.880 ;
        RECT 214.590 40.600 214.895 41.060 ;
        RECT 215.140 40.680 216.210 40.850 ;
        RECT 212.460 39.360 212.670 40.260 ;
        RECT 212.840 39.530 213.530 40.090 ;
        RECT 214.165 39.700 214.375 40.350 ;
        RECT 215.140 40.325 215.460 40.680 ;
        RECT 215.135 40.150 215.460 40.325 ;
        RECT 214.545 39.850 215.460 40.150 ;
        RECT 215.630 40.110 215.870 40.510 ;
        RECT 216.040 40.450 216.210 40.680 ;
        RECT 216.380 40.620 216.570 41.060 ;
        RECT 216.740 40.610 217.690 40.890 ;
        RECT 217.910 40.700 218.260 40.870 ;
        RECT 216.040 40.280 216.570 40.450 ;
        RECT 214.545 39.820 215.285 39.850 ;
        RECT 212.460 39.140 213.415 39.360 ;
        RECT 212.690 38.510 212.960 38.970 ;
        RECT 213.130 38.680 213.415 39.140 ;
        RECT 213.700 38.510 213.990 39.675 ;
        RECT 214.165 38.820 214.420 39.700 ;
        RECT 214.590 38.510 214.895 39.650 ;
        RECT 215.115 39.230 215.285 39.820 ;
        RECT 215.630 39.740 216.170 40.110 ;
        RECT 216.350 40.000 216.570 40.280 ;
        RECT 216.740 39.830 216.910 40.610 ;
        RECT 216.505 39.660 216.910 39.830 ;
        RECT 217.080 39.820 217.430 40.440 ;
        RECT 216.505 39.570 216.675 39.660 ;
        RECT 217.600 39.650 217.810 40.440 ;
        RECT 215.455 39.400 216.675 39.570 ;
        RECT 217.135 39.490 217.810 39.650 ;
        RECT 215.115 39.060 215.915 39.230 ;
        RECT 215.235 38.510 215.565 38.890 ;
        RECT 215.745 38.770 215.915 39.060 ;
        RECT 216.505 39.020 216.675 39.400 ;
        RECT 216.845 39.480 217.810 39.490 ;
        RECT 218.000 40.310 218.260 40.700 ;
        RECT 218.470 40.600 218.800 41.060 ;
        RECT 219.675 40.670 220.530 40.840 ;
        RECT 220.735 40.670 221.230 40.840 ;
        RECT 221.400 40.700 221.730 41.060 ;
        RECT 218.000 39.620 218.170 40.310 ;
        RECT 218.340 39.960 218.510 40.140 ;
        RECT 218.680 40.130 219.470 40.380 ;
        RECT 219.675 39.960 219.845 40.670 ;
        RECT 220.015 40.160 220.370 40.380 ;
        RECT 218.340 39.790 220.030 39.960 ;
        RECT 216.845 39.190 217.305 39.480 ;
        RECT 218.000 39.450 219.500 39.620 ;
        RECT 218.000 39.310 218.170 39.450 ;
        RECT 217.610 39.140 218.170 39.310 ;
        RECT 216.085 38.510 216.335 38.970 ;
        RECT 216.505 38.680 217.375 39.020 ;
        RECT 217.610 38.680 217.780 39.140 ;
        RECT 218.615 39.110 219.690 39.280 ;
        RECT 217.950 38.510 218.320 38.970 ;
        RECT 218.615 38.770 218.785 39.110 ;
        RECT 218.955 38.510 219.285 38.940 ;
        RECT 219.520 38.770 219.690 39.110 ;
        RECT 219.860 39.010 220.030 39.790 ;
        RECT 220.200 39.570 220.370 40.160 ;
        RECT 220.540 39.760 220.890 40.380 ;
        RECT 220.200 39.180 220.665 39.570 ;
        RECT 221.060 39.310 221.230 40.670 ;
        RECT 221.400 39.480 221.860 40.530 ;
        RECT 220.835 39.140 221.230 39.310 ;
        RECT 220.835 39.010 221.005 39.140 ;
        RECT 219.860 38.680 220.540 39.010 ;
        RECT 220.755 38.680 221.005 39.010 ;
        RECT 221.175 38.510 221.425 38.970 ;
        RECT 221.595 38.695 221.920 39.480 ;
        RECT 222.090 38.680 222.260 40.800 ;
        RECT 222.430 40.680 222.760 41.060 ;
        RECT 222.930 40.510 223.185 40.800 ;
        RECT 222.435 40.340 223.185 40.510 ;
        RECT 222.435 39.350 222.665 40.340 ;
        RECT 223.360 40.290 225.030 41.060 ;
        RECT 222.835 39.520 223.185 40.170 ;
        RECT 223.360 39.770 224.110 40.290 ;
        RECT 225.475 40.250 225.720 40.855 ;
        RECT 225.940 40.525 226.450 41.060 ;
        RECT 224.280 39.600 225.030 40.120 ;
        RECT 222.435 39.180 223.185 39.350 ;
        RECT 222.430 38.510 222.760 39.010 ;
        RECT 222.930 38.680 223.185 39.180 ;
        RECT 223.360 38.510 225.030 39.600 ;
        RECT 225.200 40.080 226.430 40.250 ;
        RECT 225.200 39.270 225.540 40.080 ;
        RECT 225.710 39.515 226.460 39.705 ;
        RECT 225.200 38.860 225.715 39.270 ;
        RECT 225.950 38.510 226.120 39.270 ;
        RECT 226.290 38.850 226.460 39.515 ;
        RECT 226.630 39.530 226.820 40.890 ;
        RECT 226.990 40.720 227.265 40.890 ;
        RECT 226.990 40.550 227.270 40.720 ;
        RECT 226.990 39.730 227.265 40.550 ;
        RECT 227.455 40.525 227.985 40.890 ;
        RECT 228.410 40.660 228.740 41.060 ;
        RECT 227.810 40.490 227.985 40.525 ;
        RECT 227.470 39.530 227.640 40.330 ;
        RECT 226.630 39.360 227.640 39.530 ;
        RECT 227.810 40.320 228.740 40.490 ;
        RECT 228.910 40.320 229.165 40.890 ;
        RECT 227.810 39.190 227.980 40.320 ;
        RECT 228.570 40.150 228.740 40.320 ;
        RECT 226.855 39.020 227.980 39.190 ;
        RECT 228.150 39.820 228.345 40.150 ;
        RECT 228.570 39.820 228.825 40.150 ;
        RECT 228.150 38.850 228.320 39.820 ;
        RECT 228.995 39.650 229.165 40.320 ;
        RECT 226.290 38.680 228.320 38.850 ;
        RECT 228.490 38.510 228.660 39.650 ;
        RECT 228.830 38.680 229.165 39.650 ;
        RECT 229.345 40.320 229.600 40.890 ;
        RECT 229.770 40.660 230.100 41.060 ;
        RECT 230.525 40.525 231.055 40.890 ;
        RECT 230.525 40.490 230.700 40.525 ;
        RECT 229.770 40.320 230.700 40.490 ;
        RECT 231.245 40.380 231.520 40.890 ;
        RECT 229.345 39.650 229.515 40.320 ;
        RECT 229.770 40.150 229.940 40.320 ;
        RECT 229.685 39.820 229.940 40.150 ;
        RECT 230.165 39.820 230.360 40.150 ;
        RECT 229.345 38.680 229.680 39.650 ;
        RECT 229.850 38.510 230.020 39.650 ;
        RECT 230.190 38.850 230.360 39.820 ;
        RECT 230.530 39.190 230.700 40.320 ;
        RECT 230.870 39.530 231.040 40.330 ;
        RECT 231.240 40.210 231.520 40.380 ;
        RECT 231.245 39.730 231.520 40.210 ;
        RECT 231.690 39.530 231.880 40.890 ;
        RECT 232.060 40.525 232.570 41.060 ;
        RECT 232.790 40.250 233.035 40.855 ;
        RECT 233.945 40.320 234.200 40.890 ;
        RECT 234.370 40.660 234.700 41.060 ;
        RECT 235.125 40.525 235.655 40.890 ;
        RECT 235.125 40.490 235.300 40.525 ;
        RECT 234.370 40.320 235.300 40.490 ;
        RECT 235.845 40.380 236.120 40.890 ;
        RECT 232.080 40.080 233.310 40.250 ;
        RECT 230.870 39.360 231.880 39.530 ;
        RECT 232.050 39.515 232.800 39.705 ;
        RECT 230.530 39.020 231.655 39.190 ;
        RECT 232.050 38.850 232.220 39.515 ;
        RECT 232.970 39.270 233.310 40.080 ;
        RECT 230.190 38.680 232.220 38.850 ;
        RECT 232.390 38.510 232.560 39.270 ;
        RECT 232.795 38.860 233.310 39.270 ;
        RECT 233.945 39.650 234.115 40.320 ;
        RECT 234.370 40.150 234.540 40.320 ;
        RECT 234.285 39.820 234.540 40.150 ;
        RECT 234.765 39.820 234.960 40.150 ;
        RECT 233.945 38.680 234.280 39.650 ;
        RECT 234.450 38.510 234.620 39.650 ;
        RECT 234.790 38.850 234.960 39.820 ;
        RECT 235.130 39.190 235.300 40.320 ;
        RECT 235.470 39.530 235.640 40.330 ;
        RECT 235.840 40.210 236.120 40.380 ;
        RECT 235.845 39.730 236.120 40.210 ;
        RECT 236.290 39.530 236.480 40.890 ;
        RECT 236.660 40.525 237.170 41.060 ;
        RECT 237.390 40.250 237.635 40.855 ;
        RECT 238.080 40.310 239.290 41.060 ;
        RECT 239.460 40.335 239.750 41.060 ;
        RECT 239.955 40.320 240.570 40.890 ;
        RECT 240.740 40.550 240.955 41.060 ;
        RECT 241.185 40.550 241.465 40.880 ;
        RECT 241.645 40.550 241.885 41.060 ;
        RECT 236.680 40.080 237.910 40.250 ;
        RECT 235.470 39.360 236.480 39.530 ;
        RECT 236.650 39.515 237.400 39.705 ;
        RECT 235.130 39.020 236.255 39.190 ;
        RECT 236.650 38.850 236.820 39.515 ;
        RECT 237.570 39.270 237.910 40.080 ;
        RECT 238.080 39.770 238.600 40.310 ;
        RECT 238.770 39.600 239.290 40.140 ;
        RECT 234.790 38.680 236.820 38.850 ;
        RECT 236.990 38.510 237.160 39.270 ;
        RECT 237.395 38.860 237.910 39.270 ;
        RECT 238.080 38.510 239.290 39.600 ;
        RECT 239.460 38.510 239.750 39.675 ;
        RECT 239.955 39.300 240.270 40.320 ;
        RECT 240.440 39.650 240.610 40.150 ;
        RECT 240.860 39.820 241.125 40.380 ;
        RECT 241.295 39.650 241.465 40.550 ;
        RECT 241.635 39.820 241.990 40.380 ;
        RECT 242.225 40.320 242.480 40.890 ;
        RECT 242.650 40.660 242.980 41.060 ;
        RECT 243.405 40.525 243.935 40.890 ;
        RECT 244.125 40.720 244.400 40.890 ;
        RECT 244.120 40.550 244.400 40.720 ;
        RECT 243.405 40.490 243.580 40.525 ;
        RECT 242.650 40.320 243.580 40.490 ;
        RECT 242.225 39.650 242.395 40.320 ;
        RECT 242.650 40.150 242.820 40.320 ;
        RECT 242.565 39.820 242.820 40.150 ;
        RECT 243.045 39.820 243.240 40.150 ;
        RECT 240.440 39.480 241.865 39.650 ;
        RECT 239.955 38.680 240.490 39.300 ;
        RECT 240.660 38.510 240.990 39.310 ;
        RECT 241.475 39.305 241.865 39.480 ;
        RECT 242.225 38.680 242.560 39.650 ;
        RECT 242.730 38.510 242.900 39.650 ;
        RECT 243.070 38.850 243.240 39.820 ;
        RECT 243.410 39.190 243.580 40.320 ;
        RECT 243.750 39.530 243.920 40.330 ;
        RECT 244.125 39.730 244.400 40.550 ;
        RECT 244.570 39.530 244.760 40.890 ;
        RECT 244.940 40.525 245.450 41.060 ;
        RECT 245.670 40.250 245.915 40.855 ;
        RECT 246.365 40.320 246.620 40.890 ;
        RECT 246.790 40.660 247.120 41.060 ;
        RECT 247.545 40.525 248.075 40.890 ;
        RECT 247.545 40.490 247.720 40.525 ;
        RECT 246.790 40.320 247.720 40.490 ;
        RECT 244.960 40.080 246.190 40.250 ;
        RECT 243.750 39.360 244.760 39.530 ;
        RECT 244.930 39.515 245.680 39.705 ;
        RECT 243.410 39.020 244.535 39.190 ;
        RECT 244.930 38.850 245.100 39.515 ;
        RECT 245.850 39.270 246.190 40.080 ;
        RECT 243.070 38.680 245.100 38.850 ;
        RECT 245.270 38.510 245.440 39.270 ;
        RECT 245.675 38.860 246.190 39.270 ;
        RECT 246.365 39.650 246.535 40.320 ;
        RECT 246.790 40.150 246.960 40.320 ;
        RECT 246.705 39.820 246.960 40.150 ;
        RECT 247.185 39.820 247.380 40.150 ;
        RECT 246.365 38.680 246.700 39.650 ;
        RECT 246.870 38.510 247.040 39.650 ;
        RECT 247.210 38.850 247.380 39.820 ;
        RECT 247.550 39.190 247.720 40.320 ;
        RECT 247.890 39.530 248.060 40.330 ;
        RECT 248.265 40.040 248.540 40.890 ;
        RECT 248.260 39.870 248.540 40.040 ;
        RECT 248.265 39.730 248.540 39.870 ;
        RECT 248.710 39.530 248.900 40.890 ;
        RECT 249.080 40.525 249.590 41.060 ;
        RECT 249.810 40.250 250.055 40.855 ;
        RECT 250.500 40.320 250.885 40.890 ;
        RECT 251.055 40.600 251.380 41.060 ;
        RECT 251.900 40.430 252.180 40.890 ;
        RECT 249.100 40.080 250.330 40.250 ;
        RECT 247.890 39.360 248.900 39.530 ;
        RECT 249.070 39.515 249.820 39.705 ;
        RECT 247.550 39.020 248.675 39.190 ;
        RECT 249.070 38.850 249.240 39.515 ;
        RECT 249.990 39.270 250.330 40.080 ;
        RECT 247.210 38.680 249.240 38.850 ;
        RECT 249.410 38.510 249.580 39.270 ;
        RECT 249.815 38.860 250.330 39.270 ;
        RECT 250.500 39.650 250.780 40.320 ;
        RECT 251.055 40.260 252.180 40.430 ;
        RECT 251.055 40.150 251.505 40.260 ;
        RECT 250.950 39.820 251.505 40.150 ;
        RECT 252.370 40.090 252.770 40.890 ;
        RECT 253.170 40.600 253.440 41.060 ;
        RECT 253.610 40.430 253.895 40.890 ;
        RECT 250.500 38.680 250.885 39.650 ;
        RECT 251.055 39.360 251.505 39.820 ;
        RECT 251.675 39.530 252.770 40.090 ;
        RECT 251.055 39.140 252.180 39.360 ;
        RECT 251.055 38.510 251.380 38.970 ;
        RECT 251.900 38.680 252.180 39.140 ;
        RECT 252.370 38.680 252.770 39.530 ;
        RECT 252.940 40.260 253.895 40.430 ;
        RECT 254.180 40.290 255.850 41.060 ;
        RECT 252.940 39.360 253.150 40.260 ;
        RECT 253.320 39.530 254.010 40.090 ;
        RECT 254.180 39.770 254.930 40.290 ;
        RECT 256.490 40.250 256.760 41.060 ;
        RECT 256.930 40.250 257.260 40.890 ;
        RECT 257.430 40.250 257.670 41.060 ;
        RECT 255.100 39.600 255.850 40.120 ;
        RECT 256.480 39.820 256.830 40.070 ;
        RECT 257.000 39.650 257.170 40.250 ;
        RECT 257.865 40.240 258.140 41.060 ;
        RECT 258.310 40.420 258.640 40.890 ;
        RECT 258.810 40.590 258.980 41.060 ;
        RECT 259.150 40.420 259.480 40.890 ;
        RECT 259.650 40.590 259.820 41.060 ;
        RECT 259.990 40.420 260.320 40.890 ;
        RECT 260.490 40.590 260.660 41.060 ;
        RECT 260.830 40.420 261.160 40.890 ;
        RECT 261.330 40.590 261.615 41.060 ;
        RECT 258.310 40.240 261.830 40.420 ;
        RECT 257.340 39.820 257.690 40.070 ;
        RECT 257.915 39.870 259.575 40.070 ;
        RECT 259.895 39.870 261.260 40.070 ;
        RECT 261.430 39.700 261.830 40.240 ;
        RECT 252.940 39.140 253.895 39.360 ;
        RECT 253.170 38.510 253.440 38.970 ;
        RECT 253.610 38.680 253.895 39.140 ;
        RECT 254.180 38.510 255.850 39.600 ;
        RECT 256.490 38.510 256.820 39.650 ;
        RECT 257.000 39.480 257.680 39.650 ;
        RECT 257.350 38.695 257.680 39.480 ;
        RECT 257.865 39.480 259.900 39.690 ;
        RECT 257.865 38.680 258.140 39.480 ;
        RECT 258.310 38.510 258.640 39.310 ;
        RECT 258.810 38.680 258.980 39.480 ;
        RECT 259.150 38.510 259.400 39.310 ;
        RECT 259.570 38.850 259.900 39.480 ;
        RECT 260.070 39.400 261.830 39.700 ;
        RECT 262.000 40.115 262.340 40.890 ;
        RECT 262.510 40.600 262.680 41.060 ;
        RECT 262.920 40.625 263.280 40.890 ;
        RECT 262.920 40.620 263.275 40.625 ;
        RECT 262.920 40.610 263.270 40.620 ;
        RECT 262.920 40.605 263.265 40.610 ;
        RECT 262.920 40.595 263.260 40.605 ;
        RECT 263.910 40.600 264.080 41.060 ;
        RECT 262.920 40.590 263.255 40.595 ;
        RECT 262.920 40.580 263.245 40.590 ;
        RECT 262.920 40.570 263.235 40.580 ;
        RECT 262.920 40.430 263.220 40.570 ;
        RECT 262.510 40.240 263.220 40.430 ;
        RECT 263.410 40.430 263.740 40.510 ;
        RECT 264.250 40.430 264.590 40.890 ;
        RECT 263.410 40.240 264.590 40.430 ;
        RECT 265.220 40.335 265.510 41.060 ;
        RECT 265.680 40.320 266.065 40.890 ;
        RECT 266.235 40.600 266.560 41.060 ;
        RECT 267.080 40.430 267.360 40.890 ;
        RECT 260.070 39.020 260.240 39.400 ;
        RECT 260.410 38.850 260.740 39.210 ;
        RECT 260.910 39.020 261.080 39.400 ;
        RECT 261.250 38.850 261.665 39.230 ;
        RECT 259.570 38.680 261.665 38.850 ;
        RECT 262.000 38.680 262.280 40.115 ;
        RECT 262.510 39.670 262.795 40.240 ;
        RECT 262.980 39.840 263.450 40.070 ;
        RECT 263.620 40.050 263.950 40.070 ;
        RECT 263.620 39.870 264.070 40.050 ;
        RECT 264.260 39.870 264.590 40.070 ;
        RECT 262.510 39.455 263.660 39.670 ;
        RECT 262.450 38.510 263.160 39.285 ;
        RECT 263.330 38.680 263.660 39.455 ;
        RECT 263.855 38.755 264.070 39.870 ;
        RECT 264.360 39.530 264.590 39.870 ;
        RECT 264.250 38.510 264.580 39.230 ;
        RECT 265.220 38.510 265.510 39.675 ;
        RECT 265.680 39.650 265.960 40.320 ;
        RECT 266.235 40.260 267.360 40.430 ;
        RECT 266.235 40.150 266.685 40.260 ;
        RECT 266.130 39.820 266.685 40.150 ;
        RECT 267.550 40.090 267.950 40.890 ;
        RECT 268.350 40.600 268.620 41.060 ;
        RECT 268.790 40.430 269.075 40.890 ;
        RECT 270.350 40.660 270.680 41.060 ;
        RECT 270.850 40.490 271.020 40.760 ;
        RECT 271.190 40.660 271.520 41.060 ;
        RECT 271.690 40.490 271.945 40.760 ;
        RECT 265.680 38.680 266.065 39.650 ;
        RECT 266.235 39.360 266.685 39.820 ;
        RECT 266.855 39.530 267.950 40.090 ;
        RECT 266.235 39.140 267.360 39.360 ;
        RECT 266.235 38.510 266.560 38.970 ;
        RECT 267.080 38.680 267.360 39.140 ;
        RECT 267.550 38.680 267.950 39.530 ;
        RECT 268.120 40.260 269.075 40.430 ;
        RECT 268.120 39.360 268.330 40.260 ;
        RECT 268.500 39.530 269.190 40.090 ;
        RECT 270.280 39.480 270.550 40.490 ;
        RECT 270.720 40.320 271.945 40.490 ;
        RECT 272.125 40.350 272.380 40.880 ;
        RECT 272.550 40.600 272.855 41.060 ;
        RECT 273.100 40.680 274.170 40.850 ;
        RECT 270.720 39.650 270.890 40.320 ;
        RECT 271.060 39.820 271.440 40.150 ;
        RECT 271.610 39.820 271.945 40.150 ;
        RECT 270.720 39.480 271.035 39.650 ;
        RECT 268.120 39.140 269.075 39.360 ;
        RECT 268.350 38.510 268.620 38.970 ;
        RECT 268.790 38.680 269.075 39.140 ;
        RECT 270.285 38.510 270.600 39.310 ;
        RECT 270.865 38.865 271.035 39.480 ;
        RECT 271.205 39.140 271.440 39.820 ;
        RECT 272.125 39.700 272.335 40.350 ;
        RECT 273.100 40.325 273.420 40.680 ;
        RECT 273.095 40.150 273.420 40.325 ;
        RECT 272.505 39.850 273.420 40.150 ;
        RECT 273.590 40.110 273.830 40.510 ;
        RECT 274.000 40.450 274.170 40.680 ;
        RECT 274.340 40.620 274.530 41.060 ;
        RECT 274.700 40.610 275.650 40.890 ;
        RECT 275.870 40.700 276.220 40.870 ;
        RECT 274.000 40.280 274.530 40.450 ;
        RECT 272.505 39.820 273.245 39.850 ;
        RECT 271.610 38.865 271.945 39.650 ;
        RECT 270.865 38.695 271.945 38.865 ;
        RECT 272.125 38.820 272.380 39.700 ;
        RECT 272.550 38.510 272.855 39.650 ;
        RECT 273.075 39.230 273.245 39.820 ;
        RECT 273.590 39.740 274.130 40.110 ;
        RECT 274.310 40.000 274.530 40.280 ;
        RECT 274.700 39.830 274.870 40.610 ;
        RECT 274.465 39.660 274.870 39.830 ;
        RECT 275.040 39.820 275.390 40.440 ;
        RECT 274.465 39.570 274.635 39.660 ;
        RECT 275.560 39.650 275.770 40.440 ;
        RECT 273.415 39.400 274.635 39.570 ;
        RECT 275.095 39.490 275.770 39.650 ;
        RECT 273.075 39.060 273.875 39.230 ;
        RECT 273.195 38.510 273.525 38.890 ;
        RECT 273.705 38.770 273.875 39.060 ;
        RECT 274.465 39.020 274.635 39.400 ;
        RECT 274.805 39.480 275.770 39.490 ;
        RECT 275.960 40.310 276.220 40.700 ;
        RECT 276.430 40.600 276.760 41.060 ;
        RECT 277.635 40.670 278.490 40.840 ;
        RECT 278.695 40.670 279.190 40.840 ;
        RECT 279.360 40.700 279.690 41.060 ;
        RECT 275.960 39.620 276.130 40.310 ;
        RECT 276.300 39.960 276.470 40.140 ;
        RECT 276.640 40.130 277.430 40.380 ;
        RECT 277.635 39.960 277.805 40.670 ;
        RECT 277.975 40.160 278.330 40.380 ;
        RECT 276.300 39.790 277.990 39.960 ;
        RECT 274.805 39.190 275.265 39.480 ;
        RECT 275.960 39.450 277.460 39.620 ;
        RECT 275.960 39.310 276.130 39.450 ;
        RECT 275.570 39.140 276.130 39.310 ;
        RECT 274.045 38.510 274.295 38.970 ;
        RECT 274.465 38.680 275.335 39.020 ;
        RECT 275.570 38.680 275.740 39.140 ;
        RECT 276.575 39.110 277.650 39.280 ;
        RECT 275.910 38.510 276.280 38.970 ;
        RECT 276.575 38.770 276.745 39.110 ;
        RECT 276.915 38.510 277.245 38.940 ;
        RECT 277.480 38.770 277.650 39.110 ;
        RECT 277.820 39.010 277.990 39.790 ;
        RECT 278.160 39.570 278.330 40.160 ;
        RECT 278.500 39.760 278.850 40.380 ;
        RECT 278.160 39.180 278.625 39.570 ;
        RECT 279.020 39.310 279.190 40.670 ;
        RECT 279.360 39.480 279.820 40.530 ;
        RECT 278.795 39.140 279.190 39.310 ;
        RECT 278.795 39.010 278.965 39.140 ;
        RECT 277.820 38.680 278.500 39.010 ;
        RECT 278.715 38.680 278.965 39.010 ;
        RECT 279.135 38.510 279.385 38.970 ;
        RECT 279.555 38.695 279.880 39.480 ;
        RECT 280.050 38.680 280.220 40.800 ;
        RECT 280.390 40.680 280.720 41.060 ;
        RECT 280.890 40.510 281.145 40.800 ;
        RECT 280.395 40.340 281.145 40.510 ;
        RECT 281.325 40.350 281.580 40.880 ;
        RECT 281.750 40.600 282.055 41.060 ;
        RECT 282.300 40.680 283.370 40.850 ;
        RECT 280.395 39.350 280.625 40.340 ;
        RECT 280.795 39.520 281.145 40.170 ;
        RECT 281.325 39.700 281.535 40.350 ;
        RECT 282.300 40.325 282.620 40.680 ;
        RECT 282.295 40.150 282.620 40.325 ;
        RECT 281.705 39.850 282.620 40.150 ;
        RECT 282.790 40.110 283.030 40.510 ;
        RECT 283.200 40.450 283.370 40.680 ;
        RECT 283.540 40.620 283.730 41.060 ;
        RECT 283.900 40.610 284.850 40.890 ;
        RECT 285.070 40.700 285.420 40.870 ;
        RECT 283.200 40.280 283.730 40.450 ;
        RECT 281.705 39.820 282.445 39.850 ;
        RECT 280.395 39.180 281.145 39.350 ;
        RECT 280.390 38.510 280.720 39.010 ;
        RECT 280.890 38.680 281.145 39.180 ;
        RECT 281.325 38.820 281.580 39.700 ;
        RECT 281.750 38.510 282.055 39.650 ;
        RECT 282.275 39.230 282.445 39.820 ;
        RECT 282.790 39.740 283.330 40.110 ;
        RECT 283.510 40.000 283.730 40.280 ;
        RECT 283.900 39.830 284.070 40.610 ;
        RECT 283.665 39.660 284.070 39.830 ;
        RECT 284.240 39.820 284.590 40.440 ;
        RECT 283.665 39.570 283.835 39.660 ;
        RECT 284.760 39.650 284.970 40.440 ;
        RECT 282.615 39.400 283.835 39.570 ;
        RECT 284.295 39.490 284.970 39.650 ;
        RECT 282.275 39.060 283.075 39.230 ;
        RECT 282.395 38.510 282.725 38.890 ;
        RECT 282.905 38.770 283.075 39.060 ;
        RECT 283.665 39.020 283.835 39.400 ;
        RECT 284.005 39.480 284.970 39.490 ;
        RECT 285.160 40.310 285.420 40.700 ;
        RECT 285.630 40.600 285.960 41.060 ;
        RECT 286.835 40.670 287.690 40.840 ;
        RECT 287.895 40.670 288.390 40.840 ;
        RECT 288.560 40.700 288.890 41.060 ;
        RECT 285.160 39.620 285.330 40.310 ;
        RECT 285.500 39.960 285.670 40.140 ;
        RECT 285.840 40.130 286.630 40.380 ;
        RECT 286.835 39.960 287.005 40.670 ;
        RECT 287.175 40.160 287.530 40.380 ;
        RECT 285.500 39.790 287.190 39.960 ;
        RECT 284.005 39.190 284.465 39.480 ;
        RECT 285.160 39.450 286.660 39.620 ;
        RECT 285.160 39.310 285.330 39.450 ;
        RECT 284.770 39.140 285.330 39.310 ;
        RECT 283.245 38.510 283.495 38.970 ;
        RECT 283.665 38.680 284.535 39.020 ;
        RECT 284.770 38.680 284.940 39.140 ;
        RECT 285.775 39.110 286.850 39.280 ;
        RECT 285.110 38.510 285.480 38.970 ;
        RECT 285.775 38.770 285.945 39.110 ;
        RECT 286.115 38.510 286.445 38.940 ;
        RECT 286.680 38.770 286.850 39.110 ;
        RECT 287.020 39.010 287.190 39.790 ;
        RECT 287.360 39.570 287.530 40.160 ;
        RECT 287.700 39.760 288.050 40.380 ;
        RECT 287.360 39.180 287.825 39.570 ;
        RECT 288.220 39.310 288.390 40.670 ;
        RECT 288.560 39.480 289.020 40.530 ;
        RECT 287.995 39.140 288.390 39.310 ;
        RECT 287.995 39.010 288.165 39.140 ;
        RECT 287.020 38.680 287.700 39.010 ;
        RECT 287.915 38.680 288.165 39.010 ;
        RECT 288.335 38.510 288.585 38.970 ;
        RECT 288.755 38.695 289.080 39.480 ;
        RECT 289.250 38.680 289.420 40.800 ;
        RECT 289.590 40.680 289.920 41.060 ;
        RECT 290.090 40.510 290.345 40.800 ;
        RECT 289.595 40.340 290.345 40.510 ;
        RECT 289.595 39.350 289.825 40.340 ;
        RECT 290.980 40.335 291.270 41.060 ;
        RECT 291.440 40.515 296.785 41.060 ;
        RECT 289.995 39.520 290.345 40.170 ;
        RECT 293.025 39.685 293.365 40.515 ;
        RECT 297.885 40.510 298.140 40.800 ;
        RECT 298.310 40.680 298.640 41.060 ;
        RECT 297.885 40.340 298.635 40.510 ;
        RECT 289.595 39.180 290.345 39.350 ;
        RECT 289.590 38.510 289.920 39.010 ;
        RECT 290.090 38.680 290.345 39.180 ;
        RECT 290.980 38.510 291.270 39.675 ;
        RECT 294.845 38.945 295.195 40.195 ;
        RECT 297.885 39.520 298.235 40.170 ;
        RECT 298.405 39.350 298.635 40.340 ;
        RECT 297.885 39.180 298.635 39.350 ;
        RECT 291.440 38.510 296.785 38.945 ;
        RECT 297.885 38.680 298.140 39.180 ;
        RECT 298.310 38.510 298.640 39.010 ;
        RECT 298.810 38.680 298.980 40.800 ;
        RECT 299.340 40.700 299.670 41.060 ;
        RECT 299.840 40.670 300.335 40.840 ;
        RECT 300.540 40.670 301.395 40.840 ;
        RECT 299.210 39.480 299.670 40.530 ;
        RECT 299.150 38.695 299.475 39.480 ;
        RECT 299.840 39.310 300.010 40.670 ;
        RECT 300.180 39.760 300.530 40.380 ;
        RECT 300.700 40.160 301.055 40.380 ;
        RECT 300.700 39.570 300.870 40.160 ;
        RECT 301.225 39.960 301.395 40.670 ;
        RECT 302.270 40.600 302.600 41.060 ;
        RECT 302.810 40.700 303.160 40.870 ;
        RECT 301.600 40.130 302.390 40.380 ;
        RECT 302.810 40.310 303.070 40.700 ;
        RECT 303.380 40.610 304.330 40.890 ;
        RECT 304.500 40.620 304.690 41.060 ;
        RECT 304.860 40.680 305.930 40.850 ;
        RECT 302.560 39.960 302.730 40.140 ;
        RECT 299.840 39.140 300.235 39.310 ;
        RECT 300.405 39.180 300.870 39.570 ;
        RECT 301.040 39.790 302.730 39.960 ;
        RECT 300.065 39.010 300.235 39.140 ;
        RECT 301.040 39.010 301.210 39.790 ;
        RECT 302.900 39.620 303.070 40.310 ;
        RECT 301.570 39.450 303.070 39.620 ;
        RECT 303.260 39.650 303.470 40.440 ;
        RECT 303.640 39.820 303.990 40.440 ;
        RECT 304.160 39.830 304.330 40.610 ;
        RECT 304.860 40.450 305.030 40.680 ;
        RECT 304.500 40.280 305.030 40.450 ;
        RECT 304.500 40.000 304.720 40.280 ;
        RECT 305.200 40.110 305.440 40.510 ;
        RECT 304.160 39.660 304.565 39.830 ;
        RECT 304.900 39.740 305.440 40.110 ;
        RECT 305.610 40.325 305.930 40.680 ;
        RECT 306.175 40.600 306.480 41.060 ;
        RECT 306.650 40.350 306.905 40.880 ;
        RECT 305.610 40.150 305.935 40.325 ;
        RECT 305.610 39.850 306.525 40.150 ;
        RECT 305.785 39.820 306.525 39.850 ;
        RECT 303.260 39.490 303.935 39.650 ;
        RECT 304.395 39.570 304.565 39.660 ;
        RECT 303.260 39.480 304.225 39.490 ;
        RECT 302.900 39.310 303.070 39.450 ;
        RECT 299.645 38.510 299.895 38.970 ;
        RECT 300.065 38.680 300.315 39.010 ;
        RECT 300.530 38.680 301.210 39.010 ;
        RECT 301.380 39.110 302.455 39.280 ;
        RECT 302.900 39.140 303.460 39.310 ;
        RECT 303.765 39.190 304.225 39.480 ;
        RECT 304.395 39.400 305.615 39.570 ;
        RECT 301.380 38.770 301.550 39.110 ;
        RECT 301.785 38.510 302.115 38.940 ;
        RECT 302.285 38.770 302.455 39.110 ;
        RECT 302.750 38.510 303.120 38.970 ;
        RECT 303.290 38.680 303.460 39.140 ;
        RECT 304.395 39.020 304.565 39.400 ;
        RECT 305.785 39.230 305.955 39.820 ;
        RECT 306.695 39.700 306.905 40.350 ;
        RECT 307.170 40.510 307.340 40.890 ;
        RECT 307.555 40.680 307.885 41.060 ;
        RECT 307.170 40.340 307.885 40.510 ;
        RECT 307.080 39.790 307.435 40.160 ;
        RECT 307.715 40.150 307.885 40.340 ;
        RECT 308.055 40.315 308.310 40.890 ;
        RECT 307.715 39.820 307.970 40.150 ;
        RECT 303.695 38.680 304.565 39.020 ;
        RECT 305.155 39.060 305.955 39.230 ;
        RECT 304.735 38.510 304.985 38.970 ;
        RECT 305.155 38.770 305.325 39.060 ;
        RECT 305.505 38.510 305.835 38.890 ;
        RECT 306.175 38.510 306.480 39.650 ;
        RECT 306.650 38.820 306.905 39.700 ;
        RECT 307.715 39.610 307.885 39.820 ;
        RECT 307.170 39.440 307.885 39.610 ;
        RECT 308.140 39.585 308.310 40.315 ;
        RECT 308.485 40.220 308.745 41.060 ;
        RECT 309.840 40.310 311.050 41.060 ;
        RECT 307.170 38.680 307.340 39.440 ;
        RECT 307.555 38.510 307.885 39.270 ;
        RECT 308.055 38.680 308.310 39.585 ;
        RECT 308.485 38.510 308.745 39.660 ;
        RECT 309.840 39.600 310.360 40.140 ;
        RECT 310.530 39.770 311.050 40.310 ;
        RECT 309.840 38.510 311.050 39.600 ;
        RECT 162.095 38.340 311.135 38.510 ;
        RECT 162.180 37.250 163.390 38.340 ;
        RECT 163.560 37.250 167.070 38.340 ;
        RECT 167.815 37.710 168.100 38.170 ;
        RECT 168.270 37.880 168.540 38.340 ;
        RECT 167.815 37.490 168.770 37.710 ;
        RECT 162.180 36.540 162.700 37.080 ;
        RECT 162.870 36.710 163.390 37.250 ;
        RECT 163.560 36.560 165.210 37.080 ;
        RECT 165.380 36.730 167.070 37.250 ;
        RECT 167.700 36.760 168.390 37.320 ;
        RECT 168.560 36.590 168.770 37.490 ;
        RECT 162.180 35.790 163.390 36.540 ;
        RECT 163.560 35.790 167.070 36.560 ;
        RECT 167.815 36.420 168.770 36.590 ;
        RECT 168.940 37.320 169.340 38.170 ;
        RECT 169.530 37.710 169.810 38.170 ;
        RECT 170.330 37.880 170.655 38.340 ;
        RECT 169.530 37.490 170.655 37.710 ;
        RECT 168.940 36.760 170.035 37.320 ;
        RECT 170.205 37.030 170.655 37.490 ;
        RECT 170.825 37.200 171.210 38.170 ;
        RECT 171.495 37.710 171.780 38.170 ;
        RECT 171.950 37.880 172.220 38.340 ;
        RECT 171.495 37.490 172.450 37.710 ;
        RECT 167.815 35.960 168.100 36.420 ;
        RECT 168.270 35.790 168.540 36.250 ;
        RECT 168.940 35.960 169.340 36.760 ;
        RECT 170.205 36.700 170.760 37.030 ;
        RECT 170.205 36.590 170.655 36.700 ;
        RECT 169.530 36.420 170.655 36.590 ;
        RECT 170.930 36.530 171.210 37.200 ;
        RECT 171.380 36.760 172.070 37.320 ;
        RECT 172.240 36.590 172.450 37.490 ;
        RECT 169.530 35.960 169.810 36.420 ;
        RECT 170.330 35.790 170.655 36.250 ;
        RECT 170.825 35.960 171.210 36.530 ;
        RECT 171.495 36.420 172.450 36.590 ;
        RECT 172.620 37.320 173.020 38.170 ;
        RECT 173.210 37.710 173.490 38.170 ;
        RECT 174.010 37.880 174.335 38.340 ;
        RECT 173.210 37.490 174.335 37.710 ;
        RECT 172.620 36.760 173.715 37.320 ;
        RECT 173.885 37.030 174.335 37.490 ;
        RECT 174.505 37.200 174.890 38.170 ;
        RECT 171.495 35.960 171.780 36.420 ;
        RECT 171.950 35.790 172.220 36.250 ;
        RECT 172.620 35.960 173.020 36.760 ;
        RECT 173.885 36.700 174.440 37.030 ;
        RECT 173.885 36.590 174.335 36.700 ;
        RECT 173.210 36.420 174.335 36.590 ;
        RECT 174.610 36.530 174.890 37.200 ;
        RECT 175.060 37.175 175.350 38.340 ;
        RECT 175.525 37.200 175.860 38.170 ;
        RECT 176.030 37.200 176.200 38.340 ;
        RECT 176.370 38.000 178.400 38.170 ;
        RECT 173.210 35.960 173.490 36.420 ;
        RECT 174.010 35.790 174.335 36.250 ;
        RECT 174.505 35.960 174.890 36.530 ;
        RECT 175.525 36.530 175.695 37.200 ;
        RECT 176.370 37.030 176.540 38.000 ;
        RECT 175.865 36.700 176.120 37.030 ;
        RECT 176.345 36.700 176.540 37.030 ;
        RECT 176.710 37.660 177.835 37.830 ;
        RECT 175.950 36.530 176.120 36.700 ;
        RECT 176.710 36.530 176.880 37.660 ;
        RECT 175.060 35.790 175.350 36.515 ;
        RECT 175.525 35.960 175.780 36.530 ;
        RECT 175.950 36.360 176.880 36.530 ;
        RECT 177.050 37.320 178.060 37.490 ;
        RECT 177.050 36.520 177.220 37.320 ;
        RECT 177.425 36.640 177.700 37.120 ;
        RECT 177.420 36.470 177.700 36.640 ;
        RECT 176.705 36.325 176.880 36.360 ;
        RECT 175.950 35.790 176.280 36.190 ;
        RECT 176.705 35.960 177.235 36.325 ;
        RECT 177.425 35.960 177.700 36.470 ;
        RECT 177.870 35.960 178.060 37.320 ;
        RECT 178.230 37.335 178.400 38.000 ;
        RECT 178.570 37.580 178.740 38.340 ;
        RECT 178.975 37.580 179.490 37.990 ;
        RECT 178.230 37.145 178.980 37.335 ;
        RECT 179.150 36.770 179.490 37.580 ;
        RECT 179.660 37.250 181.330 38.340 ;
        RECT 182.075 37.710 182.360 38.170 ;
        RECT 182.530 37.880 182.800 38.340 ;
        RECT 182.075 37.490 183.030 37.710 ;
        RECT 178.260 36.600 179.490 36.770 ;
        RECT 178.240 35.790 178.750 36.325 ;
        RECT 178.970 35.995 179.215 36.600 ;
        RECT 179.660 36.560 180.410 37.080 ;
        RECT 180.580 36.730 181.330 37.250 ;
        RECT 181.960 36.760 182.650 37.320 ;
        RECT 182.820 36.590 183.030 37.490 ;
        RECT 179.660 35.790 181.330 36.560 ;
        RECT 182.075 36.420 183.030 36.590 ;
        RECT 183.200 37.320 183.600 38.170 ;
        RECT 183.790 37.710 184.070 38.170 ;
        RECT 184.590 37.880 184.915 38.340 ;
        RECT 183.790 37.490 184.915 37.710 ;
        RECT 183.200 36.760 184.295 37.320 ;
        RECT 184.465 37.030 184.915 37.490 ;
        RECT 185.085 37.200 185.470 38.170 ;
        RECT 182.075 35.960 182.360 36.420 ;
        RECT 182.530 35.790 182.800 36.250 ;
        RECT 183.200 35.960 183.600 36.760 ;
        RECT 184.465 36.700 185.020 37.030 ;
        RECT 184.465 36.590 184.915 36.700 ;
        RECT 183.790 36.420 184.915 36.590 ;
        RECT 185.190 36.530 185.470 37.200 ;
        RECT 183.790 35.960 184.070 36.420 ;
        RECT 184.590 35.790 184.915 36.250 ;
        RECT 185.085 35.960 185.470 36.530 ;
        RECT 185.645 37.150 185.900 38.030 ;
        RECT 186.070 37.200 186.375 38.340 ;
        RECT 186.715 37.960 187.045 38.340 ;
        RECT 187.225 37.790 187.395 38.080 ;
        RECT 187.565 37.880 187.815 38.340 ;
        RECT 186.595 37.620 187.395 37.790 ;
        RECT 187.985 37.830 188.855 38.170 ;
        RECT 185.645 36.500 185.855 37.150 ;
        RECT 186.595 37.030 186.765 37.620 ;
        RECT 187.985 37.450 188.155 37.830 ;
        RECT 189.090 37.710 189.260 38.170 ;
        RECT 189.430 37.880 189.800 38.340 ;
        RECT 190.095 37.740 190.265 38.080 ;
        RECT 190.435 37.910 190.765 38.340 ;
        RECT 191.000 37.740 191.170 38.080 ;
        RECT 186.935 37.280 188.155 37.450 ;
        RECT 188.325 37.370 188.785 37.660 ;
        RECT 189.090 37.540 189.650 37.710 ;
        RECT 190.095 37.570 191.170 37.740 ;
        RECT 191.340 37.840 192.020 38.170 ;
        RECT 192.235 37.840 192.485 38.170 ;
        RECT 192.655 37.880 192.905 38.340 ;
        RECT 189.480 37.400 189.650 37.540 ;
        RECT 188.325 37.360 189.290 37.370 ;
        RECT 187.985 37.190 188.155 37.280 ;
        RECT 188.615 37.200 189.290 37.360 ;
        RECT 186.025 37.000 186.765 37.030 ;
        RECT 186.025 36.700 186.940 37.000 ;
        RECT 186.615 36.525 186.940 36.700 ;
        RECT 185.645 35.970 185.900 36.500 ;
        RECT 186.070 35.790 186.375 36.250 ;
        RECT 186.620 36.170 186.940 36.525 ;
        RECT 187.110 36.740 187.650 37.110 ;
        RECT 187.985 37.020 188.390 37.190 ;
        RECT 187.110 36.340 187.350 36.740 ;
        RECT 187.830 36.570 188.050 36.850 ;
        RECT 187.520 36.400 188.050 36.570 ;
        RECT 187.520 36.170 187.690 36.400 ;
        RECT 188.220 36.240 188.390 37.020 ;
        RECT 188.560 36.410 188.910 37.030 ;
        RECT 189.080 36.410 189.290 37.200 ;
        RECT 189.480 37.230 190.980 37.400 ;
        RECT 189.480 36.540 189.650 37.230 ;
        RECT 191.340 37.060 191.510 37.840 ;
        RECT 192.315 37.710 192.485 37.840 ;
        RECT 189.820 36.890 191.510 37.060 ;
        RECT 191.680 37.280 192.145 37.670 ;
        RECT 192.315 37.540 192.710 37.710 ;
        RECT 189.820 36.710 189.990 36.890 ;
        RECT 186.620 36.000 187.690 36.170 ;
        RECT 187.860 35.790 188.050 36.230 ;
        RECT 188.220 35.960 189.170 36.240 ;
        RECT 189.480 36.150 189.740 36.540 ;
        RECT 190.160 36.470 190.950 36.720 ;
        RECT 189.390 35.980 189.740 36.150 ;
        RECT 189.950 35.790 190.280 36.250 ;
        RECT 191.155 36.180 191.325 36.890 ;
        RECT 191.680 36.690 191.850 37.280 ;
        RECT 191.495 36.470 191.850 36.690 ;
        RECT 192.020 36.470 192.370 37.090 ;
        RECT 192.540 36.180 192.710 37.540 ;
        RECT 193.075 37.370 193.400 38.155 ;
        RECT 192.880 36.320 193.340 37.370 ;
        RECT 191.155 36.010 192.010 36.180 ;
        RECT 192.215 36.010 192.710 36.180 ;
        RECT 192.880 35.790 193.210 36.150 ;
        RECT 193.570 36.050 193.740 38.170 ;
        RECT 193.910 37.840 194.240 38.340 ;
        RECT 194.410 37.670 194.665 38.170 ;
        RECT 193.915 37.500 194.665 37.670 ;
        RECT 194.955 37.710 195.240 38.170 ;
        RECT 195.410 37.880 195.680 38.340 ;
        RECT 193.915 36.510 194.145 37.500 ;
        RECT 194.955 37.490 195.910 37.710 ;
        RECT 194.315 36.680 194.665 37.330 ;
        RECT 194.840 36.760 195.530 37.320 ;
        RECT 195.700 36.590 195.910 37.490 ;
        RECT 193.915 36.340 194.665 36.510 ;
        RECT 193.910 35.790 194.240 36.170 ;
        RECT 194.410 36.050 194.665 36.340 ;
        RECT 194.955 36.420 195.910 36.590 ;
        RECT 196.080 37.320 196.480 38.170 ;
        RECT 196.670 37.710 196.950 38.170 ;
        RECT 197.470 37.880 197.795 38.340 ;
        RECT 196.670 37.490 197.795 37.710 ;
        RECT 196.080 36.760 197.175 37.320 ;
        RECT 197.345 37.030 197.795 37.490 ;
        RECT 197.965 37.200 198.350 38.170 ;
        RECT 198.520 37.250 200.190 38.340 ;
        RECT 194.955 35.960 195.240 36.420 ;
        RECT 195.410 35.790 195.680 36.250 ;
        RECT 196.080 35.960 196.480 36.760 ;
        RECT 197.345 36.700 197.900 37.030 ;
        RECT 197.345 36.590 197.795 36.700 ;
        RECT 196.670 36.420 197.795 36.590 ;
        RECT 198.070 36.530 198.350 37.200 ;
        RECT 196.670 35.960 196.950 36.420 ;
        RECT 197.470 35.790 197.795 36.250 ;
        RECT 197.965 35.960 198.350 36.530 ;
        RECT 198.520 36.560 199.270 37.080 ;
        RECT 199.440 36.730 200.190 37.250 ;
        RECT 200.820 37.175 201.110 38.340 ;
        RECT 201.280 37.250 202.950 38.340 ;
        RECT 201.280 36.560 202.030 37.080 ;
        RECT 202.200 36.730 202.950 37.250 ;
        RECT 203.585 37.200 203.920 38.170 ;
        RECT 204.090 37.200 204.260 38.340 ;
        RECT 204.430 38.000 206.460 38.170 ;
        RECT 198.520 35.790 200.190 36.560 ;
        RECT 200.820 35.790 201.110 36.515 ;
        RECT 201.280 35.790 202.950 36.560 ;
        RECT 203.585 36.530 203.755 37.200 ;
        RECT 204.430 37.030 204.600 38.000 ;
        RECT 203.925 36.700 204.180 37.030 ;
        RECT 204.405 36.700 204.600 37.030 ;
        RECT 204.770 37.660 205.895 37.830 ;
        RECT 204.010 36.530 204.180 36.700 ;
        RECT 204.770 36.530 204.940 37.660 ;
        RECT 203.585 35.960 203.840 36.530 ;
        RECT 204.010 36.360 204.940 36.530 ;
        RECT 205.110 37.320 206.120 37.490 ;
        RECT 205.110 36.520 205.280 37.320 ;
        RECT 205.485 36.980 205.760 37.120 ;
        RECT 205.480 36.810 205.760 36.980 ;
        RECT 204.765 36.325 204.940 36.360 ;
        RECT 204.010 35.790 204.340 36.190 ;
        RECT 204.765 35.960 205.295 36.325 ;
        RECT 205.485 35.960 205.760 36.810 ;
        RECT 205.930 35.960 206.120 37.320 ;
        RECT 206.290 37.335 206.460 38.000 ;
        RECT 206.630 37.580 206.800 38.340 ;
        RECT 207.035 37.580 207.550 37.990 ;
        RECT 206.290 37.145 207.040 37.335 ;
        RECT 207.210 36.770 207.550 37.580 ;
        RECT 206.320 36.600 207.550 36.770 ;
        RECT 207.720 37.200 208.105 38.170 ;
        RECT 208.275 37.880 208.600 38.340 ;
        RECT 209.120 37.710 209.400 38.170 ;
        RECT 208.275 37.490 209.400 37.710 ;
        RECT 206.300 35.790 206.810 36.325 ;
        RECT 207.030 35.995 207.275 36.600 ;
        RECT 207.720 36.530 208.000 37.200 ;
        RECT 208.275 37.030 208.725 37.490 ;
        RECT 209.590 37.320 209.990 38.170 ;
        RECT 210.390 37.880 210.660 38.340 ;
        RECT 210.830 37.710 211.115 38.170 ;
        RECT 208.170 36.700 208.725 37.030 ;
        RECT 208.895 36.760 209.990 37.320 ;
        RECT 208.275 36.590 208.725 36.700 ;
        RECT 207.720 35.960 208.105 36.530 ;
        RECT 208.275 36.420 209.400 36.590 ;
        RECT 208.275 35.790 208.600 36.250 ;
        RECT 209.120 35.960 209.400 36.420 ;
        RECT 209.590 35.960 209.990 36.760 ;
        RECT 210.160 37.490 211.115 37.710 ;
        RECT 210.160 36.590 210.370 37.490 ;
        RECT 211.455 37.470 211.740 38.340 ;
        RECT 211.910 37.710 212.170 38.170 ;
        RECT 212.345 37.880 212.600 38.340 ;
        RECT 212.770 37.710 213.030 38.170 ;
        RECT 211.910 37.540 213.030 37.710 ;
        RECT 213.200 37.540 213.510 38.340 ;
        RECT 210.540 36.760 211.230 37.320 ;
        RECT 211.910 37.290 212.170 37.540 ;
        RECT 213.680 37.370 213.990 38.170 ;
        RECT 211.415 37.120 212.170 37.290 ;
        RECT 212.960 37.200 213.990 37.370 ;
        RECT 211.415 36.610 211.820 37.120 ;
        RECT 212.960 36.950 213.130 37.200 ;
        RECT 211.990 36.780 213.130 36.950 ;
        RECT 210.160 36.420 211.115 36.590 ;
        RECT 211.415 36.440 213.065 36.610 ;
        RECT 213.300 36.460 213.650 37.030 ;
        RECT 210.390 35.790 210.660 36.250 ;
        RECT 210.830 35.960 211.115 36.420 ;
        RECT 211.460 35.790 211.740 36.270 ;
        RECT 211.910 36.050 212.170 36.440 ;
        RECT 212.345 35.790 212.600 36.270 ;
        RECT 212.770 36.050 213.065 36.440 ;
        RECT 213.820 36.290 213.990 37.200 ;
        RECT 214.620 37.580 215.135 37.990 ;
        RECT 215.370 37.580 215.540 38.340 ;
        RECT 215.710 38.000 217.740 38.170 ;
        RECT 214.620 36.770 214.960 37.580 ;
        RECT 215.710 37.335 215.880 38.000 ;
        RECT 216.275 37.660 217.400 37.830 ;
        RECT 215.130 37.145 215.880 37.335 ;
        RECT 216.050 37.320 217.060 37.490 ;
        RECT 214.620 36.600 215.850 36.770 ;
        RECT 213.245 35.790 213.520 36.270 ;
        RECT 213.690 35.960 213.990 36.290 ;
        RECT 214.895 35.995 215.140 36.600 ;
        RECT 215.360 35.790 215.870 36.325 ;
        RECT 216.050 35.960 216.240 37.320 ;
        RECT 216.410 36.980 216.685 37.120 ;
        RECT 216.410 36.810 216.690 36.980 ;
        RECT 216.410 35.960 216.685 36.810 ;
        RECT 216.890 36.520 217.060 37.320 ;
        RECT 217.230 36.530 217.400 37.660 ;
        RECT 217.570 37.030 217.740 38.000 ;
        RECT 217.910 37.200 218.080 38.340 ;
        RECT 218.250 37.200 218.585 38.170 ;
        RECT 219.335 37.710 219.620 38.170 ;
        RECT 219.790 37.880 220.060 38.340 ;
        RECT 219.335 37.490 220.290 37.710 ;
        RECT 217.570 36.700 217.765 37.030 ;
        RECT 217.990 36.700 218.245 37.030 ;
        RECT 217.990 36.530 218.160 36.700 ;
        RECT 218.415 36.530 218.585 37.200 ;
        RECT 219.220 36.760 219.910 37.320 ;
        RECT 220.080 36.590 220.290 37.490 ;
        RECT 217.230 36.360 218.160 36.530 ;
        RECT 217.230 36.325 217.405 36.360 ;
        RECT 216.875 35.960 217.405 36.325 ;
        RECT 217.830 35.790 218.160 36.190 ;
        RECT 218.330 35.960 218.585 36.530 ;
        RECT 219.335 36.420 220.290 36.590 ;
        RECT 220.460 37.320 220.860 38.170 ;
        RECT 221.050 37.710 221.330 38.170 ;
        RECT 221.850 37.880 222.175 38.340 ;
        RECT 221.050 37.490 222.175 37.710 ;
        RECT 220.460 36.760 221.555 37.320 ;
        RECT 221.725 37.030 222.175 37.490 ;
        RECT 222.345 37.200 222.730 38.170 ;
        RECT 223.015 37.710 223.300 38.170 ;
        RECT 223.470 37.880 223.740 38.340 ;
        RECT 223.015 37.490 223.970 37.710 ;
        RECT 219.335 35.960 219.620 36.420 ;
        RECT 219.790 35.790 220.060 36.250 ;
        RECT 220.460 35.960 220.860 36.760 ;
        RECT 221.725 36.700 222.280 37.030 ;
        RECT 221.725 36.590 222.175 36.700 ;
        RECT 221.050 36.420 222.175 36.590 ;
        RECT 222.450 36.530 222.730 37.200 ;
        RECT 222.900 36.760 223.590 37.320 ;
        RECT 223.760 36.590 223.970 37.490 ;
        RECT 221.050 35.960 221.330 36.420 ;
        RECT 221.850 35.790 222.175 36.250 ;
        RECT 222.345 35.960 222.730 36.530 ;
        RECT 223.015 36.420 223.970 36.590 ;
        RECT 224.140 37.320 224.540 38.170 ;
        RECT 224.730 37.710 225.010 38.170 ;
        RECT 225.530 37.880 225.855 38.340 ;
        RECT 224.730 37.490 225.855 37.710 ;
        RECT 224.140 36.760 225.235 37.320 ;
        RECT 225.405 37.030 225.855 37.490 ;
        RECT 226.025 37.200 226.410 38.170 ;
        RECT 223.015 35.960 223.300 36.420 ;
        RECT 223.470 35.790 223.740 36.250 ;
        RECT 224.140 35.960 224.540 36.760 ;
        RECT 225.405 36.700 225.960 37.030 ;
        RECT 225.405 36.590 225.855 36.700 ;
        RECT 224.730 36.420 225.855 36.590 ;
        RECT 226.130 36.530 226.410 37.200 ;
        RECT 226.580 37.175 226.870 38.340 ;
        RECT 227.040 37.250 229.630 38.340 ;
        RECT 230.265 37.670 230.520 38.170 ;
        RECT 230.690 37.840 231.020 38.340 ;
        RECT 230.265 37.500 231.015 37.670 ;
        RECT 224.730 35.960 225.010 36.420 ;
        RECT 225.530 35.790 225.855 36.250 ;
        RECT 226.025 35.960 226.410 36.530 ;
        RECT 227.040 36.560 228.250 37.080 ;
        RECT 228.420 36.730 229.630 37.250 ;
        RECT 230.265 36.680 230.615 37.330 ;
        RECT 226.580 35.790 226.870 36.515 ;
        RECT 227.040 35.790 229.630 36.560 ;
        RECT 230.785 36.510 231.015 37.500 ;
        RECT 230.265 36.340 231.015 36.510 ;
        RECT 230.265 36.050 230.520 36.340 ;
        RECT 230.690 35.790 231.020 36.170 ;
        RECT 231.190 36.050 231.360 38.170 ;
        RECT 231.530 37.370 231.855 38.155 ;
        RECT 232.025 37.880 232.275 38.340 ;
        RECT 232.445 37.840 232.695 38.170 ;
        RECT 232.910 37.840 233.590 38.170 ;
        RECT 232.445 37.710 232.615 37.840 ;
        RECT 232.220 37.540 232.615 37.710 ;
        RECT 231.590 36.320 232.050 37.370 ;
        RECT 232.220 36.180 232.390 37.540 ;
        RECT 232.785 37.280 233.250 37.670 ;
        RECT 232.560 36.470 232.910 37.090 ;
        RECT 233.080 36.690 233.250 37.280 ;
        RECT 233.420 37.060 233.590 37.840 ;
        RECT 233.760 37.740 233.930 38.080 ;
        RECT 234.165 37.910 234.495 38.340 ;
        RECT 234.665 37.740 234.835 38.080 ;
        RECT 235.130 37.880 235.500 38.340 ;
        RECT 233.760 37.570 234.835 37.740 ;
        RECT 235.670 37.710 235.840 38.170 ;
        RECT 236.075 37.830 236.945 38.170 ;
        RECT 237.115 37.880 237.365 38.340 ;
        RECT 235.280 37.540 235.840 37.710 ;
        RECT 235.280 37.400 235.450 37.540 ;
        RECT 233.950 37.230 235.450 37.400 ;
        RECT 236.145 37.370 236.605 37.660 ;
        RECT 233.420 36.890 235.110 37.060 ;
        RECT 233.080 36.470 233.435 36.690 ;
        RECT 233.605 36.180 233.775 36.890 ;
        RECT 233.980 36.470 234.770 36.720 ;
        RECT 234.940 36.710 235.110 36.890 ;
        RECT 235.280 36.540 235.450 37.230 ;
        RECT 231.720 35.790 232.050 36.150 ;
        RECT 232.220 36.010 232.715 36.180 ;
        RECT 232.920 36.010 233.775 36.180 ;
        RECT 234.650 35.790 234.980 36.250 ;
        RECT 235.190 36.150 235.450 36.540 ;
        RECT 235.640 37.360 236.605 37.370 ;
        RECT 236.775 37.450 236.945 37.830 ;
        RECT 237.535 37.790 237.705 38.080 ;
        RECT 237.885 37.960 238.215 38.340 ;
        RECT 237.535 37.620 238.335 37.790 ;
        RECT 235.640 37.200 236.315 37.360 ;
        RECT 236.775 37.280 237.995 37.450 ;
        RECT 235.640 36.410 235.850 37.200 ;
        RECT 236.775 37.190 236.945 37.280 ;
        RECT 236.020 36.410 236.370 37.030 ;
        RECT 236.540 37.020 236.945 37.190 ;
        RECT 236.540 36.240 236.710 37.020 ;
        RECT 236.880 36.570 237.100 36.850 ;
        RECT 237.280 36.740 237.820 37.110 ;
        RECT 238.165 37.030 238.335 37.620 ;
        RECT 238.555 37.200 238.860 38.340 ;
        RECT 239.030 37.150 239.280 38.030 ;
        RECT 239.450 37.200 239.700 38.340 ;
        RECT 240.845 37.670 241.100 38.170 ;
        RECT 241.270 37.840 241.600 38.340 ;
        RECT 240.845 37.500 241.595 37.670 ;
        RECT 238.165 37.000 238.905 37.030 ;
        RECT 236.880 36.400 237.410 36.570 ;
        RECT 235.190 35.980 235.540 36.150 ;
        RECT 235.760 35.960 236.710 36.240 ;
        RECT 236.880 35.790 237.070 36.230 ;
        RECT 237.240 36.170 237.410 36.400 ;
        RECT 237.580 36.340 237.820 36.740 ;
        RECT 237.990 36.700 238.905 37.000 ;
        RECT 237.990 36.525 238.315 36.700 ;
        RECT 237.990 36.170 238.310 36.525 ;
        RECT 239.075 36.500 239.280 37.150 ;
        RECT 240.845 36.680 241.195 37.330 ;
        RECT 237.240 36.000 238.310 36.170 ;
        RECT 238.555 35.790 238.860 36.250 ;
        RECT 239.030 35.970 239.280 36.500 ;
        RECT 239.450 35.790 239.700 36.545 ;
        RECT 241.365 36.510 241.595 37.500 ;
        RECT 240.845 36.340 241.595 36.510 ;
        RECT 240.845 36.050 241.100 36.340 ;
        RECT 241.270 35.790 241.600 36.170 ;
        RECT 241.770 36.050 241.940 38.170 ;
        RECT 242.110 37.370 242.435 38.155 ;
        RECT 242.605 37.880 242.855 38.340 ;
        RECT 243.025 37.840 243.275 38.170 ;
        RECT 243.490 37.840 244.170 38.170 ;
        RECT 243.025 37.710 243.195 37.840 ;
        RECT 242.800 37.540 243.195 37.710 ;
        RECT 242.170 36.320 242.630 37.370 ;
        RECT 242.800 36.180 242.970 37.540 ;
        RECT 243.365 37.280 243.830 37.670 ;
        RECT 243.140 36.470 243.490 37.090 ;
        RECT 243.660 36.690 243.830 37.280 ;
        RECT 244.000 37.060 244.170 37.840 ;
        RECT 244.340 37.740 244.510 38.080 ;
        RECT 244.745 37.910 245.075 38.340 ;
        RECT 245.245 37.740 245.415 38.080 ;
        RECT 245.710 37.880 246.080 38.340 ;
        RECT 244.340 37.570 245.415 37.740 ;
        RECT 246.250 37.710 246.420 38.170 ;
        RECT 246.655 37.830 247.525 38.170 ;
        RECT 247.695 37.880 247.945 38.340 ;
        RECT 245.860 37.540 246.420 37.710 ;
        RECT 245.860 37.400 246.030 37.540 ;
        RECT 244.530 37.230 246.030 37.400 ;
        RECT 246.725 37.370 247.185 37.660 ;
        RECT 244.000 36.890 245.690 37.060 ;
        RECT 243.660 36.470 244.015 36.690 ;
        RECT 244.185 36.180 244.355 36.890 ;
        RECT 244.560 36.470 245.350 36.720 ;
        RECT 245.520 36.710 245.690 36.890 ;
        RECT 245.860 36.540 246.030 37.230 ;
        RECT 242.300 35.790 242.630 36.150 ;
        RECT 242.800 36.010 243.295 36.180 ;
        RECT 243.500 36.010 244.355 36.180 ;
        RECT 245.230 35.790 245.560 36.250 ;
        RECT 245.770 36.150 246.030 36.540 ;
        RECT 246.220 37.360 247.185 37.370 ;
        RECT 247.355 37.450 247.525 37.830 ;
        RECT 248.115 37.790 248.285 38.080 ;
        RECT 248.465 37.960 248.795 38.340 ;
        RECT 248.115 37.620 248.915 37.790 ;
        RECT 246.220 37.200 246.895 37.360 ;
        RECT 247.355 37.280 248.575 37.450 ;
        RECT 246.220 36.410 246.430 37.200 ;
        RECT 247.355 37.190 247.525 37.280 ;
        RECT 246.600 36.410 246.950 37.030 ;
        RECT 247.120 37.020 247.525 37.190 ;
        RECT 247.120 36.240 247.290 37.020 ;
        RECT 247.460 36.570 247.680 36.850 ;
        RECT 247.860 36.740 248.400 37.110 ;
        RECT 248.745 37.030 248.915 37.620 ;
        RECT 249.135 37.200 249.440 38.340 ;
        RECT 249.610 37.150 249.865 38.030 ;
        RECT 250.040 37.250 251.710 38.340 ;
        RECT 248.745 37.000 249.485 37.030 ;
        RECT 247.460 36.400 247.990 36.570 ;
        RECT 245.770 35.980 246.120 36.150 ;
        RECT 246.340 35.960 247.290 36.240 ;
        RECT 247.460 35.790 247.650 36.230 ;
        RECT 247.820 36.170 247.990 36.400 ;
        RECT 248.160 36.340 248.400 36.740 ;
        RECT 248.570 36.700 249.485 37.000 ;
        RECT 248.570 36.525 248.895 36.700 ;
        RECT 248.570 36.170 248.890 36.525 ;
        RECT 249.655 36.500 249.865 37.150 ;
        RECT 247.820 36.000 248.890 36.170 ;
        RECT 249.135 35.790 249.440 36.250 ;
        RECT 249.610 35.970 249.865 36.500 ;
        RECT 250.040 36.560 250.790 37.080 ;
        RECT 250.960 36.730 251.710 37.250 ;
        RECT 252.340 37.175 252.630 38.340 ;
        RECT 252.800 37.250 254.470 38.340 ;
        RECT 252.800 36.560 253.550 37.080 ;
        RECT 253.720 36.730 254.470 37.250 ;
        RECT 255.105 37.150 255.360 38.030 ;
        RECT 255.530 37.200 255.835 38.340 ;
        RECT 256.175 37.960 256.505 38.340 ;
        RECT 256.685 37.790 256.855 38.080 ;
        RECT 257.025 37.880 257.275 38.340 ;
        RECT 256.055 37.620 256.855 37.790 ;
        RECT 257.445 37.830 258.315 38.170 ;
        RECT 250.040 35.790 251.710 36.560 ;
        RECT 252.340 35.790 252.630 36.515 ;
        RECT 252.800 35.790 254.470 36.560 ;
        RECT 255.105 36.500 255.315 37.150 ;
        RECT 256.055 37.030 256.225 37.620 ;
        RECT 257.445 37.450 257.615 37.830 ;
        RECT 258.550 37.710 258.720 38.170 ;
        RECT 258.890 37.880 259.260 38.340 ;
        RECT 259.555 37.740 259.725 38.080 ;
        RECT 259.895 37.910 260.225 38.340 ;
        RECT 260.460 37.740 260.630 38.080 ;
        RECT 256.395 37.280 257.615 37.450 ;
        RECT 257.785 37.370 258.245 37.660 ;
        RECT 258.550 37.540 259.110 37.710 ;
        RECT 259.555 37.570 260.630 37.740 ;
        RECT 260.800 37.840 261.480 38.170 ;
        RECT 261.695 37.840 261.945 38.170 ;
        RECT 262.115 37.880 262.365 38.340 ;
        RECT 258.940 37.400 259.110 37.540 ;
        RECT 257.785 37.360 258.750 37.370 ;
        RECT 257.445 37.190 257.615 37.280 ;
        RECT 258.075 37.200 258.750 37.360 ;
        RECT 255.485 37.000 256.225 37.030 ;
        RECT 255.485 36.700 256.400 37.000 ;
        RECT 256.075 36.525 256.400 36.700 ;
        RECT 255.105 35.970 255.360 36.500 ;
        RECT 255.530 35.790 255.835 36.250 ;
        RECT 256.080 36.170 256.400 36.525 ;
        RECT 256.570 36.740 257.110 37.110 ;
        RECT 257.445 37.020 257.850 37.190 ;
        RECT 256.570 36.340 256.810 36.740 ;
        RECT 257.290 36.570 257.510 36.850 ;
        RECT 256.980 36.400 257.510 36.570 ;
        RECT 256.980 36.170 257.150 36.400 ;
        RECT 257.680 36.240 257.850 37.020 ;
        RECT 258.020 36.410 258.370 37.030 ;
        RECT 258.540 36.410 258.750 37.200 ;
        RECT 258.940 37.230 260.440 37.400 ;
        RECT 258.940 36.540 259.110 37.230 ;
        RECT 260.800 37.060 260.970 37.840 ;
        RECT 261.775 37.710 261.945 37.840 ;
        RECT 259.280 36.890 260.970 37.060 ;
        RECT 261.140 37.280 261.605 37.670 ;
        RECT 261.775 37.540 262.170 37.710 ;
        RECT 259.280 36.710 259.450 36.890 ;
        RECT 256.080 36.000 257.150 36.170 ;
        RECT 257.320 35.790 257.510 36.230 ;
        RECT 257.680 35.960 258.630 36.240 ;
        RECT 258.940 36.150 259.200 36.540 ;
        RECT 259.620 36.470 260.410 36.720 ;
        RECT 258.850 35.980 259.200 36.150 ;
        RECT 259.410 35.790 259.740 36.250 ;
        RECT 260.615 36.180 260.785 36.890 ;
        RECT 261.140 36.690 261.310 37.280 ;
        RECT 260.955 36.470 261.310 36.690 ;
        RECT 261.480 36.470 261.830 37.090 ;
        RECT 262.000 36.180 262.170 37.540 ;
        RECT 262.535 37.370 262.860 38.155 ;
        RECT 262.340 36.320 262.800 37.370 ;
        RECT 260.615 36.010 261.470 36.180 ;
        RECT 261.675 36.010 262.170 36.180 ;
        RECT 262.340 35.790 262.670 36.150 ;
        RECT 263.030 36.050 263.200 38.170 ;
        RECT 263.370 37.840 263.700 38.340 ;
        RECT 263.870 37.670 264.125 38.170 ;
        RECT 263.375 37.500 264.125 37.670 ;
        RECT 263.375 36.510 263.605 37.500 ;
        RECT 264.300 37.370 264.610 38.170 ;
        RECT 264.780 37.540 265.090 38.340 ;
        RECT 265.260 37.710 265.520 38.170 ;
        RECT 265.690 37.880 265.945 38.340 ;
        RECT 266.120 37.710 266.380 38.170 ;
        RECT 265.260 37.540 266.380 37.710 ;
        RECT 263.775 36.680 264.125 37.330 ;
        RECT 264.300 37.200 265.330 37.370 ;
        RECT 263.375 36.340 264.125 36.510 ;
        RECT 263.370 35.790 263.700 36.170 ;
        RECT 263.870 36.050 264.125 36.340 ;
        RECT 264.300 36.290 264.470 37.200 ;
        RECT 264.640 36.460 264.990 37.030 ;
        RECT 265.160 36.950 265.330 37.200 ;
        RECT 266.120 37.290 266.380 37.540 ;
        RECT 266.550 37.470 266.835 38.340 ;
        RECT 267.060 37.470 267.335 38.170 ;
        RECT 267.505 37.795 267.760 38.340 ;
        RECT 267.930 37.830 268.410 38.170 ;
        RECT 268.585 37.785 269.190 38.340 ;
        RECT 268.575 37.685 269.190 37.785 ;
        RECT 268.575 37.660 268.760 37.685 ;
        RECT 266.120 37.120 266.875 37.290 ;
        RECT 265.160 36.780 266.300 36.950 ;
        RECT 266.470 36.610 266.875 37.120 ;
        RECT 265.225 36.440 266.875 36.610 ;
        RECT 267.060 36.440 267.230 37.470 ;
        RECT 267.505 37.340 268.260 37.590 ;
        RECT 268.430 37.415 268.760 37.660 ;
        RECT 267.505 37.305 268.275 37.340 ;
        RECT 267.505 37.295 268.290 37.305 ;
        RECT 267.400 37.280 268.295 37.295 ;
        RECT 267.400 37.265 268.315 37.280 ;
        RECT 267.400 37.255 268.335 37.265 ;
        RECT 267.400 37.245 268.360 37.255 ;
        RECT 267.400 37.215 268.430 37.245 ;
        RECT 267.400 37.185 268.450 37.215 ;
        RECT 267.400 37.155 268.470 37.185 ;
        RECT 267.400 37.130 268.500 37.155 ;
        RECT 267.400 37.095 268.535 37.130 ;
        RECT 267.400 37.090 268.565 37.095 ;
        RECT 267.400 36.695 267.630 37.090 ;
        RECT 268.175 37.085 268.565 37.090 ;
        RECT 268.200 37.075 268.565 37.085 ;
        RECT 268.215 37.070 268.565 37.075 ;
        RECT 268.230 37.065 268.565 37.070 ;
        RECT 268.930 37.065 269.190 37.515 ;
        RECT 269.360 37.250 272.870 38.340 ;
        RECT 268.230 37.060 269.190 37.065 ;
        RECT 268.240 37.050 269.190 37.060 ;
        RECT 268.250 37.045 269.190 37.050 ;
        RECT 268.260 37.035 269.190 37.045 ;
        RECT 268.265 37.025 269.190 37.035 ;
        RECT 268.270 37.020 269.190 37.025 ;
        RECT 268.280 37.005 269.190 37.020 ;
        RECT 268.285 36.990 269.190 37.005 ;
        RECT 268.295 36.965 269.190 36.990 ;
        RECT 267.800 36.495 268.130 36.920 ;
        RECT 267.880 36.470 268.130 36.495 ;
        RECT 264.300 35.960 264.600 36.290 ;
        RECT 264.770 35.790 265.045 36.270 ;
        RECT 265.225 36.050 265.520 36.440 ;
        RECT 265.690 35.790 265.945 36.270 ;
        RECT 266.120 36.050 266.380 36.440 ;
        RECT 266.550 35.790 266.830 36.270 ;
        RECT 267.060 35.960 267.320 36.440 ;
        RECT 267.490 35.790 267.740 36.330 ;
        RECT 267.910 36.010 268.130 36.470 ;
        RECT 268.300 36.895 269.190 36.965 ;
        RECT 268.300 36.170 268.470 36.895 ;
        RECT 268.640 36.340 269.190 36.725 ;
        RECT 269.360 36.560 271.010 37.080 ;
        RECT 271.180 36.730 272.870 37.250 ;
        RECT 273.960 37.915 274.495 38.130 ;
        RECT 275.420 37.915 275.760 38.340 ;
        RECT 276.265 37.915 276.595 38.340 ;
        RECT 277.105 37.915 277.465 38.340 ;
        RECT 268.300 36.000 269.190 36.170 ;
        RECT 269.360 35.790 272.870 36.560 ;
        RECT 273.960 36.530 274.165 37.915 ;
        RECT 277.670 37.745 277.930 37.925 ;
        RECT 274.395 37.575 277.930 37.745 ;
        RECT 274.395 37.030 274.625 37.575 ;
        RECT 277.250 37.515 277.930 37.575 ;
        RECT 274.335 36.700 274.625 37.030 ;
        RECT 274.815 36.700 275.125 37.405 ;
        RECT 275.295 37.120 275.615 37.405 ;
        RECT 275.795 37.120 277.080 37.405 ;
        RECT 275.295 36.700 275.480 37.120 ;
        RECT 275.650 36.780 276.740 36.950 ;
        RECT 275.650 36.595 275.820 36.780 ;
        RECT 276.910 36.610 277.080 37.120 ;
        RECT 275.615 36.530 275.820 36.595 ;
        RECT 273.960 36.425 275.820 36.530 ;
        RECT 275.990 36.440 277.080 36.610 ;
        RECT 277.250 36.610 277.420 37.515 ;
        RECT 277.590 36.780 277.930 37.345 ;
        RECT 278.100 37.175 278.390 38.340 ;
        RECT 278.560 37.200 278.945 38.170 ;
        RECT 279.115 37.880 279.440 38.340 ;
        RECT 279.960 37.710 280.240 38.170 ;
        RECT 279.115 37.490 280.240 37.710 ;
        RECT 277.250 36.440 277.930 36.610 ;
        RECT 278.560 36.530 278.840 37.200 ;
        RECT 279.115 37.030 279.565 37.490 ;
        RECT 280.430 37.320 280.830 38.170 ;
        RECT 281.230 37.880 281.500 38.340 ;
        RECT 281.670 37.710 281.955 38.170 ;
        RECT 279.010 36.700 279.565 37.030 ;
        RECT 279.735 36.760 280.830 37.320 ;
        RECT 279.115 36.590 279.565 36.700 ;
        RECT 273.960 36.360 275.765 36.425 ;
        RECT 273.960 36.310 274.355 36.360 ;
        RECT 274.100 36.010 274.355 36.310 ;
        RECT 274.525 35.790 274.915 36.190 ;
        RECT 275.085 36.010 275.255 36.360 ;
        RECT 275.990 36.290 276.160 36.440 ;
        RECT 275.425 35.790 275.755 36.190 ;
        RECT 275.925 35.960 276.160 36.290 ;
        RECT 276.345 35.790 276.515 36.270 ;
        RECT 276.685 35.990 277.015 36.440 ;
        RECT 277.225 35.790 277.395 36.270 ;
        RECT 277.670 35.995 277.930 36.440 ;
        RECT 278.100 35.790 278.390 36.515 ;
        RECT 278.560 35.960 278.945 36.530 ;
        RECT 279.115 36.420 280.240 36.590 ;
        RECT 279.115 35.790 279.440 36.250 ;
        RECT 279.960 35.960 280.240 36.420 ;
        RECT 280.430 35.960 280.830 36.760 ;
        RECT 281.000 37.490 281.955 37.710 ;
        RECT 281.000 36.590 281.210 37.490 ;
        RECT 282.240 37.470 282.515 38.170 ;
        RECT 282.725 37.795 282.940 38.340 ;
        RECT 283.110 37.830 283.585 38.170 ;
        RECT 283.755 37.835 284.370 38.340 ;
        RECT 283.755 37.660 283.950 37.835 ;
        RECT 281.380 36.760 282.070 37.320 ;
        RECT 281.000 36.420 281.955 36.590 ;
        RECT 281.230 35.790 281.500 36.250 ;
        RECT 281.670 35.960 281.955 36.420 ;
        RECT 282.240 36.440 282.410 37.470 ;
        RECT 282.685 37.300 283.400 37.595 ;
        RECT 283.620 37.470 283.950 37.660 ;
        RECT 284.120 37.300 284.370 37.665 ;
        RECT 282.580 37.130 284.370 37.300 ;
        RECT 282.580 36.700 282.810 37.130 ;
        RECT 282.240 35.960 282.500 36.440 ;
        RECT 282.980 36.430 283.390 36.950 ;
        RECT 282.670 35.790 283.000 36.250 ;
        RECT 283.190 36.010 283.390 36.430 ;
        RECT 283.560 36.275 283.815 37.130 ;
        RECT 284.610 36.950 284.780 38.170 ;
        RECT 285.030 37.830 285.290 38.340 ;
        RECT 285.460 37.905 290.805 38.340 ;
        RECT 290.980 37.905 296.325 38.340 ;
        RECT 296.500 37.905 301.845 38.340 ;
        RECT 283.985 36.700 284.780 36.950 ;
        RECT 284.950 36.780 285.290 37.660 ;
        RECT 284.530 36.610 284.780 36.700 ;
        RECT 283.560 36.010 284.350 36.275 ;
        RECT 284.530 36.190 284.860 36.610 ;
        RECT 285.030 35.790 285.290 36.610 ;
        RECT 287.045 36.335 287.385 37.165 ;
        RECT 288.865 36.655 289.215 37.905 ;
        RECT 292.565 36.335 292.905 37.165 ;
        RECT 294.385 36.655 294.735 37.905 ;
        RECT 298.085 36.335 298.425 37.165 ;
        RECT 299.905 36.655 300.255 37.905 ;
        RECT 302.020 37.250 303.690 38.340 ;
        RECT 302.020 36.560 302.770 37.080 ;
        RECT 302.940 36.730 303.690 37.250 ;
        RECT 303.860 37.175 304.150 38.340 ;
        RECT 304.870 37.410 305.040 38.170 ;
        RECT 305.220 37.580 305.550 38.340 ;
        RECT 304.870 37.240 305.535 37.410 ;
        RECT 305.720 37.265 305.990 38.170 ;
        RECT 306.275 37.710 306.560 38.170 ;
        RECT 306.730 37.880 307.000 38.340 ;
        RECT 306.275 37.490 307.230 37.710 ;
        RECT 305.365 37.095 305.535 37.240 ;
        RECT 304.800 36.690 305.130 37.060 ;
        RECT 305.365 36.765 305.650 37.095 ;
        RECT 285.460 35.790 290.805 36.335 ;
        RECT 290.980 35.790 296.325 36.335 ;
        RECT 296.500 35.790 301.845 36.335 ;
        RECT 302.020 35.790 303.690 36.560 ;
        RECT 303.860 35.790 304.150 36.515 ;
        RECT 305.365 36.510 305.535 36.765 ;
        RECT 304.870 36.340 305.535 36.510 ;
        RECT 305.820 36.465 305.990 37.265 ;
        RECT 306.160 36.760 306.850 37.320 ;
        RECT 307.020 36.590 307.230 37.490 ;
        RECT 304.870 35.960 305.040 36.340 ;
        RECT 305.220 35.790 305.550 36.170 ;
        RECT 305.730 35.960 305.990 36.465 ;
        RECT 306.275 36.420 307.230 36.590 ;
        RECT 307.400 37.320 307.800 38.170 ;
        RECT 307.990 37.710 308.270 38.170 ;
        RECT 308.790 37.880 309.115 38.340 ;
        RECT 307.990 37.490 309.115 37.710 ;
        RECT 307.400 36.760 308.495 37.320 ;
        RECT 308.665 37.030 309.115 37.490 ;
        RECT 309.285 37.200 309.670 38.170 ;
        RECT 306.275 35.960 306.560 36.420 ;
        RECT 306.730 35.790 307.000 36.250 ;
        RECT 307.400 35.960 307.800 36.760 ;
        RECT 308.665 36.700 309.220 37.030 ;
        RECT 308.665 36.590 309.115 36.700 ;
        RECT 307.990 36.420 309.115 36.590 ;
        RECT 309.390 36.530 309.670 37.200 ;
        RECT 309.840 37.250 311.050 38.340 ;
        RECT 309.840 36.710 310.360 37.250 ;
        RECT 310.530 36.540 311.050 37.080 ;
        RECT 307.990 35.960 308.270 36.420 ;
        RECT 308.790 35.790 309.115 36.250 ;
        RECT 309.285 35.960 309.670 36.530 ;
        RECT 309.840 35.790 311.050 36.540 ;
        RECT 162.095 35.620 311.135 35.790 ;
        RECT 162.180 34.870 163.390 35.620 ;
        RECT 162.180 34.330 162.700 34.870 ;
        RECT 163.560 34.850 165.230 35.620 ;
        RECT 165.865 34.910 166.120 35.440 ;
        RECT 166.290 35.160 166.595 35.620 ;
        RECT 166.840 35.240 167.910 35.410 ;
        RECT 162.870 34.160 163.390 34.700 ;
        RECT 163.560 34.330 164.310 34.850 ;
        RECT 164.480 34.160 165.230 34.680 ;
        RECT 162.180 33.070 163.390 34.160 ;
        RECT 163.560 33.070 165.230 34.160 ;
        RECT 165.865 34.260 166.075 34.910 ;
        RECT 166.840 34.885 167.160 35.240 ;
        RECT 166.835 34.710 167.160 34.885 ;
        RECT 166.245 34.410 167.160 34.710 ;
        RECT 167.330 34.670 167.570 35.070 ;
        RECT 167.740 35.010 167.910 35.240 ;
        RECT 168.080 35.180 168.270 35.620 ;
        RECT 168.440 35.170 169.390 35.450 ;
        RECT 169.610 35.260 169.960 35.430 ;
        RECT 167.740 34.840 168.270 35.010 ;
        RECT 166.245 34.380 166.985 34.410 ;
        RECT 165.865 33.380 166.120 34.260 ;
        RECT 166.290 33.070 166.595 34.210 ;
        RECT 166.815 33.790 166.985 34.380 ;
        RECT 167.330 34.300 167.870 34.670 ;
        RECT 168.050 34.560 168.270 34.840 ;
        RECT 168.440 34.390 168.610 35.170 ;
        RECT 168.205 34.220 168.610 34.390 ;
        RECT 168.780 34.380 169.130 35.000 ;
        RECT 168.205 34.130 168.375 34.220 ;
        RECT 169.300 34.210 169.510 35.000 ;
        RECT 167.155 33.960 168.375 34.130 ;
        RECT 168.835 34.050 169.510 34.210 ;
        RECT 166.815 33.620 167.615 33.790 ;
        RECT 166.935 33.070 167.265 33.450 ;
        RECT 167.445 33.330 167.615 33.620 ;
        RECT 168.205 33.580 168.375 33.960 ;
        RECT 168.545 34.040 169.510 34.050 ;
        RECT 169.700 34.870 169.960 35.260 ;
        RECT 170.170 35.160 170.500 35.620 ;
        RECT 171.375 35.230 172.230 35.400 ;
        RECT 172.435 35.230 172.930 35.400 ;
        RECT 173.100 35.260 173.430 35.620 ;
        RECT 169.700 34.180 169.870 34.870 ;
        RECT 170.040 34.520 170.210 34.700 ;
        RECT 170.380 34.690 171.170 34.940 ;
        RECT 171.375 34.520 171.545 35.230 ;
        RECT 171.715 34.720 172.070 34.940 ;
        RECT 170.040 34.350 171.730 34.520 ;
        RECT 168.545 33.750 169.005 34.040 ;
        RECT 169.700 34.010 171.200 34.180 ;
        RECT 169.700 33.870 169.870 34.010 ;
        RECT 169.310 33.700 169.870 33.870 ;
        RECT 167.785 33.070 168.035 33.530 ;
        RECT 168.205 33.240 169.075 33.580 ;
        RECT 169.310 33.240 169.480 33.700 ;
        RECT 170.315 33.670 171.390 33.840 ;
        RECT 169.650 33.070 170.020 33.530 ;
        RECT 170.315 33.330 170.485 33.670 ;
        RECT 170.655 33.070 170.985 33.500 ;
        RECT 171.220 33.330 171.390 33.670 ;
        RECT 171.560 33.570 171.730 34.350 ;
        RECT 171.900 34.130 172.070 34.720 ;
        RECT 172.240 34.320 172.590 34.940 ;
        RECT 171.900 33.740 172.365 34.130 ;
        RECT 172.760 33.870 172.930 35.230 ;
        RECT 173.100 34.040 173.560 35.090 ;
        RECT 172.535 33.700 172.930 33.870 ;
        RECT 172.535 33.570 172.705 33.700 ;
        RECT 171.560 33.240 172.240 33.570 ;
        RECT 172.455 33.240 172.705 33.570 ;
        RECT 172.875 33.070 173.125 33.530 ;
        RECT 173.295 33.255 173.620 34.040 ;
        RECT 173.790 33.240 173.960 35.360 ;
        RECT 174.130 35.240 174.460 35.620 ;
        RECT 174.630 35.070 174.885 35.360 ;
        RECT 174.135 34.900 174.885 35.070 ;
        RECT 174.135 33.910 174.365 34.900 ;
        RECT 175.065 34.880 175.320 35.450 ;
        RECT 175.490 35.220 175.820 35.620 ;
        RECT 176.245 35.085 176.775 35.450 ;
        RECT 176.245 35.050 176.420 35.085 ;
        RECT 175.490 34.880 176.420 35.050 ;
        RECT 174.535 34.080 174.885 34.730 ;
        RECT 175.065 34.210 175.235 34.880 ;
        RECT 175.490 34.710 175.660 34.880 ;
        RECT 175.405 34.380 175.660 34.710 ;
        RECT 175.885 34.380 176.080 34.710 ;
        RECT 174.135 33.740 174.885 33.910 ;
        RECT 174.130 33.070 174.460 33.570 ;
        RECT 174.630 33.240 174.885 33.740 ;
        RECT 175.065 33.240 175.400 34.210 ;
        RECT 175.570 33.070 175.740 34.210 ;
        RECT 175.910 33.410 176.080 34.380 ;
        RECT 176.250 33.750 176.420 34.880 ;
        RECT 176.590 34.090 176.760 34.890 ;
        RECT 176.965 34.600 177.240 35.450 ;
        RECT 176.960 34.430 177.240 34.600 ;
        RECT 176.965 34.290 177.240 34.430 ;
        RECT 177.410 34.090 177.600 35.450 ;
        RECT 177.780 35.085 178.290 35.620 ;
        RECT 178.510 34.810 178.755 35.415 ;
        RECT 179.935 34.810 180.180 35.415 ;
        RECT 180.400 35.085 180.910 35.620 ;
        RECT 177.800 34.640 179.030 34.810 ;
        RECT 176.590 33.920 177.600 34.090 ;
        RECT 177.770 34.075 178.520 34.265 ;
        RECT 176.250 33.580 177.375 33.750 ;
        RECT 177.770 33.410 177.940 34.075 ;
        RECT 178.690 33.830 179.030 34.640 ;
        RECT 175.910 33.240 177.940 33.410 ;
        RECT 178.110 33.070 178.280 33.830 ;
        RECT 178.515 33.420 179.030 33.830 ;
        RECT 179.660 34.640 180.890 34.810 ;
        RECT 179.660 33.830 180.000 34.640 ;
        RECT 180.170 34.075 180.920 34.265 ;
        RECT 179.660 33.420 180.175 33.830 ;
        RECT 180.410 33.070 180.580 33.830 ;
        RECT 180.750 33.410 180.920 34.075 ;
        RECT 181.090 34.090 181.280 35.450 ;
        RECT 181.450 34.940 181.725 35.450 ;
        RECT 181.915 35.085 182.445 35.450 ;
        RECT 182.870 35.220 183.200 35.620 ;
        RECT 182.270 35.050 182.445 35.085 ;
        RECT 181.450 34.770 181.730 34.940 ;
        RECT 181.450 34.290 181.725 34.770 ;
        RECT 181.930 34.090 182.100 34.890 ;
        RECT 181.090 33.920 182.100 34.090 ;
        RECT 182.270 34.880 183.200 35.050 ;
        RECT 183.370 34.880 183.625 35.450 ;
        RECT 182.270 33.750 182.440 34.880 ;
        RECT 183.030 34.710 183.200 34.880 ;
        RECT 181.315 33.580 182.440 33.750 ;
        RECT 182.610 34.380 182.805 34.710 ;
        RECT 183.030 34.380 183.285 34.710 ;
        RECT 182.610 33.410 182.780 34.380 ;
        RECT 183.455 34.210 183.625 34.880 ;
        RECT 184.075 34.810 184.320 35.415 ;
        RECT 184.540 35.085 185.050 35.620 ;
        RECT 180.750 33.240 182.780 33.410 ;
        RECT 182.950 33.070 183.120 34.210 ;
        RECT 183.290 33.240 183.625 34.210 ;
        RECT 183.800 34.640 185.030 34.810 ;
        RECT 183.800 33.830 184.140 34.640 ;
        RECT 184.310 34.075 185.060 34.265 ;
        RECT 183.800 33.420 184.315 33.830 ;
        RECT 184.550 33.070 184.720 33.830 ;
        RECT 184.890 33.410 185.060 34.075 ;
        RECT 185.230 34.090 185.420 35.450 ;
        RECT 185.590 35.280 185.865 35.450 ;
        RECT 185.590 35.110 185.870 35.280 ;
        RECT 185.590 34.290 185.865 35.110 ;
        RECT 186.055 35.085 186.585 35.450 ;
        RECT 187.010 35.220 187.340 35.620 ;
        RECT 186.410 35.050 186.585 35.085 ;
        RECT 186.070 34.090 186.240 34.890 ;
        RECT 185.230 33.920 186.240 34.090 ;
        RECT 186.410 34.880 187.340 35.050 ;
        RECT 187.510 34.880 187.765 35.450 ;
        RECT 187.940 34.895 188.230 35.620 ;
        RECT 188.405 34.910 188.660 35.440 ;
        RECT 188.830 35.160 189.135 35.620 ;
        RECT 189.380 35.240 190.450 35.410 ;
        RECT 186.410 33.750 186.580 34.880 ;
        RECT 187.170 34.710 187.340 34.880 ;
        RECT 185.455 33.580 186.580 33.750 ;
        RECT 186.750 34.380 186.945 34.710 ;
        RECT 187.170 34.380 187.425 34.710 ;
        RECT 186.750 33.410 186.920 34.380 ;
        RECT 187.595 34.210 187.765 34.880 ;
        RECT 188.405 34.260 188.615 34.910 ;
        RECT 189.380 34.885 189.700 35.240 ;
        RECT 189.375 34.710 189.700 34.885 ;
        RECT 188.785 34.410 189.700 34.710 ;
        RECT 189.870 34.670 190.110 35.070 ;
        RECT 190.280 35.010 190.450 35.240 ;
        RECT 190.620 35.180 190.810 35.620 ;
        RECT 190.980 35.170 191.930 35.450 ;
        RECT 192.150 35.260 192.500 35.430 ;
        RECT 190.280 34.840 190.810 35.010 ;
        RECT 188.785 34.380 189.525 34.410 ;
        RECT 184.890 33.240 186.920 33.410 ;
        RECT 187.090 33.070 187.260 34.210 ;
        RECT 187.430 33.240 187.765 34.210 ;
        RECT 187.940 33.070 188.230 34.235 ;
        RECT 188.405 33.380 188.660 34.260 ;
        RECT 188.830 33.070 189.135 34.210 ;
        RECT 189.355 33.790 189.525 34.380 ;
        RECT 189.870 34.300 190.410 34.670 ;
        RECT 190.590 34.560 190.810 34.840 ;
        RECT 190.980 34.390 191.150 35.170 ;
        RECT 190.745 34.220 191.150 34.390 ;
        RECT 191.320 34.380 191.670 35.000 ;
        RECT 190.745 34.130 190.915 34.220 ;
        RECT 191.840 34.210 192.050 35.000 ;
        RECT 189.695 33.960 190.915 34.130 ;
        RECT 191.375 34.050 192.050 34.210 ;
        RECT 189.355 33.620 190.155 33.790 ;
        RECT 189.475 33.070 189.805 33.450 ;
        RECT 189.985 33.330 190.155 33.620 ;
        RECT 190.745 33.580 190.915 33.960 ;
        RECT 191.085 34.040 192.050 34.050 ;
        RECT 192.240 34.870 192.500 35.260 ;
        RECT 192.710 35.160 193.040 35.620 ;
        RECT 193.915 35.230 194.770 35.400 ;
        RECT 194.975 35.230 195.470 35.400 ;
        RECT 195.640 35.260 195.970 35.620 ;
        RECT 192.240 34.180 192.410 34.870 ;
        RECT 192.580 34.520 192.750 34.700 ;
        RECT 192.920 34.690 193.710 34.940 ;
        RECT 193.915 34.520 194.085 35.230 ;
        RECT 194.255 34.720 194.610 34.940 ;
        RECT 192.580 34.350 194.270 34.520 ;
        RECT 191.085 33.750 191.545 34.040 ;
        RECT 192.240 34.010 193.740 34.180 ;
        RECT 192.240 33.870 192.410 34.010 ;
        RECT 191.850 33.700 192.410 33.870 ;
        RECT 190.325 33.070 190.575 33.530 ;
        RECT 190.745 33.240 191.615 33.580 ;
        RECT 191.850 33.240 192.020 33.700 ;
        RECT 192.855 33.670 193.930 33.840 ;
        RECT 192.190 33.070 192.560 33.530 ;
        RECT 192.855 33.330 193.025 33.670 ;
        RECT 193.195 33.070 193.525 33.500 ;
        RECT 193.760 33.330 193.930 33.670 ;
        RECT 194.100 33.570 194.270 34.350 ;
        RECT 194.440 34.130 194.610 34.720 ;
        RECT 194.780 34.320 195.130 34.940 ;
        RECT 194.440 33.740 194.905 34.130 ;
        RECT 195.300 33.870 195.470 35.230 ;
        RECT 195.640 34.040 196.100 35.090 ;
        RECT 195.075 33.700 195.470 33.870 ;
        RECT 195.075 33.570 195.245 33.700 ;
        RECT 194.100 33.240 194.780 33.570 ;
        RECT 194.995 33.240 195.245 33.570 ;
        RECT 195.415 33.070 195.665 33.530 ;
        RECT 195.835 33.255 196.160 34.040 ;
        RECT 196.330 33.240 196.500 35.360 ;
        RECT 196.670 35.240 197.000 35.620 ;
        RECT 197.170 35.070 197.425 35.360 ;
        RECT 196.675 34.900 197.425 35.070 ;
        RECT 196.675 33.910 196.905 34.900 ;
        RECT 197.600 34.850 200.190 35.620 ;
        RECT 200.365 35.070 200.620 35.360 ;
        RECT 200.790 35.240 201.120 35.620 ;
        RECT 200.365 34.900 201.115 35.070 ;
        RECT 197.075 34.080 197.425 34.730 ;
        RECT 197.600 34.330 198.810 34.850 ;
        RECT 198.980 34.160 200.190 34.680 ;
        RECT 196.675 33.740 197.425 33.910 ;
        RECT 196.670 33.070 197.000 33.570 ;
        RECT 197.170 33.240 197.425 33.740 ;
        RECT 197.600 33.070 200.190 34.160 ;
        RECT 200.365 34.080 200.715 34.730 ;
        RECT 200.885 33.910 201.115 34.900 ;
        RECT 200.365 33.740 201.115 33.910 ;
        RECT 200.365 33.240 200.620 33.740 ;
        RECT 200.790 33.070 201.120 33.570 ;
        RECT 201.290 33.240 201.460 35.360 ;
        RECT 201.820 35.260 202.150 35.620 ;
        RECT 202.320 35.230 202.815 35.400 ;
        RECT 203.020 35.230 203.875 35.400 ;
        RECT 201.690 34.040 202.150 35.090 ;
        RECT 201.630 33.255 201.955 34.040 ;
        RECT 202.320 33.870 202.490 35.230 ;
        RECT 202.660 34.320 203.010 34.940 ;
        RECT 203.180 34.720 203.535 34.940 ;
        RECT 203.180 34.130 203.350 34.720 ;
        RECT 203.705 34.520 203.875 35.230 ;
        RECT 204.750 35.160 205.080 35.620 ;
        RECT 205.290 35.260 205.640 35.430 ;
        RECT 204.080 34.690 204.870 34.940 ;
        RECT 205.290 34.870 205.550 35.260 ;
        RECT 205.860 35.170 206.810 35.450 ;
        RECT 206.980 35.180 207.170 35.620 ;
        RECT 207.340 35.240 208.410 35.410 ;
        RECT 205.040 34.520 205.210 34.700 ;
        RECT 202.320 33.700 202.715 33.870 ;
        RECT 202.885 33.740 203.350 34.130 ;
        RECT 203.520 34.350 205.210 34.520 ;
        RECT 202.545 33.570 202.715 33.700 ;
        RECT 203.520 33.570 203.690 34.350 ;
        RECT 205.380 34.180 205.550 34.870 ;
        RECT 204.050 34.010 205.550 34.180 ;
        RECT 205.740 34.210 205.950 35.000 ;
        RECT 206.120 34.380 206.470 35.000 ;
        RECT 206.640 34.390 206.810 35.170 ;
        RECT 207.340 35.010 207.510 35.240 ;
        RECT 206.980 34.840 207.510 35.010 ;
        RECT 206.980 34.560 207.200 34.840 ;
        RECT 207.680 34.670 207.920 35.070 ;
        RECT 206.640 34.220 207.045 34.390 ;
        RECT 207.380 34.300 207.920 34.670 ;
        RECT 208.090 34.885 208.410 35.240 ;
        RECT 208.655 35.160 208.960 35.620 ;
        RECT 209.130 34.910 209.385 35.440 ;
        RECT 208.090 34.710 208.415 34.885 ;
        RECT 208.090 34.410 209.005 34.710 ;
        RECT 208.265 34.380 209.005 34.410 ;
        RECT 205.740 34.050 206.415 34.210 ;
        RECT 206.875 34.130 207.045 34.220 ;
        RECT 205.740 34.040 206.705 34.050 ;
        RECT 205.380 33.870 205.550 34.010 ;
        RECT 202.125 33.070 202.375 33.530 ;
        RECT 202.545 33.240 202.795 33.570 ;
        RECT 203.010 33.240 203.690 33.570 ;
        RECT 203.860 33.670 204.935 33.840 ;
        RECT 205.380 33.700 205.940 33.870 ;
        RECT 206.245 33.750 206.705 34.040 ;
        RECT 206.875 33.960 208.095 34.130 ;
        RECT 203.860 33.330 204.030 33.670 ;
        RECT 204.265 33.070 204.595 33.500 ;
        RECT 204.765 33.330 204.935 33.670 ;
        RECT 205.230 33.070 205.600 33.530 ;
        RECT 205.770 33.240 205.940 33.700 ;
        RECT 206.875 33.580 207.045 33.960 ;
        RECT 208.265 33.790 208.435 34.380 ;
        RECT 209.175 34.260 209.385 34.910 ;
        RECT 210.135 34.990 210.420 35.450 ;
        RECT 210.590 35.160 210.860 35.620 ;
        RECT 210.135 34.820 211.090 34.990 ;
        RECT 206.175 33.240 207.045 33.580 ;
        RECT 207.635 33.620 208.435 33.790 ;
        RECT 207.215 33.070 207.465 33.530 ;
        RECT 207.635 33.330 207.805 33.620 ;
        RECT 207.985 33.070 208.315 33.450 ;
        RECT 208.655 33.070 208.960 34.210 ;
        RECT 209.130 33.380 209.385 34.260 ;
        RECT 210.020 34.090 210.710 34.650 ;
        RECT 210.880 33.920 211.090 34.820 ;
        RECT 210.135 33.700 211.090 33.920 ;
        RECT 211.260 34.650 211.660 35.450 ;
        RECT 211.850 34.990 212.130 35.450 ;
        RECT 212.650 35.160 212.975 35.620 ;
        RECT 211.850 34.820 212.975 34.990 ;
        RECT 213.145 34.880 213.530 35.450 ;
        RECT 213.700 34.895 213.990 35.620 ;
        RECT 212.525 34.710 212.975 34.820 ;
        RECT 211.260 34.090 212.355 34.650 ;
        RECT 212.525 34.380 213.080 34.710 ;
        RECT 210.135 33.240 210.420 33.700 ;
        RECT 210.590 33.070 210.860 33.530 ;
        RECT 211.260 33.240 211.660 34.090 ;
        RECT 212.525 33.920 212.975 34.380 ;
        RECT 213.250 34.210 213.530 34.880 ;
        RECT 214.165 34.880 214.420 35.450 ;
        RECT 214.590 35.220 214.920 35.620 ;
        RECT 215.345 35.085 215.875 35.450 ;
        RECT 215.345 35.050 215.520 35.085 ;
        RECT 214.590 34.880 215.520 35.050 ;
        RECT 211.850 33.700 212.975 33.920 ;
        RECT 211.850 33.240 212.130 33.700 ;
        RECT 212.650 33.070 212.975 33.530 ;
        RECT 213.145 33.240 213.530 34.210 ;
        RECT 213.700 33.070 213.990 34.235 ;
        RECT 214.165 34.210 214.335 34.880 ;
        RECT 214.590 34.710 214.760 34.880 ;
        RECT 214.505 34.380 214.760 34.710 ;
        RECT 214.985 34.380 215.180 34.710 ;
        RECT 214.165 33.240 214.500 34.210 ;
        RECT 214.670 33.070 214.840 34.210 ;
        RECT 215.010 33.410 215.180 34.380 ;
        RECT 215.350 33.750 215.520 34.880 ;
        RECT 215.690 34.090 215.860 34.890 ;
        RECT 216.065 34.600 216.340 35.450 ;
        RECT 216.060 34.430 216.340 34.600 ;
        RECT 216.065 34.290 216.340 34.430 ;
        RECT 216.510 34.090 216.700 35.450 ;
        RECT 216.880 35.085 217.390 35.620 ;
        RECT 217.610 34.810 217.855 35.415 ;
        RECT 218.305 34.910 218.560 35.440 ;
        RECT 218.730 35.160 219.035 35.620 ;
        RECT 219.280 35.240 220.350 35.410 ;
        RECT 216.900 34.640 218.130 34.810 ;
        RECT 215.690 33.920 216.700 34.090 ;
        RECT 216.870 34.075 217.620 34.265 ;
        RECT 215.350 33.580 216.475 33.750 ;
        RECT 216.870 33.410 217.040 34.075 ;
        RECT 217.790 33.830 218.130 34.640 ;
        RECT 215.010 33.240 217.040 33.410 ;
        RECT 217.210 33.070 217.380 33.830 ;
        RECT 217.615 33.420 218.130 33.830 ;
        RECT 218.305 34.260 218.515 34.910 ;
        RECT 219.280 34.885 219.600 35.240 ;
        RECT 219.275 34.710 219.600 34.885 ;
        RECT 218.685 34.410 219.600 34.710 ;
        RECT 219.770 34.670 220.010 35.070 ;
        RECT 220.180 35.010 220.350 35.240 ;
        RECT 220.520 35.180 220.710 35.620 ;
        RECT 220.880 35.170 221.830 35.450 ;
        RECT 222.050 35.260 222.400 35.430 ;
        RECT 220.180 34.840 220.710 35.010 ;
        RECT 218.685 34.380 219.425 34.410 ;
        RECT 218.305 33.380 218.560 34.260 ;
        RECT 218.730 33.070 219.035 34.210 ;
        RECT 219.255 33.790 219.425 34.380 ;
        RECT 219.770 34.300 220.310 34.670 ;
        RECT 220.490 34.560 220.710 34.840 ;
        RECT 220.880 34.390 221.050 35.170 ;
        RECT 220.645 34.220 221.050 34.390 ;
        RECT 221.220 34.380 221.570 35.000 ;
        RECT 220.645 34.130 220.815 34.220 ;
        RECT 221.740 34.210 221.950 35.000 ;
        RECT 219.595 33.960 220.815 34.130 ;
        RECT 221.275 34.050 221.950 34.210 ;
        RECT 219.255 33.620 220.055 33.790 ;
        RECT 219.375 33.070 219.705 33.450 ;
        RECT 219.885 33.330 220.055 33.620 ;
        RECT 220.645 33.580 220.815 33.960 ;
        RECT 220.985 34.040 221.950 34.050 ;
        RECT 222.140 34.870 222.400 35.260 ;
        RECT 222.610 35.160 222.940 35.620 ;
        RECT 223.815 35.230 224.670 35.400 ;
        RECT 224.875 35.230 225.370 35.400 ;
        RECT 225.540 35.260 225.870 35.620 ;
        RECT 222.140 34.180 222.310 34.870 ;
        RECT 222.480 34.520 222.650 34.700 ;
        RECT 222.820 34.690 223.610 34.940 ;
        RECT 223.815 34.520 223.985 35.230 ;
        RECT 224.155 34.720 224.510 34.940 ;
        RECT 222.480 34.350 224.170 34.520 ;
        RECT 220.985 33.750 221.445 34.040 ;
        RECT 222.140 34.010 223.640 34.180 ;
        RECT 222.140 33.870 222.310 34.010 ;
        RECT 221.750 33.700 222.310 33.870 ;
        RECT 220.225 33.070 220.475 33.530 ;
        RECT 220.645 33.240 221.515 33.580 ;
        RECT 221.750 33.240 221.920 33.700 ;
        RECT 222.755 33.670 223.830 33.840 ;
        RECT 222.090 33.070 222.460 33.530 ;
        RECT 222.755 33.330 222.925 33.670 ;
        RECT 223.095 33.070 223.425 33.500 ;
        RECT 223.660 33.330 223.830 33.670 ;
        RECT 224.000 33.570 224.170 34.350 ;
        RECT 224.340 34.130 224.510 34.720 ;
        RECT 224.680 34.320 225.030 34.940 ;
        RECT 224.340 33.740 224.805 34.130 ;
        RECT 225.200 33.870 225.370 35.230 ;
        RECT 225.540 34.040 226.000 35.090 ;
        RECT 224.975 33.700 225.370 33.870 ;
        RECT 224.975 33.570 225.145 33.700 ;
        RECT 224.000 33.240 224.680 33.570 ;
        RECT 224.895 33.240 225.145 33.570 ;
        RECT 225.315 33.070 225.565 33.530 ;
        RECT 225.735 33.255 226.060 34.040 ;
        RECT 226.230 33.240 226.400 35.360 ;
        RECT 226.570 35.240 226.900 35.620 ;
        RECT 227.070 35.070 227.325 35.360 ;
        RECT 226.575 34.900 227.325 35.070 ;
        RECT 226.575 33.910 226.805 34.900 ;
        RECT 227.500 34.850 229.170 35.620 ;
        RECT 229.345 35.070 229.600 35.360 ;
        RECT 229.770 35.240 230.100 35.620 ;
        RECT 229.345 34.900 230.095 35.070 ;
        RECT 226.975 34.080 227.325 34.730 ;
        RECT 227.500 34.330 228.250 34.850 ;
        RECT 228.420 34.160 229.170 34.680 ;
        RECT 226.575 33.740 227.325 33.910 ;
        RECT 226.570 33.070 226.900 33.570 ;
        RECT 227.070 33.240 227.325 33.740 ;
        RECT 227.500 33.070 229.170 34.160 ;
        RECT 229.345 34.080 229.695 34.730 ;
        RECT 229.865 33.910 230.095 34.900 ;
        RECT 229.345 33.740 230.095 33.910 ;
        RECT 229.345 33.240 229.600 33.740 ;
        RECT 229.770 33.070 230.100 33.570 ;
        RECT 230.270 33.240 230.440 35.360 ;
        RECT 230.800 35.260 231.130 35.620 ;
        RECT 231.300 35.230 231.795 35.400 ;
        RECT 232.000 35.230 232.855 35.400 ;
        RECT 230.670 34.040 231.130 35.090 ;
        RECT 230.610 33.255 230.935 34.040 ;
        RECT 231.300 33.870 231.470 35.230 ;
        RECT 231.640 34.320 231.990 34.940 ;
        RECT 232.160 34.720 232.515 34.940 ;
        RECT 232.160 34.130 232.330 34.720 ;
        RECT 232.685 34.520 232.855 35.230 ;
        RECT 233.730 35.160 234.060 35.620 ;
        RECT 234.270 35.260 234.620 35.430 ;
        RECT 233.060 34.690 233.850 34.940 ;
        RECT 234.270 34.870 234.530 35.260 ;
        RECT 234.840 35.170 235.790 35.450 ;
        RECT 235.960 35.180 236.150 35.620 ;
        RECT 236.320 35.240 237.390 35.410 ;
        RECT 234.020 34.520 234.190 34.700 ;
        RECT 231.300 33.700 231.695 33.870 ;
        RECT 231.865 33.740 232.330 34.130 ;
        RECT 232.500 34.350 234.190 34.520 ;
        RECT 231.525 33.570 231.695 33.700 ;
        RECT 232.500 33.570 232.670 34.350 ;
        RECT 234.360 34.180 234.530 34.870 ;
        RECT 233.030 34.010 234.530 34.180 ;
        RECT 234.720 34.210 234.930 35.000 ;
        RECT 235.100 34.380 235.450 35.000 ;
        RECT 235.620 34.390 235.790 35.170 ;
        RECT 236.320 35.010 236.490 35.240 ;
        RECT 235.960 34.840 236.490 35.010 ;
        RECT 235.960 34.560 236.180 34.840 ;
        RECT 236.660 34.670 236.900 35.070 ;
        RECT 235.620 34.220 236.025 34.390 ;
        RECT 236.360 34.300 236.900 34.670 ;
        RECT 237.070 34.885 237.390 35.240 ;
        RECT 237.635 35.160 237.940 35.620 ;
        RECT 238.110 34.910 238.365 35.440 ;
        RECT 237.070 34.710 237.395 34.885 ;
        RECT 237.070 34.410 237.985 34.710 ;
        RECT 237.245 34.380 237.985 34.410 ;
        RECT 234.720 34.050 235.395 34.210 ;
        RECT 235.855 34.130 236.025 34.220 ;
        RECT 234.720 34.040 235.685 34.050 ;
        RECT 234.360 33.870 234.530 34.010 ;
        RECT 231.105 33.070 231.355 33.530 ;
        RECT 231.525 33.240 231.775 33.570 ;
        RECT 231.990 33.240 232.670 33.570 ;
        RECT 232.840 33.670 233.915 33.840 ;
        RECT 234.360 33.700 234.920 33.870 ;
        RECT 235.225 33.750 235.685 34.040 ;
        RECT 235.855 33.960 237.075 34.130 ;
        RECT 232.840 33.330 233.010 33.670 ;
        RECT 233.245 33.070 233.575 33.500 ;
        RECT 233.745 33.330 233.915 33.670 ;
        RECT 234.210 33.070 234.580 33.530 ;
        RECT 234.750 33.240 234.920 33.700 ;
        RECT 235.855 33.580 236.025 33.960 ;
        RECT 237.245 33.790 237.415 34.380 ;
        RECT 238.155 34.260 238.365 34.910 ;
        RECT 239.460 34.895 239.750 35.620 ;
        RECT 240.385 35.070 240.640 35.360 ;
        RECT 240.810 35.240 241.140 35.620 ;
        RECT 240.385 34.900 241.135 35.070 ;
        RECT 235.155 33.240 236.025 33.580 ;
        RECT 236.615 33.620 237.415 33.790 ;
        RECT 236.195 33.070 236.445 33.530 ;
        RECT 236.615 33.330 236.785 33.620 ;
        RECT 236.965 33.070 237.295 33.450 ;
        RECT 237.635 33.070 237.940 34.210 ;
        RECT 238.110 33.380 238.365 34.260 ;
        RECT 239.460 33.070 239.750 34.235 ;
        RECT 240.385 34.080 240.735 34.730 ;
        RECT 240.905 33.910 241.135 34.900 ;
        RECT 240.385 33.740 241.135 33.910 ;
        RECT 240.385 33.240 240.640 33.740 ;
        RECT 240.810 33.070 241.140 33.570 ;
        RECT 241.310 33.240 241.480 35.360 ;
        RECT 241.840 35.260 242.170 35.620 ;
        RECT 242.340 35.230 242.835 35.400 ;
        RECT 243.040 35.230 243.895 35.400 ;
        RECT 241.710 34.040 242.170 35.090 ;
        RECT 241.650 33.255 241.975 34.040 ;
        RECT 242.340 33.870 242.510 35.230 ;
        RECT 242.680 34.320 243.030 34.940 ;
        RECT 243.200 34.720 243.555 34.940 ;
        RECT 243.200 34.130 243.370 34.720 ;
        RECT 243.725 34.520 243.895 35.230 ;
        RECT 244.770 35.160 245.100 35.620 ;
        RECT 245.310 35.260 245.660 35.430 ;
        RECT 244.100 34.690 244.890 34.940 ;
        RECT 245.310 34.870 245.570 35.260 ;
        RECT 245.880 35.170 246.830 35.450 ;
        RECT 247.000 35.180 247.190 35.620 ;
        RECT 247.360 35.240 248.430 35.410 ;
        RECT 245.060 34.520 245.230 34.700 ;
        RECT 242.340 33.700 242.735 33.870 ;
        RECT 242.905 33.740 243.370 34.130 ;
        RECT 243.540 34.350 245.230 34.520 ;
        RECT 242.565 33.570 242.735 33.700 ;
        RECT 243.540 33.570 243.710 34.350 ;
        RECT 245.400 34.180 245.570 34.870 ;
        RECT 244.070 34.010 245.570 34.180 ;
        RECT 245.760 34.210 245.970 35.000 ;
        RECT 246.140 34.380 246.490 35.000 ;
        RECT 246.660 34.390 246.830 35.170 ;
        RECT 247.360 35.010 247.530 35.240 ;
        RECT 247.000 34.840 247.530 35.010 ;
        RECT 247.000 34.560 247.220 34.840 ;
        RECT 247.700 34.670 247.940 35.070 ;
        RECT 246.660 34.220 247.065 34.390 ;
        RECT 247.400 34.300 247.940 34.670 ;
        RECT 248.110 34.885 248.430 35.240 ;
        RECT 248.675 35.160 248.980 35.620 ;
        RECT 249.150 34.910 249.405 35.440 ;
        RECT 249.580 35.075 254.925 35.620 ;
        RECT 248.110 34.710 248.435 34.885 ;
        RECT 248.110 34.410 249.025 34.710 ;
        RECT 248.285 34.380 249.025 34.410 ;
        RECT 245.760 34.050 246.435 34.210 ;
        RECT 246.895 34.130 247.065 34.220 ;
        RECT 245.760 34.040 246.725 34.050 ;
        RECT 245.400 33.870 245.570 34.010 ;
        RECT 242.145 33.070 242.395 33.530 ;
        RECT 242.565 33.240 242.815 33.570 ;
        RECT 243.030 33.240 243.710 33.570 ;
        RECT 243.880 33.670 244.955 33.840 ;
        RECT 245.400 33.700 245.960 33.870 ;
        RECT 246.265 33.750 246.725 34.040 ;
        RECT 246.895 33.960 248.115 34.130 ;
        RECT 243.880 33.330 244.050 33.670 ;
        RECT 244.285 33.070 244.615 33.500 ;
        RECT 244.785 33.330 244.955 33.670 ;
        RECT 245.250 33.070 245.620 33.530 ;
        RECT 245.790 33.240 245.960 33.700 ;
        RECT 246.895 33.580 247.065 33.960 ;
        RECT 248.285 33.790 248.455 34.380 ;
        RECT 249.195 34.260 249.405 34.910 ;
        RECT 246.195 33.240 247.065 33.580 ;
        RECT 247.655 33.620 248.455 33.790 ;
        RECT 247.235 33.070 247.485 33.530 ;
        RECT 247.655 33.330 247.825 33.620 ;
        RECT 248.005 33.070 248.335 33.450 ;
        RECT 248.675 33.070 248.980 34.210 ;
        RECT 249.150 33.380 249.405 34.260 ;
        RECT 251.165 34.245 251.505 35.075 ;
        RECT 255.565 35.070 255.820 35.360 ;
        RECT 255.990 35.240 256.320 35.620 ;
        RECT 255.565 34.900 256.315 35.070 ;
        RECT 252.985 33.505 253.335 34.755 ;
        RECT 255.565 34.080 255.915 34.730 ;
        RECT 256.085 33.910 256.315 34.900 ;
        RECT 255.565 33.740 256.315 33.910 ;
        RECT 249.580 33.070 254.925 33.505 ;
        RECT 255.565 33.240 255.820 33.740 ;
        RECT 255.990 33.070 256.320 33.570 ;
        RECT 256.490 33.240 256.660 35.360 ;
        RECT 257.020 35.260 257.350 35.620 ;
        RECT 257.520 35.230 258.015 35.400 ;
        RECT 258.220 35.230 259.075 35.400 ;
        RECT 256.890 34.040 257.350 35.090 ;
        RECT 256.830 33.255 257.155 34.040 ;
        RECT 257.520 33.870 257.690 35.230 ;
        RECT 257.860 34.320 258.210 34.940 ;
        RECT 258.380 34.720 258.735 34.940 ;
        RECT 258.380 34.130 258.550 34.720 ;
        RECT 258.905 34.520 259.075 35.230 ;
        RECT 259.950 35.160 260.280 35.620 ;
        RECT 260.490 35.260 260.840 35.430 ;
        RECT 259.280 34.690 260.070 34.940 ;
        RECT 260.490 34.870 260.750 35.260 ;
        RECT 261.060 35.170 262.010 35.450 ;
        RECT 262.180 35.180 262.370 35.620 ;
        RECT 262.540 35.240 263.610 35.410 ;
        RECT 260.240 34.520 260.410 34.700 ;
        RECT 257.520 33.700 257.915 33.870 ;
        RECT 258.085 33.740 258.550 34.130 ;
        RECT 258.720 34.350 260.410 34.520 ;
        RECT 257.745 33.570 257.915 33.700 ;
        RECT 258.720 33.570 258.890 34.350 ;
        RECT 260.580 34.180 260.750 34.870 ;
        RECT 259.250 34.010 260.750 34.180 ;
        RECT 260.940 34.210 261.150 35.000 ;
        RECT 261.320 34.380 261.670 35.000 ;
        RECT 261.840 34.390 262.010 35.170 ;
        RECT 262.540 35.010 262.710 35.240 ;
        RECT 262.180 34.840 262.710 35.010 ;
        RECT 262.180 34.560 262.400 34.840 ;
        RECT 262.880 34.670 263.120 35.070 ;
        RECT 261.840 34.220 262.245 34.390 ;
        RECT 262.580 34.300 263.120 34.670 ;
        RECT 263.290 34.885 263.610 35.240 ;
        RECT 263.855 35.160 264.160 35.620 ;
        RECT 264.330 34.910 264.585 35.440 ;
        RECT 263.290 34.710 263.615 34.885 ;
        RECT 263.290 34.410 264.205 34.710 ;
        RECT 263.465 34.380 264.205 34.410 ;
        RECT 260.940 34.050 261.615 34.210 ;
        RECT 262.075 34.130 262.245 34.220 ;
        RECT 260.940 34.040 261.905 34.050 ;
        RECT 260.580 33.870 260.750 34.010 ;
        RECT 257.325 33.070 257.575 33.530 ;
        RECT 257.745 33.240 257.995 33.570 ;
        RECT 258.210 33.240 258.890 33.570 ;
        RECT 259.060 33.670 260.135 33.840 ;
        RECT 260.580 33.700 261.140 33.870 ;
        RECT 261.445 33.750 261.905 34.040 ;
        RECT 262.075 33.960 263.295 34.130 ;
        RECT 259.060 33.330 259.230 33.670 ;
        RECT 259.465 33.070 259.795 33.500 ;
        RECT 259.965 33.330 260.135 33.670 ;
        RECT 260.430 33.070 260.800 33.530 ;
        RECT 260.970 33.240 261.140 33.700 ;
        RECT 262.075 33.580 262.245 33.960 ;
        RECT 263.465 33.790 263.635 34.380 ;
        RECT 264.375 34.260 264.585 34.910 ;
        RECT 265.220 34.895 265.510 35.620 ;
        RECT 265.680 35.160 266.240 35.450 ;
        RECT 266.410 35.160 266.660 35.620 ;
        RECT 261.375 33.240 262.245 33.580 ;
        RECT 262.835 33.620 263.635 33.790 ;
        RECT 262.415 33.070 262.665 33.530 ;
        RECT 262.835 33.330 263.005 33.620 ;
        RECT 263.185 33.070 263.515 33.450 ;
        RECT 263.855 33.070 264.160 34.210 ;
        RECT 264.330 33.380 264.585 34.260 ;
        RECT 265.220 33.070 265.510 34.235 ;
        RECT 265.680 33.790 265.930 35.160 ;
        RECT 267.280 34.990 267.610 35.350 ;
        RECT 267.980 35.075 273.325 35.620 ;
        RECT 273.500 35.075 278.845 35.620 ;
        RECT 279.020 35.075 284.365 35.620 ;
        RECT 284.540 35.075 289.885 35.620 ;
        RECT 266.220 34.800 267.610 34.990 ;
        RECT 266.220 34.710 266.390 34.800 ;
        RECT 266.100 34.380 266.390 34.710 ;
        RECT 266.560 34.380 266.900 34.630 ;
        RECT 267.120 34.380 267.795 34.630 ;
        RECT 266.220 34.130 266.390 34.380 ;
        RECT 266.220 33.960 267.160 34.130 ;
        RECT 267.530 34.020 267.795 34.380 ;
        RECT 269.565 34.245 269.905 35.075 ;
        RECT 265.680 33.240 266.140 33.790 ;
        RECT 266.330 33.070 266.660 33.790 ;
        RECT 266.860 33.410 267.160 33.960 ;
        RECT 267.330 33.070 267.610 33.740 ;
        RECT 271.385 33.505 271.735 34.755 ;
        RECT 275.085 34.245 275.425 35.075 ;
        RECT 276.905 33.505 277.255 34.755 ;
        RECT 280.605 34.245 280.945 35.075 ;
        RECT 282.425 33.505 282.775 34.755 ;
        RECT 286.125 34.245 286.465 35.075 ;
        RECT 290.980 34.895 291.270 35.620 ;
        RECT 291.440 35.075 296.785 35.620 ;
        RECT 287.945 33.505 288.295 34.755 ;
        RECT 293.025 34.245 293.365 35.075 ;
        RECT 296.960 34.850 299.550 35.620 ;
        RECT 299.725 34.910 299.980 35.440 ;
        RECT 300.150 35.160 300.455 35.620 ;
        RECT 300.700 35.240 301.770 35.410 ;
        RECT 267.980 33.070 273.325 33.505 ;
        RECT 273.500 33.070 278.845 33.505 ;
        RECT 279.020 33.070 284.365 33.505 ;
        RECT 284.540 33.070 289.885 33.505 ;
        RECT 290.980 33.070 291.270 34.235 ;
        RECT 294.845 33.505 295.195 34.755 ;
        RECT 296.960 34.330 298.170 34.850 ;
        RECT 298.340 34.160 299.550 34.680 ;
        RECT 291.440 33.070 296.785 33.505 ;
        RECT 296.960 33.070 299.550 34.160 ;
        RECT 299.725 34.260 299.935 34.910 ;
        RECT 300.700 34.885 301.020 35.240 ;
        RECT 300.695 34.710 301.020 34.885 ;
        RECT 300.105 34.410 301.020 34.710 ;
        RECT 301.190 34.670 301.430 35.070 ;
        RECT 301.600 35.010 301.770 35.240 ;
        RECT 301.940 35.180 302.130 35.620 ;
        RECT 302.300 35.170 303.250 35.450 ;
        RECT 303.470 35.260 303.820 35.430 ;
        RECT 301.600 34.840 302.130 35.010 ;
        RECT 300.105 34.380 300.845 34.410 ;
        RECT 299.725 33.380 299.980 34.260 ;
        RECT 300.150 33.070 300.455 34.210 ;
        RECT 300.675 33.790 300.845 34.380 ;
        RECT 301.190 34.300 301.730 34.670 ;
        RECT 301.910 34.560 302.130 34.840 ;
        RECT 302.300 34.390 302.470 35.170 ;
        RECT 302.065 34.220 302.470 34.390 ;
        RECT 302.640 34.380 302.990 35.000 ;
        RECT 302.065 34.130 302.235 34.220 ;
        RECT 303.160 34.210 303.370 35.000 ;
        RECT 301.015 33.960 302.235 34.130 ;
        RECT 302.695 34.050 303.370 34.210 ;
        RECT 300.675 33.620 301.475 33.790 ;
        RECT 300.795 33.070 301.125 33.450 ;
        RECT 301.305 33.330 301.475 33.620 ;
        RECT 302.065 33.580 302.235 33.960 ;
        RECT 302.405 34.040 303.370 34.050 ;
        RECT 303.560 34.870 303.820 35.260 ;
        RECT 304.030 35.160 304.360 35.620 ;
        RECT 305.235 35.230 306.090 35.400 ;
        RECT 306.295 35.230 306.790 35.400 ;
        RECT 306.960 35.260 307.290 35.620 ;
        RECT 303.560 34.180 303.730 34.870 ;
        RECT 303.900 34.520 304.070 34.700 ;
        RECT 304.240 34.690 305.030 34.940 ;
        RECT 305.235 34.520 305.405 35.230 ;
        RECT 305.575 34.720 305.930 34.940 ;
        RECT 303.900 34.350 305.590 34.520 ;
        RECT 302.405 33.750 302.865 34.040 ;
        RECT 303.560 34.010 305.060 34.180 ;
        RECT 303.560 33.870 303.730 34.010 ;
        RECT 303.170 33.700 303.730 33.870 ;
        RECT 301.645 33.070 301.895 33.530 ;
        RECT 302.065 33.240 302.935 33.580 ;
        RECT 303.170 33.240 303.340 33.700 ;
        RECT 304.175 33.670 305.250 33.840 ;
        RECT 303.510 33.070 303.880 33.530 ;
        RECT 304.175 33.330 304.345 33.670 ;
        RECT 304.515 33.070 304.845 33.500 ;
        RECT 305.080 33.330 305.250 33.670 ;
        RECT 305.420 33.570 305.590 34.350 ;
        RECT 305.760 34.130 305.930 34.720 ;
        RECT 306.100 34.320 306.450 34.940 ;
        RECT 305.760 33.740 306.225 34.130 ;
        RECT 306.620 33.870 306.790 35.230 ;
        RECT 306.960 34.040 307.420 35.090 ;
        RECT 306.395 33.700 306.790 33.870 ;
        RECT 306.395 33.570 306.565 33.700 ;
        RECT 305.420 33.240 306.100 33.570 ;
        RECT 306.315 33.240 306.565 33.570 ;
        RECT 306.735 33.070 306.985 33.530 ;
        RECT 307.155 33.255 307.480 34.040 ;
        RECT 307.650 33.240 307.820 35.360 ;
        RECT 307.990 35.240 308.320 35.620 ;
        RECT 308.490 35.070 308.745 35.360 ;
        RECT 307.995 34.900 308.745 35.070 ;
        RECT 307.995 33.910 308.225 34.900 ;
        RECT 309.840 34.870 311.050 35.620 ;
        RECT 308.395 34.080 308.745 34.730 ;
        RECT 309.840 34.160 310.360 34.700 ;
        RECT 310.530 34.330 311.050 34.870 ;
        RECT 307.995 33.740 308.745 33.910 ;
        RECT 307.990 33.070 308.320 33.570 ;
        RECT 308.490 33.240 308.745 33.740 ;
        RECT 309.840 33.070 311.050 34.160 ;
        RECT 162.095 32.900 311.135 33.070 ;
        RECT 162.180 31.810 163.390 32.900 ;
        RECT 163.560 31.810 165.230 32.900 ;
        RECT 165.865 32.230 166.120 32.730 ;
        RECT 166.290 32.400 166.620 32.900 ;
        RECT 165.865 32.060 166.615 32.230 ;
        RECT 162.180 31.100 162.700 31.640 ;
        RECT 162.870 31.270 163.390 31.810 ;
        RECT 163.560 31.120 164.310 31.640 ;
        RECT 164.480 31.290 165.230 31.810 ;
        RECT 165.865 31.240 166.215 31.890 ;
        RECT 162.180 30.350 163.390 31.100 ;
        RECT 163.560 30.350 165.230 31.120 ;
        RECT 166.385 31.070 166.615 32.060 ;
        RECT 165.865 30.900 166.615 31.070 ;
        RECT 165.865 30.610 166.120 30.900 ;
        RECT 166.290 30.350 166.620 30.730 ;
        RECT 166.790 30.610 166.960 32.730 ;
        RECT 167.130 31.930 167.455 32.715 ;
        RECT 167.625 32.440 167.875 32.900 ;
        RECT 168.045 32.400 168.295 32.730 ;
        RECT 168.510 32.400 169.190 32.730 ;
        RECT 168.045 32.270 168.215 32.400 ;
        RECT 167.820 32.100 168.215 32.270 ;
        RECT 167.190 30.880 167.650 31.930 ;
        RECT 167.820 30.740 167.990 32.100 ;
        RECT 168.385 31.840 168.850 32.230 ;
        RECT 168.160 31.030 168.510 31.650 ;
        RECT 168.680 31.250 168.850 31.840 ;
        RECT 169.020 31.620 169.190 32.400 ;
        RECT 169.360 32.300 169.530 32.640 ;
        RECT 169.765 32.470 170.095 32.900 ;
        RECT 170.265 32.300 170.435 32.640 ;
        RECT 170.730 32.440 171.100 32.900 ;
        RECT 169.360 32.130 170.435 32.300 ;
        RECT 171.270 32.270 171.440 32.730 ;
        RECT 171.675 32.390 172.545 32.730 ;
        RECT 172.715 32.440 172.965 32.900 ;
        RECT 170.880 32.100 171.440 32.270 ;
        RECT 170.880 31.960 171.050 32.100 ;
        RECT 169.550 31.790 171.050 31.960 ;
        RECT 171.745 31.930 172.205 32.220 ;
        RECT 169.020 31.450 170.710 31.620 ;
        RECT 168.680 31.030 169.035 31.250 ;
        RECT 169.205 30.740 169.375 31.450 ;
        RECT 169.580 31.030 170.370 31.280 ;
        RECT 170.540 31.270 170.710 31.450 ;
        RECT 170.880 31.100 171.050 31.790 ;
        RECT 167.320 30.350 167.650 30.710 ;
        RECT 167.820 30.570 168.315 30.740 ;
        RECT 168.520 30.570 169.375 30.740 ;
        RECT 170.250 30.350 170.580 30.810 ;
        RECT 170.790 30.710 171.050 31.100 ;
        RECT 171.240 31.920 172.205 31.930 ;
        RECT 172.375 32.010 172.545 32.390 ;
        RECT 173.135 32.350 173.305 32.640 ;
        RECT 173.485 32.520 173.815 32.900 ;
        RECT 173.135 32.180 173.935 32.350 ;
        RECT 171.240 31.760 171.915 31.920 ;
        RECT 172.375 31.840 173.595 32.010 ;
        RECT 171.240 30.970 171.450 31.760 ;
        RECT 172.375 31.750 172.545 31.840 ;
        RECT 171.620 30.970 171.970 31.590 ;
        RECT 172.140 31.580 172.545 31.750 ;
        RECT 172.140 30.800 172.310 31.580 ;
        RECT 172.480 31.130 172.700 31.410 ;
        RECT 172.880 31.300 173.420 31.670 ;
        RECT 173.765 31.590 173.935 32.180 ;
        RECT 174.155 31.760 174.460 32.900 ;
        RECT 174.630 31.710 174.885 32.590 ;
        RECT 175.060 31.735 175.350 32.900 ;
        RECT 175.525 31.760 175.860 32.730 ;
        RECT 176.030 31.760 176.200 32.900 ;
        RECT 176.370 32.560 178.400 32.730 ;
        RECT 173.765 31.560 174.505 31.590 ;
        RECT 172.480 30.960 173.010 31.130 ;
        RECT 170.790 30.540 171.140 30.710 ;
        RECT 171.360 30.520 172.310 30.800 ;
        RECT 172.480 30.350 172.670 30.790 ;
        RECT 172.840 30.730 173.010 30.960 ;
        RECT 173.180 30.900 173.420 31.300 ;
        RECT 173.590 31.260 174.505 31.560 ;
        RECT 173.590 31.085 173.915 31.260 ;
        RECT 173.590 30.730 173.910 31.085 ;
        RECT 174.675 31.060 174.885 31.710 ;
        RECT 175.525 31.090 175.695 31.760 ;
        RECT 176.370 31.590 176.540 32.560 ;
        RECT 175.865 31.260 176.120 31.590 ;
        RECT 176.345 31.260 176.540 31.590 ;
        RECT 176.710 32.220 177.835 32.390 ;
        RECT 175.950 31.090 176.120 31.260 ;
        RECT 176.710 31.090 176.880 32.220 ;
        RECT 172.840 30.560 173.910 30.730 ;
        RECT 174.155 30.350 174.460 30.810 ;
        RECT 174.630 30.530 174.885 31.060 ;
        RECT 175.060 30.350 175.350 31.075 ;
        RECT 175.525 30.520 175.780 31.090 ;
        RECT 175.950 30.920 176.880 31.090 ;
        RECT 177.050 31.880 178.060 32.050 ;
        RECT 177.050 31.080 177.220 31.880 ;
        RECT 177.425 31.540 177.700 31.680 ;
        RECT 177.420 31.370 177.700 31.540 ;
        RECT 176.705 30.885 176.880 30.920 ;
        RECT 175.950 30.350 176.280 30.750 ;
        RECT 176.705 30.520 177.235 30.885 ;
        RECT 177.425 30.520 177.700 31.370 ;
        RECT 177.870 30.520 178.060 31.880 ;
        RECT 178.230 31.895 178.400 32.560 ;
        RECT 178.570 32.140 178.740 32.900 ;
        RECT 178.975 32.140 179.490 32.550 ;
        RECT 178.230 31.705 178.980 31.895 ;
        RECT 179.150 31.330 179.490 32.140 ;
        RECT 179.660 31.810 181.330 32.900 ;
        RECT 178.260 31.160 179.490 31.330 ;
        RECT 178.240 30.350 178.750 30.885 ;
        RECT 178.970 30.555 179.215 31.160 ;
        RECT 179.660 31.120 180.410 31.640 ;
        RECT 180.580 31.290 181.330 31.810 ;
        RECT 181.965 31.710 182.220 32.590 ;
        RECT 182.390 31.760 182.695 32.900 ;
        RECT 183.035 32.520 183.365 32.900 ;
        RECT 183.545 32.350 183.715 32.640 ;
        RECT 183.885 32.440 184.135 32.900 ;
        RECT 182.915 32.180 183.715 32.350 ;
        RECT 184.305 32.390 185.175 32.730 ;
        RECT 179.660 30.350 181.330 31.120 ;
        RECT 181.965 31.060 182.175 31.710 ;
        RECT 182.915 31.590 183.085 32.180 ;
        RECT 184.305 32.010 184.475 32.390 ;
        RECT 185.410 32.270 185.580 32.730 ;
        RECT 185.750 32.440 186.120 32.900 ;
        RECT 186.415 32.300 186.585 32.640 ;
        RECT 186.755 32.470 187.085 32.900 ;
        RECT 187.320 32.300 187.490 32.640 ;
        RECT 183.255 31.840 184.475 32.010 ;
        RECT 184.645 31.930 185.105 32.220 ;
        RECT 185.410 32.100 185.970 32.270 ;
        RECT 186.415 32.130 187.490 32.300 ;
        RECT 187.660 32.400 188.340 32.730 ;
        RECT 188.555 32.400 188.805 32.730 ;
        RECT 188.975 32.440 189.225 32.900 ;
        RECT 185.800 31.960 185.970 32.100 ;
        RECT 184.645 31.920 185.610 31.930 ;
        RECT 184.305 31.750 184.475 31.840 ;
        RECT 184.935 31.760 185.610 31.920 ;
        RECT 182.345 31.560 183.085 31.590 ;
        RECT 182.345 31.260 183.260 31.560 ;
        RECT 182.935 31.085 183.260 31.260 ;
        RECT 181.965 30.530 182.220 31.060 ;
        RECT 182.390 30.350 182.695 30.810 ;
        RECT 182.940 30.730 183.260 31.085 ;
        RECT 183.430 31.300 183.970 31.670 ;
        RECT 184.305 31.580 184.710 31.750 ;
        RECT 183.430 30.900 183.670 31.300 ;
        RECT 184.150 31.130 184.370 31.410 ;
        RECT 183.840 30.960 184.370 31.130 ;
        RECT 183.840 30.730 184.010 30.960 ;
        RECT 184.540 30.800 184.710 31.580 ;
        RECT 184.880 30.970 185.230 31.590 ;
        RECT 185.400 30.970 185.610 31.760 ;
        RECT 185.800 31.790 187.300 31.960 ;
        RECT 185.800 31.100 185.970 31.790 ;
        RECT 187.660 31.620 187.830 32.400 ;
        RECT 188.635 32.270 188.805 32.400 ;
        RECT 186.140 31.450 187.830 31.620 ;
        RECT 188.000 31.840 188.465 32.230 ;
        RECT 188.635 32.100 189.030 32.270 ;
        RECT 186.140 31.270 186.310 31.450 ;
        RECT 182.940 30.560 184.010 30.730 ;
        RECT 184.180 30.350 184.370 30.790 ;
        RECT 184.540 30.520 185.490 30.800 ;
        RECT 185.800 30.710 186.060 31.100 ;
        RECT 186.480 31.030 187.270 31.280 ;
        RECT 185.710 30.540 186.060 30.710 ;
        RECT 186.270 30.350 186.600 30.810 ;
        RECT 187.475 30.740 187.645 31.450 ;
        RECT 188.000 31.250 188.170 31.840 ;
        RECT 187.815 31.030 188.170 31.250 ;
        RECT 188.340 31.030 188.690 31.650 ;
        RECT 188.860 30.740 189.030 32.100 ;
        RECT 189.395 31.930 189.720 32.715 ;
        RECT 189.200 30.880 189.660 31.930 ;
        RECT 187.475 30.570 188.330 30.740 ;
        RECT 188.535 30.570 189.030 30.740 ;
        RECT 189.200 30.350 189.530 30.710 ;
        RECT 189.890 30.610 190.060 32.730 ;
        RECT 190.230 32.400 190.560 32.900 ;
        RECT 190.730 32.230 190.985 32.730 ;
        RECT 190.235 32.060 190.985 32.230 ;
        RECT 190.235 31.070 190.465 32.060 ;
        RECT 190.635 31.240 190.985 31.890 ;
        RECT 191.165 31.760 191.500 32.730 ;
        RECT 191.670 31.760 191.840 32.900 ;
        RECT 192.010 32.560 194.040 32.730 ;
        RECT 191.165 31.090 191.335 31.760 ;
        RECT 192.010 31.590 192.180 32.560 ;
        RECT 191.505 31.260 191.760 31.590 ;
        RECT 191.985 31.260 192.180 31.590 ;
        RECT 192.350 32.220 193.475 32.390 ;
        RECT 191.590 31.090 191.760 31.260 ;
        RECT 192.350 31.090 192.520 32.220 ;
        RECT 190.235 30.900 190.985 31.070 ;
        RECT 190.230 30.350 190.560 30.730 ;
        RECT 190.730 30.610 190.985 30.900 ;
        RECT 191.165 30.520 191.420 31.090 ;
        RECT 191.590 30.920 192.520 31.090 ;
        RECT 192.690 31.880 193.700 32.050 ;
        RECT 192.690 31.080 192.860 31.880 ;
        RECT 193.065 31.200 193.340 31.680 ;
        RECT 193.060 31.030 193.340 31.200 ;
        RECT 192.345 30.885 192.520 30.920 ;
        RECT 191.590 30.350 191.920 30.750 ;
        RECT 192.345 30.520 192.875 30.885 ;
        RECT 193.065 30.520 193.340 31.030 ;
        RECT 193.510 30.520 193.700 31.880 ;
        RECT 193.870 31.895 194.040 32.560 ;
        RECT 194.210 32.140 194.380 32.900 ;
        RECT 194.615 32.140 195.130 32.550 ;
        RECT 193.870 31.705 194.620 31.895 ;
        RECT 194.790 31.330 195.130 32.140 ;
        RECT 195.300 31.810 197.890 32.900 ;
        RECT 198.115 32.030 198.400 32.900 ;
        RECT 198.570 32.270 198.830 32.730 ;
        RECT 199.005 32.440 199.260 32.900 ;
        RECT 199.430 32.270 199.690 32.730 ;
        RECT 198.570 32.100 199.690 32.270 ;
        RECT 199.860 32.100 200.170 32.900 ;
        RECT 198.570 31.850 198.830 32.100 ;
        RECT 200.340 31.930 200.650 32.730 ;
        RECT 193.900 31.160 195.130 31.330 ;
        RECT 193.880 30.350 194.390 30.885 ;
        RECT 194.610 30.555 194.855 31.160 ;
        RECT 195.300 31.120 196.510 31.640 ;
        RECT 196.680 31.290 197.890 31.810 ;
        RECT 198.075 31.680 198.830 31.850 ;
        RECT 199.620 31.760 200.650 31.930 ;
        RECT 198.075 31.170 198.480 31.680 ;
        RECT 199.620 31.510 199.790 31.760 ;
        RECT 198.650 31.340 199.790 31.510 ;
        RECT 195.300 30.350 197.890 31.120 ;
        RECT 198.075 31.000 199.725 31.170 ;
        RECT 199.960 31.020 200.310 31.590 ;
        RECT 198.120 30.350 198.400 30.830 ;
        RECT 198.570 30.610 198.830 31.000 ;
        RECT 199.005 30.350 199.260 30.830 ;
        RECT 199.430 30.610 199.725 31.000 ;
        RECT 200.480 30.850 200.650 31.760 ;
        RECT 200.820 31.735 201.110 32.900 ;
        RECT 201.285 31.760 201.620 32.730 ;
        RECT 201.790 31.760 201.960 32.900 ;
        RECT 202.130 32.560 204.160 32.730 ;
        RECT 201.285 31.090 201.455 31.760 ;
        RECT 202.130 31.590 202.300 32.560 ;
        RECT 201.625 31.260 201.880 31.590 ;
        RECT 202.105 31.260 202.300 31.590 ;
        RECT 202.470 32.220 203.595 32.390 ;
        RECT 201.710 31.090 201.880 31.260 ;
        RECT 202.470 31.090 202.640 32.220 ;
        RECT 199.905 30.350 200.180 30.830 ;
        RECT 200.350 30.520 200.650 30.850 ;
        RECT 200.820 30.350 201.110 31.075 ;
        RECT 201.285 30.520 201.540 31.090 ;
        RECT 201.710 30.920 202.640 31.090 ;
        RECT 202.810 31.880 203.820 32.050 ;
        RECT 202.810 31.080 202.980 31.880 ;
        RECT 203.185 31.200 203.460 31.680 ;
        RECT 203.180 31.030 203.460 31.200 ;
        RECT 202.465 30.885 202.640 30.920 ;
        RECT 201.710 30.350 202.040 30.750 ;
        RECT 202.465 30.520 202.995 30.885 ;
        RECT 203.185 30.520 203.460 31.030 ;
        RECT 203.630 30.520 203.820 31.880 ;
        RECT 203.990 31.895 204.160 32.560 ;
        RECT 204.330 32.140 204.500 32.900 ;
        RECT 204.735 32.140 205.250 32.550 ;
        RECT 203.990 31.705 204.740 31.895 ;
        RECT 204.910 31.330 205.250 32.140 ;
        RECT 204.020 31.160 205.250 31.330 ;
        RECT 206.345 31.710 206.600 32.590 ;
        RECT 206.770 31.760 207.075 32.900 ;
        RECT 207.415 32.520 207.745 32.900 ;
        RECT 207.925 32.350 208.095 32.640 ;
        RECT 208.265 32.440 208.515 32.900 ;
        RECT 207.295 32.180 208.095 32.350 ;
        RECT 208.685 32.390 209.555 32.730 ;
        RECT 204.000 30.350 204.510 30.885 ;
        RECT 204.730 30.555 204.975 31.160 ;
        RECT 206.345 31.060 206.555 31.710 ;
        RECT 207.295 31.590 207.465 32.180 ;
        RECT 208.685 32.010 208.855 32.390 ;
        RECT 209.790 32.270 209.960 32.730 ;
        RECT 210.130 32.440 210.500 32.900 ;
        RECT 210.795 32.300 210.965 32.640 ;
        RECT 211.135 32.470 211.465 32.900 ;
        RECT 211.700 32.300 211.870 32.640 ;
        RECT 207.635 31.840 208.855 32.010 ;
        RECT 209.025 31.930 209.485 32.220 ;
        RECT 209.790 32.100 210.350 32.270 ;
        RECT 210.795 32.130 211.870 32.300 ;
        RECT 212.040 32.400 212.720 32.730 ;
        RECT 212.935 32.400 213.185 32.730 ;
        RECT 213.355 32.440 213.605 32.900 ;
        RECT 210.180 31.960 210.350 32.100 ;
        RECT 209.025 31.920 209.990 31.930 ;
        RECT 208.685 31.750 208.855 31.840 ;
        RECT 209.315 31.760 209.990 31.920 ;
        RECT 206.725 31.560 207.465 31.590 ;
        RECT 206.725 31.260 207.640 31.560 ;
        RECT 207.315 31.085 207.640 31.260 ;
        RECT 206.345 30.530 206.600 31.060 ;
        RECT 206.770 30.350 207.075 30.810 ;
        RECT 207.320 30.730 207.640 31.085 ;
        RECT 207.810 31.300 208.350 31.670 ;
        RECT 208.685 31.580 209.090 31.750 ;
        RECT 207.810 30.900 208.050 31.300 ;
        RECT 208.530 31.130 208.750 31.410 ;
        RECT 208.220 30.960 208.750 31.130 ;
        RECT 208.220 30.730 208.390 30.960 ;
        RECT 208.920 30.800 209.090 31.580 ;
        RECT 209.260 30.970 209.610 31.590 ;
        RECT 209.780 30.970 209.990 31.760 ;
        RECT 210.180 31.790 211.680 31.960 ;
        RECT 210.180 31.100 210.350 31.790 ;
        RECT 212.040 31.620 212.210 32.400 ;
        RECT 213.015 32.270 213.185 32.400 ;
        RECT 210.520 31.450 212.210 31.620 ;
        RECT 212.380 31.840 212.845 32.230 ;
        RECT 213.015 32.100 213.410 32.270 ;
        RECT 210.520 31.270 210.690 31.450 ;
        RECT 207.320 30.560 208.390 30.730 ;
        RECT 208.560 30.350 208.750 30.790 ;
        RECT 208.920 30.520 209.870 30.800 ;
        RECT 210.180 30.710 210.440 31.100 ;
        RECT 210.860 31.030 211.650 31.280 ;
        RECT 210.090 30.540 210.440 30.710 ;
        RECT 210.650 30.350 210.980 30.810 ;
        RECT 211.855 30.740 212.025 31.450 ;
        RECT 212.380 31.250 212.550 31.840 ;
        RECT 212.195 31.030 212.550 31.250 ;
        RECT 212.720 31.030 213.070 31.650 ;
        RECT 213.240 30.740 213.410 32.100 ;
        RECT 213.775 31.930 214.100 32.715 ;
        RECT 213.580 30.880 214.040 31.930 ;
        RECT 211.855 30.570 212.710 30.740 ;
        RECT 212.915 30.570 213.410 30.740 ;
        RECT 213.580 30.350 213.910 30.710 ;
        RECT 214.270 30.610 214.440 32.730 ;
        RECT 214.610 32.400 214.940 32.900 ;
        RECT 215.110 32.230 215.365 32.730 ;
        RECT 214.615 32.060 215.365 32.230 ;
        RECT 214.615 31.070 214.845 32.060 ;
        RECT 215.015 31.240 215.365 31.890 ;
        RECT 215.540 31.810 217.210 32.900 ;
        RECT 217.495 32.270 217.780 32.730 ;
        RECT 217.950 32.440 218.220 32.900 ;
        RECT 217.495 32.050 218.450 32.270 ;
        RECT 215.540 31.120 216.290 31.640 ;
        RECT 216.460 31.290 217.210 31.810 ;
        RECT 217.380 31.320 218.070 31.880 ;
        RECT 218.240 31.150 218.450 32.050 ;
        RECT 214.615 30.900 215.365 31.070 ;
        RECT 214.610 30.350 214.940 30.730 ;
        RECT 215.110 30.610 215.365 30.900 ;
        RECT 215.540 30.350 217.210 31.120 ;
        RECT 217.495 30.980 218.450 31.150 ;
        RECT 218.620 31.880 219.020 32.730 ;
        RECT 219.210 32.270 219.490 32.730 ;
        RECT 220.010 32.440 220.335 32.900 ;
        RECT 219.210 32.050 220.335 32.270 ;
        RECT 218.620 31.320 219.715 31.880 ;
        RECT 219.885 31.590 220.335 32.050 ;
        RECT 220.505 31.760 220.890 32.730 ;
        RECT 221.060 31.810 222.270 32.900 ;
        RECT 217.495 30.520 217.780 30.980 ;
        RECT 217.950 30.350 218.220 30.810 ;
        RECT 218.620 30.520 219.020 31.320 ;
        RECT 219.885 31.260 220.440 31.590 ;
        RECT 219.885 31.150 220.335 31.260 ;
        RECT 219.210 30.980 220.335 31.150 ;
        RECT 220.610 31.090 220.890 31.760 ;
        RECT 219.210 30.520 219.490 30.980 ;
        RECT 220.010 30.350 220.335 30.810 ;
        RECT 220.505 30.520 220.890 31.090 ;
        RECT 221.060 31.100 221.580 31.640 ;
        RECT 221.750 31.270 222.270 31.810 ;
        RECT 222.445 31.760 222.780 32.730 ;
        RECT 222.950 31.760 223.120 32.900 ;
        RECT 223.290 32.560 225.320 32.730 ;
        RECT 221.060 30.350 222.270 31.100 ;
        RECT 222.445 31.090 222.615 31.760 ;
        RECT 223.290 31.590 223.460 32.560 ;
        RECT 222.785 31.260 223.040 31.590 ;
        RECT 223.265 31.260 223.460 31.590 ;
        RECT 223.630 32.220 224.755 32.390 ;
        RECT 222.870 31.090 223.040 31.260 ;
        RECT 223.630 31.090 223.800 32.220 ;
        RECT 222.445 30.520 222.700 31.090 ;
        RECT 222.870 30.920 223.800 31.090 ;
        RECT 223.970 31.880 224.980 32.050 ;
        RECT 223.970 31.080 224.140 31.880 ;
        RECT 223.625 30.885 223.800 30.920 ;
        RECT 222.870 30.350 223.200 30.750 ;
        RECT 223.625 30.520 224.155 30.885 ;
        RECT 224.345 30.860 224.620 31.680 ;
        RECT 224.340 30.690 224.620 30.860 ;
        RECT 224.345 30.520 224.620 30.690 ;
        RECT 224.790 30.520 224.980 31.880 ;
        RECT 225.150 31.895 225.320 32.560 ;
        RECT 225.490 32.140 225.660 32.900 ;
        RECT 225.895 32.140 226.410 32.550 ;
        RECT 225.150 31.705 225.900 31.895 ;
        RECT 226.070 31.330 226.410 32.140 ;
        RECT 226.580 31.735 226.870 32.900 ;
        RECT 227.045 32.230 227.300 32.730 ;
        RECT 227.470 32.400 227.800 32.900 ;
        RECT 227.045 32.060 227.795 32.230 ;
        RECT 225.180 31.160 226.410 31.330 ;
        RECT 227.045 31.240 227.395 31.890 ;
        RECT 225.160 30.350 225.670 30.885 ;
        RECT 225.890 30.555 226.135 31.160 ;
        RECT 226.580 30.350 226.870 31.075 ;
        RECT 227.565 31.070 227.795 32.060 ;
        RECT 227.045 30.900 227.795 31.070 ;
        RECT 227.045 30.610 227.300 30.900 ;
        RECT 227.470 30.350 227.800 30.730 ;
        RECT 227.970 30.610 228.140 32.730 ;
        RECT 228.310 31.930 228.635 32.715 ;
        RECT 228.805 32.440 229.055 32.900 ;
        RECT 229.225 32.400 229.475 32.730 ;
        RECT 229.690 32.400 230.370 32.730 ;
        RECT 229.225 32.270 229.395 32.400 ;
        RECT 229.000 32.100 229.395 32.270 ;
        RECT 228.370 30.880 228.830 31.930 ;
        RECT 229.000 30.740 229.170 32.100 ;
        RECT 229.565 31.840 230.030 32.230 ;
        RECT 229.340 31.030 229.690 31.650 ;
        RECT 229.860 31.250 230.030 31.840 ;
        RECT 230.200 31.620 230.370 32.400 ;
        RECT 230.540 32.300 230.710 32.640 ;
        RECT 230.945 32.470 231.275 32.900 ;
        RECT 231.445 32.300 231.615 32.640 ;
        RECT 231.910 32.440 232.280 32.900 ;
        RECT 230.540 32.130 231.615 32.300 ;
        RECT 232.450 32.270 232.620 32.730 ;
        RECT 232.855 32.390 233.725 32.730 ;
        RECT 233.895 32.440 234.145 32.900 ;
        RECT 232.060 32.100 232.620 32.270 ;
        RECT 232.060 31.960 232.230 32.100 ;
        RECT 230.730 31.790 232.230 31.960 ;
        RECT 232.925 31.930 233.385 32.220 ;
        RECT 230.200 31.450 231.890 31.620 ;
        RECT 229.860 31.030 230.215 31.250 ;
        RECT 230.385 30.740 230.555 31.450 ;
        RECT 230.760 31.030 231.550 31.280 ;
        RECT 231.720 31.270 231.890 31.450 ;
        RECT 232.060 31.100 232.230 31.790 ;
        RECT 228.500 30.350 228.830 30.710 ;
        RECT 229.000 30.570 229.495 30.740 ;
        RECT 229.700 30.570 230.555 30.740 ;
        RECT 231.430 30.350 231.760 30.810 ;
        RECT 231.970 30.710 232.230 31.100 ;
        RECT 232.420 31.920 233.385 31.930 ;
        RECT 233.555 32.010 233.725 32.390 ;
        RECT 234.315 32.350 234.485 32.640 ;
        RECT 234.665 32.520 234.995 32.900 ;
        RECT 234.315 32.180 235.115 32.350 ;
        RECT 232.420 31.760 233.095 31.920 ;
        RECT 233.555 31.840 234.775 32.010 ;
        RECT 232.420 30.970 232.630 31.760 ;
        RECT 233.555 31.750 233.725 31.840 ;
        RECT 232.800 30.970 233.150 31.590 ;
        RECT 233.320 31.580 233.725 31.750 ;
        RECT 233.320 30.800 233.490 31.580 ;
        RECT 233.660 31.130 233.880 31.410 ;
        RECT 234.060 31.300 234.600 31.670 ;
        RECT 234.945 31.590 235.115 32.180 ;
        RECT 235.335 31.760 235.640 32.900 ;
        RECT 235.810 31.710 236.065 32.590 ;
        RECT 234.945 31.560 235.685 31.590 ;
        RECT 233.660 30.960 234.190 31.130 ;
        RECT 231.970 30.540 232.320 30.710 ;
        RECT 232.540 30.520 233.490 30.800 ;
        RECT 233.660 30.350 233.850 30.790 ;
        RECT 234.020 30.730 234.190 30.960 ;
        RECT 234.360 30.900 234.600 31.300 ;
        RECT 234.770 31.260 235.685 31.560 ;
        RECT 234.770 31.085 235.095 31.260 ;
        RECT 234.770 30.730 235.090 31.085 ;
        RECT 235.855 31.060 236.065 31.710 ;
        RECT 234.020 30.560 235.090 30.730 ;
        RECT 235.335 30.350 235.640 30.810 ;
        RECT 235.810 30.530 236.065 31.060 ;
        RECT 236.240 31.760 236.625 32.730 ;
        RECT 236.795 32.440 237.120 32.900 ;
        RECT 237.640 32.270 237.920 32.730 ;
        RECT 236.795 32.050 237.920 32.270 ;
        RECT 236.240 31.090 236.520 31.760 ;
        RECT 236.795 31.590 237.245 32.050 ;
        RECT 238.110 31.880 238.510 32.730 ;
        RECT 238.910 32.440 239.180 32.900 ;
        RECT 239.350 32.270 239.635 32.730 ;
        RECT 236.690 31.260 237.245 31.590 ;
        RECT 237.415 31.320 238.510 31.880 ;
        RECT 236.795 31.150 237.245 31.260 ;
        RECT 236.240 30.520 236.625 31.090 ;
        RECT 236.795 30.980 237.920 31.150 ;
        RECT 236.795 30.350 237.120 30.810 ;
        RECT 237.640 30.520 237.920 30.980 ;
        RECT 238.110 30.520 238.510 31.320 ;
        RECT 238.680 32.050 239.635 32.270 ;
        RECT 238.680 31.150 238.890 32.050 ;
        RECT 239.975 32.030 240.260 32.900 ;
        RECT 240.430 32.270 240.690 32.730 ;
        RECT 240.865 32.440 241.120 32.900 ;
        RECT 241.290 32.270 241.550 32.730 ;
        RECT 240.430 32.100 241.550 32.270 ;
        RECT 241.720 32.100 242.030 32.900 ;
        RECT 239.060 31.320 239.750 31.880 ;
        RECT 240.430 31.850 240.690 32.100 ;
        RECT 242.200 31.930 242.510 32.730 ;
        RECT 242.685 32.475 243.020 32.900 ;
        RECT 243.190 32.295 243.375 32.700 ;
        RECT 239.935 31.680 240.690 31.850 ;
        RECT 241.480 31.760 242.510 31.930 ;
        RECT 239.935 31.170 240.340 31.680 ;
        RECT 241.480 31.510 241.650 31.760 ;
        RECT 240.510 31.340 241.650 31.510 ;
        RECT 238.680 30.980 239.635 31.150 ;
        RECT 239.935 31.000 241.585 31.170 ;
        RECT 241.820 31.020 242.170 31.590 ;
        RECT 238.910 30.350 239.180 30.810 ;
        RECT 239.350 30.520 239.635 30.980 ;
        RECT 239.980 30.350 240.260 30.830 ;
        RECT 240.430 30.610 240.690 31.000 ;
        RECT 240.865 30.350 241.120 30.830 ;
        RECT 241.290 30.610 241.585 31.000 ;
        RECT 242.340 30.850 242.510 31.760 ;
        RECT 242.710 32.120 243.375 32.295 ;
        RECT 243.580 32.120 243.910 32.900 ;
        RECT 242.710 31.090 243.050 32.120 ;
        RECT 244.080 31.930 244.350 32.700 ;
        RECT 244.520 32.465 249.865 32.900 ;
        RECT 243.220 31.760 244.350 31.930 ;
        RECT 243.220 31.260 243.470 31.760 ;
        RECT 242.710 30.920 243.395 31.090 ;
        RECT 243.650 31.010 244.010 31.590 ;
        RECT 241.765 30.350 242.040 30.830 ;
        RECT 242.210 30.520 242.510 30.850 ;
        RECT 242.685 30.350 243.020 30.750 ;
        RECT 243.190 30.520 243.395 30.920 ;
        RECT 244.180 30.850 244.350 31.760 ;
        RECT 246.105 30.895 246.445 31.725 ;
        RECT 247.925 31.215 248.275 32.465 ;
        RECT 250.040 31.810 251.710 32.900 ;
        RECT 250.040 31.120 250.790 31.640 ;
        RECT 250.960 31.290 251.710 31.810 ;
        RECT 252.340 31.735 252.630 32.900 ;
        RECT 252.800 32.465 258.145 32.900 ;
        RECT 243.605 30.350 243.880 30.830 ;
        RECT 244.090 30.520 244.350 30.850 ;
        RECT 244.520 30.350 249.865 30.895 ;
        RECT 250.040 30.350 251.710 31.120 ;
        RECT 252.340 30.350 252.630 31.075 ;
        RECT 254.385 30.895 254.725 31.725 ;
        RECT 256.205 31.215 256.555 32.465 ;
        RECT 258.320 31.810 259.990 32.900 ;
        RECT 258.320 31.120 259.070 31.640 ;
        RECT 259.240 31.290 259.990 31.810 ;
        RECT 260.160 31.760 260.440 32.900 ;
        RECT 260.610 31.750 260.940 32.730 ;
        RECT 261.110 31.760 261.370 32.900 ;
        RECT 261.540 32.465 266.885 32.900 ;
        RECT 267.060 32.465 272.405 32.900 ;
        RECT 272.580 32.465 277.925 32.900 ;
        RECT 260.170 31.320 260.505 31.590 ;
        RECT 260.675 31.150 260.845 31.750 ;
        RECT 261.015 31.340 261.350 31.590 ;
        RECT 252.800 30.350 258.145 30.895 ;
        RECT 258.320 30.350 259.990 31.120 ;
        RECT 260.160 30.350 260.470 31.150 ;
        RECT 260.675 30.520 261.370 31.150 ;
        RECT 263.125 30.895 263.465 31.725 ;
        RECT 264.945 31.215 265.295 32.465 ;
        RECT 268.645 30.895 268.985 31.725 ;
        RECT 270.465 31.215 270.815 32.465 ;
        RECT 274.165 30.895 274.505 31.725 ;
        RECT 275.985 31.215 276.335 32.465 ;
        RECT 278.100 31.735 278.390 32.900 ;
        RECT 278.560 32.465 283.905 32.900 ;
        RECT 284.080 32.465 289.425 32.900 ;
        RECT 289.600 32.465 294.945 32.900 ;
        RECT 295.120 32.465 300.465 32.900 ;
        RECT 261.540 30.350 266.885 30.895 ;
        RECT 267.060 30.350 272.405 30.895 ;
        RECT 272.580 30.350 277.925 30.895 ;
        RECT 278.100 30.350 278.390 31.075 ;
        RECT 280.145 30.895 280.485 31.725 ;
        RECT 281.965 31.215 282.315 32.465 ;
        RECT 285.665 30.895 286.005 31.725 ;
        RECT 287.485 31.215 287.835 32.465 ;
        RECT 291.185 30.895 291.525 31.725 ;
        RECT 293.005 31.215 293.355 32.465 ;
        RECT 296.705 30.895 297.045 31.725 ;
        RECT 298.525 31.215 298.875 32.465 ;
        RECT 300.640 31.810 303.230 32.900 ;
        RECT 300.640 31.120 301.850 31.640 ;
        RECT 302.020 31.290 303.230 31.810 ;
        RECT 303.860 31.735 304.150 32.900 ;
        RECT 304.320 32.465 309.665 32.900 ;
        RECT 278.560 30.350 283.905 30.895 ;
        RECT 284.080 30.350 289.425 30.895 ;
        RECT 289.600 30.350 294.945 30.895 ;
        RECT 295.120 30.350 300.465 30.895 ;
        RECT 300.640 30.350 303.230 31.120 ;
        RECT 303.860 30.350 304.150 31.075 ;
        RECT 305.905 30.895 306.245 31.725 ;
        RECT 307.725 31.215 308.075 32.465 ;
        RECT 309.840 31.810 311.050 32.900 ;
        RECT 309.840 31.270 310.360 31.810 ;
        RECT 310.530 31.100 311.050 31.640 ;
        RECT 304.320 30.350 309.665 30.895 ;
        RECT 309.840 30.350 311.050 31.100 ;
        RECT 162.095 30.180 311.135 30.350 ;
        RECT 162.180 29.430 163.390 30.180 ;
        RECT 162.180 28.890 162.700 29.430 ;
        RECT 163.565 29.340 163.825 30.180 ;
        RECT 164.000 29.435 164.255 30.010 ;
        RECT 164.425 29.800 164.755 30.180 ;
        RECT 164.970 29.630 165.140 30.010 ;
        RECT 165.400 29.635 170.745 30.180 ;
        RECT 164.425 29.460 165.140 29.630 ;
        RECT 162.870 28.720 163.390 29.260 ;
        RECT 162.180 27.630 163.390 28.720 ;
        RECT 163.565 27.630 163.825 28.780 ;
        RECT 164.000 28.705 164.170 29.435 ;
        RECT 164.425 29.270 164.595 29.460 ;
        RECT 164.340 28.940 164.595 29.270 ;
        RECT 164.425 28.730 164.595 28.940 ;
        RECT 164.875 28.910 165.230 29.280 ;
        RECT 166.985 28.805 167.325 29.635 ;
        RECT 170.920 29.410 174.430 30.180 ;
        RECT 175.175 29.550 175.460 30.010 ;
        RECT 175.630 29.720 175.900 30.180 ;
        RECT 164.000 27.800 164.255 28.705 ;
        RECT 164.425 28.560 165.140 28.730 ;
        RECT 164.425 27.630 164.755 28.390 ;
        RECT 164.970 27.800 165.140 28.560 ;
        RECT 168.805 28.065 169.155 29.315 ;
        RECT 170.920 28.890 172.570 29.410 ;
        RECT 175.175 29.380 176.130 29.550 ;
        RECT 172.740 28.720 174.430 29.240 ;
        RECT 165.400 27.630 170.745 28.065 ;
        RECT 170.920 27.630 174.430 28.720 ;
        RECT 175.060 28.650 175.750 29.210 ;
        RECT 175.920 28.480 176.130 29.380 ;
        RECT 175.175 28.260 176.130 28.480 ;
        RECT 176.300 29.210 176.700 30.010 ;
        RECT 176.890 29.550 177.170 30.010 ;
        RECT 177.690 29.720 178.015 30.180 ;
        RECT 176.890 29.380 178.015 29.550 ;
        RECT 178.185 29.440 178.570 30.010 ;
        RECT 177.565 29.270 178.015 29.380 ;
        RECT 176.300 28.650 177.395 29.210 ;
        RECT 177.565 28.940 178.120 29.270 ;
        RECT 175.175 27.800 175.460 28.260 ;
        RECT 175.630 27.630 175.900 28.090 ;
        RECT 176.300 27.800 176.700 28.650 ;
        RECT 177.565 28.480 178.015 28.940 ;
        RECT 178.290 28.770 178.570 29.440 ;
        RECT 176.890 28.260 178.015 28.480 ;
        RECT 176.890 27.800 177.170 28.260 ;
        RECT 177.690 27.630 178.015 28.090 ;
        RECT 178.185 27.800 178.570 28.770 ;
        RECT 178.745 29.470 179.000 30.000 ;
        RECT 179.170 29.720 179.475 30.180 ;
        RECT 179.720 29.800 180.790 29.970 ;
        RECT 178.745 28.820 178.955 29.470 ;
        RECT 179.720 29.445 180.040 29.800 ;
        RECT 179.715 29.270 180.040 29.445 ;
        RECT 179.125 28.970 180.040 29.270 ;
        RECT 180.210 29.230 180.450 29.630 ;
        RECT 180.620 29.570 180.790 29.800 ;
        RECT 180.960 29.740 181.150 30.180 ;
        RECT 181.320 29.730 182.270 30.010 ;
        RECT 182.490 29.820 182.840 29.990 ;
        RECT 180.620 29.400 181.150 29.570 ;
        RECT 179.125 28.940 179.865 28.970 ;
        RECT 178.745 27.940 179.000 28.820 ;
        RECT 179.170 27.630 179.475 28.770 ;
        RECT 179.695 28.350 179.865 28.940 ;
        RECT 180.210 28.860 180.750 29.230 ;
        RECT 180.930 29.120 181.150 29.400 ;
        RECT 181.320 28.950 181.490 29.730 ;
        RECT 181.085 28.780 181.490 28.950 ;
        RECT 181.660 28.940 182.010 29.560 ;
        RECT 181.085 28.690 181.255 28.780 ;
        RECT 182.180 28.770 182.390 29.560 ;
        RECT 180.035 28.520 181.255 28.690 ;
        RECT 181.715 28.610 182.390 28.770 ;
        RECT 179.695 28.180 180.495 28.350 ;
        RECT 179.815 27.630 180.145 28.010 ;
        RECT 180.325 27.890 180.495 28.180 ;
        RECT 181.085 28.140 181.255 28.520 ;
        RECT 181.425 28.600 182.390 28.610 ;
        RECT 182.580 29.430 182.840 29.820 ;
        RECT 183.050 29.720 183.380 30.180 ;
        RECT 184.255 29.790 185.110 29.960 ;
        RECT 185.315 29.790 185.810 29.960 ;
        RECT 185.980 29.820 186.310 30.180 ;
        RECT 182.580 28.740 182.750 29.430 ;
        RECT 182.920 29.080 183.090 29.260 ;
        RECT 183.260 29.250 184.050 29.500 ;
        RECT 184.255 29.080 184.425 29.790 ;
        RECT 184.595 29.280 184.950 29.500 ;
        RECT 182.920 28.910 184.610 29.080 ;
        RECT 181.425 28.310 181.885 28.600 ;
        RECT 182.580 28.570 184.080 28.740 ;
        RECT 182.580 28.430 182.750 28.570 ;
        RECT 182.190 28.260 182.750 28.430 ;
        RECT 180.665 27.630 180.915 28.090 ;
        RECT 181.085 27.800 181.955 28.140 ;
        RECT 182.190 27.800 182.360 28.260 ;
        RECT 183.195 28.230 184.270 28.400 ;
        RECT 182.530 27.630 182.900 28.090 ;
        RECT 183.195 27.890 183.365 28.230 ;
        RECT 183.535 27.630 183.865 28.060 ;
        RECT 184.100 27.890 184.270 28.230 ;
        RECT 184.440 28.130 184.610 28.910 ;
        RECT 184.780 28.690 184.950 29.280 ;
        RECT 185.120 28.880 185.470 29.500 ;
        RECT 184.780 28.300 185.245 28.690 ;
        RECT 185.640 28.430 185.810 29.790 ;
        RECT 185.980 28.600 186.440 29.650 ;
        RECT 185.415 28.260 185.810 28.430 ;
        RECT 185.415 28.130 185.585 28.260 ;
        RECT 184.440 27.800 185.120 28.130 ;
        RECT 185.335 27.800 185.585 28.130 ;
        RECT 185.755 27.630 186.005 28.090 ;
        RECT 186.175 27.815 186.500 28.600 ;
        RECT 186.670 27.800 186.840 29.920 ;
        RECT 187.010 29.800 187.340 30.180 ;
        RECT 187.510 29.630 187.765 29.920 ;
        RECT 187.015 29.460 187.765 29.630 ;
        RECT 187.015 28.470 187.245 29.460 ;
        RECT 187.940 29.455 188.230 30.180 ;
        RECT 188.400 29.635 193.745 30.180 ;
        RECT 187.415 28.640 187.765 29.290 ;
        RECT 189.985 28.805 190.325 29.635 ;
        RECT 193.920 29.410 195.590 30.180 ;
        RECT 195.765 29.470 196.020 30.000 ;
        RECT 196.190 29.720 196.495 30.180 ;
        RECT 196.740 29.800 197.810 29.970 ;
        RECT 187.015 28.300 187.765 28.470 ;
        RECT 187.010 27.630 187.340 28.130 ;
        RECT 187.510 27.800 187.765 28.300 ;
        RECT 187.940 27.630 188.230 28.795 ;
        RECT 191.805 28.065 192.155 29.315 ;
        RECT 193.920 28.890 194.670 29.410 ;
        RECT 194.840 28.720 195.590 29.240 ;
        RECT 188.400 27.630 193.745 28.065 ;
        RECT 193.920 27.630 195.590 28.720 ;
        RECT 195.765 28.820 195.975 29.470 ;
        RECT 196.740 29.445 197.060 29.800 ;
        RECT 196.735 29.270 197.060 29.445 ;
        RECT 196.145 28.970 197.060 29.270 ;
        RECT 197.230 29.230 197.470 29.630 ;
        RECT 197.640 29.570 197.810 29.800 ;
        RECT 197.980 29.740 198.170 30.180 ;
        RECT 198.340 29.730 199.290 30.010 ;
        RECT 199.510 29.820 199.860 29.990 ;
        RECT 197.640 29.400 198.170 29.570 ;
        RECT 196.145 28.940 196.885 28.970 ;
        RECT 195.765 27.940 196.020 28.820 ;
        RECT 196.190 27.630 196.495 28.770 ;
        RECT 196.715 28.350 196.885 28.940 ;
        RECT 197.230 28.860 197.770 29.230 ;
        RECT 197.950 29.120 198.170 29.400 ;
        RECT 198.340 28.950 198.510 29.730 ;
        RECT 198.105 28.780 198.510 28.950 ;
        RECT 198.680 28.940 199.030 29.560 ;
        RECT 198.105 28.690 198.275 28.780 ;
        RECT 199.200 28.770 199.410 29.560 ;
        RECT 197.055 28.520 198.275 28.690 ;
        RECT 198.735 28.610 199.410 28.770 ;
        RECT 196.715 28.180 197.515 28.350 ;
        RECT 196.835 27.630 197.165 28.010 ;
        RECT 197.345 27.890 197.515 28.180 ;
        RECT 198.105 28.140 198.275 28.520 ;
        RECT 198.445 28.600 199.410 28.610 ;
        RECT 199.600 29.430 199.860 29.820 ;
        RECT 200.070 29.720 200.400 30.180 ;
        RECT 201.275 29.790 202.130 29.960 ;
        RECT 202.335 29.790 202.830 29.960 ;
        RECT 203.000 29.820 203.330 30.180 ;
        RECT 199.600 28.740 199.770 29.430 ;
        RECT 199.940 29.080 200.110 29.260 ;
        RECT 200.280 29.250 201.070 29.500 ;
        RECT 201.275 29.080 201.445 29.790 ;
        RECT 201.615 29.280 201.970 29.500 ;
        RECT 199.940 28.910 201.630 29.080 ;
        RECT 198.445 28.310 198.905 28.600 ;
        RECT 199.600 28.570 201.100 28.740 ;
        RECT 199.600 28.430 199.770 28.570 ;
        RECT 199.210 28.260 199.770 28.430 ;
        RECT 197.685 27.630 197.935 28.090 ;
        RECT 198.105 27.800 198.975 28.140 ;
        RECT 199.210 27.800 199.380 28.260 ;
        RECT 200.215 28.230 201.290 28.400 ;
        RECT 199.550 27.630 199.920 28.090 ;
        RECT 200.215 27.890 200.385 28.230 ;
        RECT 200.555 27.630 200.885 28.060 ;
        RECT 201.120 27.890 201.290 28.230 ;
        RECT 201.460 28.130 201.630 28.910 ;
        RECT 201.800 28.690 201.970 29.280 ;
        RECT 202.140 28.880 202.490 29.500 ;
        RECT 201.800 28.300 202.265 28.690 ;
        RECT 202.660 28.430 202.830 29.790 ;
        RECT 203.000 28.600 203.460 29.650 ;
        RECT 202.435 28.260 202.830 28.430 ;
        RECT 202.435 28.130 202.605 28.260 ;
        RECT 201.460 27.800 202.140 28.130 ;
        RECT 202.355 27.800 202.605 28.130 ;
        RECT 202.775 27.630 203.025 28.090 ;
        RECT 203.195 27.815 203.520 28.600 ;
        RECT 203.690 27.800 203.860 29.920 ;
        RECT 204.030 29.800 204.360 30.180 ;
        RECT 204.530 29.630 204.785 29.920 ;
        RECT 204.035 29.460 204.785 29.630 ;
        RECT 204.035 28.470 204.265 29.460 ;
        RECT 204.960 29.440 205.345 30.010 ;
        RECT 205.515 29.720 205.840 30.180 ;
        RECT 206.360 29.550 206.640 30.010 ;
        RECT 204.435 28.640 204.785 29.290 ;
        RECT 204.960 28.770 205.240 29.440 ;
        RECT 205.515 29.380 206.640 29.550 ;
        RECT 205.515 29.270 205.965 29.380 ;
        RECT 205.410 28.940 205.965 29.270 ;
        RECT 206.830 29.210 207.230 30.010 ;
        RECT 207.630 29.720 207.900 30.180 ;
        RECT 208.070 29.550 208.355 30.010 ;
        RECT 204.035 28.300 204.785 28.470 ;
        RECT 204.030 27.630 204.360 28.130 ;
        RECT 204.530 27.800 204.785 28.300 ;
        RECT 204.960 27.800 205.345 28.770 ;
        RECT 205.515 28.480 205.965 28.940 ;
        RECT 206.135 28.650 207.230 29.210 ;
        RECT 205.515 28.260 206.640 28.480 ;
        RECT 205.515 27.630 205.840 28.090 ;
        RECT 206.360 27.800 206.640 28.260 ;
        RECT 206.830 27.800 207.230 28.650 ;
        RECT 207.400 29.380 208.355 29.550 ;
        RECT 208.640 29.410 212.150 30.180 ;
        RECT 212.320 29.430 213.530 30.180 ;
        RECT 213.700 29.455 213.990 30.180 ;
        RECT 214.160 29.635 219.505 30.180 ;
        RECT 219.680 29.635 225.025 30.180 ;
        RECT 225.200 29.635 230.545 30.180 ;
        RECT 207.400 28.480 207.610 29.380 ;
        RECT 207.780 28.650 208.470 29.210 ;
        RECT 208.640 28.890 210.290 29.410 ;
        RECT 210.460 28.720 212.150 29.240 ;
        RECT 212.320 28.890 212.840 29.430 ;
        RECT 213.010 28.720 213.530 29.260 ;
        RECT 215.745 28.805 216.085 29.635 ;
        RECT 207.400 28.260 208.355 28.480 ;
        RECT 207.630 27.630 207.900 28.090 ;
        RECT 208.070 27.800 208.355 28.260 ;
        RECT 208.640 27.630 212.150 28.720 ;
        RECT 212.320 27.630 213.530 28.720 ;
        RECT 213.700 27.630 213.990 28.795 ;
        RECT 217.565 28.065 217.915 29.315 ;
        RECT 221.265 28.805 221.605 29.635 ;
        RECT 223.085 28.065 223.435 29.315 ;
        RECT 226.785 28.805 227.125 29.635 ;
        RECT 231.640 29.440 232.025 30.010 ;
        RECT 232.195 29.720 232.520 30.180 ;
        RECT 233.040 29.550 233.320 30.010 ;
        RECT 228.605 28.065 228.955 29.315 ;
        RECT 231.640 28.770 231.920 29.440 ;
        RECT 232.195 29.380 233.320 29.550 ;
        RECT 232.195 29.270 232.645 29.380 ;
        RECT 232.090 28.940 232.645 29.270 ;
        RECT 233.510 29.210 233.910 30.010 ;
        RECT 234.310 29.720 234.580 30.180 ;
        RECT 234.750 29.550 235.035 30.010 ;
        RECT 214.160 27.630 219.505 28.065 ;
        RECT 219.680 27.630 225.025 28.065 ;
        RECT 225.200 27.630 230.545 28.065 ;
        RECT 231.640 27.800 232.025 28.770 ;
        RECT 232.195 28.480 232.645 28.940 ;
        RECT 232.815 28.650 233.910 29.210 ;
        RECT 232.195 28.260 233.320 28.480 ;
        RECT 232.195 27.630 232.520 28.090 ;
        RECT 233.040 27.800 233.320 28.260 ;
        RECT 233.510 27.800 233.910 28.650 ;
        RECT 234.080 29.380 235.035 29.550 ;
        RECT 235.320 29.410 238.830 30.180 ;
        RECT 239.460 29.455 239.750 30.180 ;
        RECT 239.920 29.635 245.265 30.180 ;
        RECT 245.440 29.635 250.785 30.180 ;
        RECT 250.960 29.635 256.305 30.180 ;
        RECT 256.480 29.635 261.825 30.180 ;
        RECT 234.080 28.480 234.290 29.380 ;
        RECT 234.460 28.650 235.150 29.210 ;
        RECT 235.320 28.890 236.970 29.410 ;
        RECT 237.140 28.720 238.830 29.240 ;
        RECT 241.505 28.805 241.845 29.635 ;
        RECT 234.080 28.260 235.035 28.480 ;
        RECT 234.310 27.630 234.580 28.090 ;
        RECT 234.750 27.800 235.035 28.260 ;
        RECT 235.320 27.630 238.830 28.720 ;
        RECT 239.460 27.630 239.750 28.795 ;
        RECT 243.325 28.065 243.675 29.315 ;
        RECT 247.025 28.805 247.365 29.635 ;
        RECT 248.845 28.065 249.195 29.315 ;
        RECT 252.545 28.805 252.885 29.635 ;
        RECT 254.365 28.065 254.715 29.315 ;
        RECT 258.065 28.805 258.405 29.635 ;
        RECT 262.000 29.410 264.590 30.180 ;
        RECT 265.220 29.455 265.510 30.180 ;
        RECT 265.680 29.635 271.025 30.180 ;
        RECT 271.200 29.635 276.545 30.180 ;
        RECT 276.720 29.635 282.065 30.180 ;
        RECT 282.240 29.635 287.585 30.180 ;
        RECT 259.885 28.065 260.235 29.315 ;
        RECT 262.000 28.890 263.210 29.410 ;
        RECT 263.380 28.720 264.590 29.240 ;
        RECT 267.265 28.805 267.605 29.635 ;
        RECT 239.920 27.630 245.265 28.065 ;
        RECT 245.440 27.630 250.785 28.065 ;
        RECT 250.960 27.630 256.305 28.065 ;
        RECT 256.480 27.630 261.825 28.065 ;
        RECT 262.000 27.630 264.590 28.720 ;
        RECT 265.220 27.630 265.510 28.795 ;
        RECT 269.085 28.065 269.435 29.315 ;
        RECT 272.785 28.805 273.125 29.635 ;
        RECT 274.605 28.065 274.955 29.315 ;
        RECT 278.305 28.805 278.645 29.635 ;
        RECT 280.125 28.065 280.475 29.315 ;
        RECT 283.825 28.805 284.165 29.635 ;
        RECT 287.760 29.410 290.350 30.180 ;
        RECT 290.980 29.455 291.270 30.180 ;
        RECT 291.440 29.635 296.785 30.180 ;
        RECT 296.960 29.635 302.305 30.180 ;
        RECT 302.480 29.635 307.825 30.180 ;
        RECT 285.645 28.065 285.995 29.315 ;
        RECT 287.760 28.890 288.970 29.410 ;
        RECT 289.140 28.720 290.350 29.240 ;
        RECT 293.025 28.805 293.365 29.635 ;
        RECT 265.680 27.630 271.025 28.065 ;
        RECT 271.200 27.630 276.545 28.065 ;
        RECT 276.720 27.630 282.065 28.065 ;
        RECT 282.240 27.630 287.585 28.065 ;
        RECT 287.760 27.630 290.350 28.720 ;
        RECT 290.980 27.630 291.270 28.795 ;
        RECT 294.845 28.065 295.195 29.315 ;
        RECT 298.545 28.805 298.885 29.635 ;
        RECT 300.365 28.065 300.715 29.315 ;
        RECT 304.065 28.805 304.405 29.635 ;
        RECT 308.000 29.410 309.670 30.180 ;
        RECT 309.840 29.430 311.050 30.180 ;
        RECT 305.885 28.065 306.235 29.315 ;
        RECT 308.000 28.890 308.750 29.410 ;
        RECT 308.920 28.720 309.670 29.240 ;
        RECT 291.440 27.630 296.785 28.065 ;
        RECT 296.960 27.630 302.305 28.065 ;
        RECT 302.480 27.630 307.825 28.065 ;
        RECT 308.000 27.630 309.670 28.720 ;
        RECT 309.840 28.720 310.360 29.260 ;
        RECT 310.530 28.890 311.050 29.430 ;
        RECT 309.840 27.630 311.050 28.720 ;
        RECT 162.095 27.460 311.135 27.630 ;
        RECT 162.180 26.370 163.390 27.460 ;
        RECT 163.560 27.025 168.905 27.460 ;
        RECT 169.080 27.025 174.425 27.460 ;
        RECT 162.180 25.660 162.700 26.200 ;
        RECT 162.870 25.830 163.390 26.370 ;
        RECT 162.180 24.910 163.390 25.660 ;
        RECT 165.145 25.455 165.485 26.285 ;
        RECT 166.965 25.775 167.315 27.025 ;
        RECT 170.665 25.455 171.005 26.285 ;
        RECT 172.485 25.775 172.835 27.025 ;
        RECT 175.060 26.295 175.350 27.460 ;
        RECT 175.520 26.370 178.110 27.460 ;
        RECT 175.520 25.680 176.730 26.200 ;
        RECT 176.900 25.850 178.110 26.370 ;
        RECT 178.280 26.320 178.665 27.290 ;
        RECT 178.835 27.000 179.160 27.460 ;
        RECT 179.680 26.830 179.960 27.290 ;
        RECT 178.835 26.610 179.960 26.830 ;
        RECT 163.560 24.910 168.905 25.455 ;
        RECT 169.080 24.910 174.425 25.455 ;
        RECT 175.060 24.910 175.350 25.635 ;
        RECT 175.520 24.910 178.110 25.680 ;
        RECT 178.280 25.650 178.560 26.320 ;
        RECT 178.835 26.150 179.285 26.610 ;
        RECT 180.150 26.440 180.550 27.290 ;
        RECT 180.950 27.000 181.220 27.460 ;
        RECT 181.390 26.830 181.675 27.290 ;
        RECT 178.730 25.820 179.285 26.150 ;
        RECT 179.455 25.880 180.550 26.440 ;
        RECT 178.835 25.710 179.285 25.820 ;
        RECT 178.280 25.080 178.665 25.650 ;
        RECT 178.835 25.540 179.960 25.710 ;
        RECT 178.835 24.910 179.160 25.370 ;
        RECT 179.680 25.080 179.960 25.540 ;
        RECT 180.150 25.080 180.550 25.880 ;
        RECT 180.720 26.610 181.675 26.830 ;
        RECT 180.720 25.710 180.930 26.610 ;
        RECT 181.100 25.880 181.790 26.440 ;
        RECT 181.960 26.370 183.170 27.460 ;
        RECT 183.455 26.830 183.740 27.290 ;
        RECT 183.910 27.000 184.180 27.460 ;
        RECT 183.455 26.610 184.410 26.830 ;
        RECT 180.720 25.540 181.675 25.710 ;
        RECT 180.950 24.910 181.220 25.370 ;
        RECT 181.390 25.080 181.675 25.540 ;
        RECT 181.960 25.660 182.480 26.200 ;
        RECT 182.650 25.830 183.170 26.370 ;
        RECT 183.340 25.880 184.030 26.440 ;
        RECT 184.200 25.710 184.410 26.610 ;
        RECT 181.960 24.910 183.170 25.660 ;
        RECT 183.455 25.540 184.410 25.710 ;
        RECT 184.580 26.440 184.980 27.290 ;
        RECT 185.170 26.830 185.450 27.290 ;
        RECT 185.970 27.000 186.295 27.460 ;
        RECT 185.170 26.610 186.295 26.830 ;
        RECT 184.580 25.880 185.675 26.440 ;
        RECT 185.845 26.150 186.295 26.610 ;
        RECT 186.465 26.320 186.850 27.290 ;
        RECT 187.020 27.025 192.365 27.460 ;
        RECT 192.540 27.025 197.885 27.460 ;
        RECT 183.455 25.080 183.740 25.540 ;
        RECT 183.910 24.910 184.180 25.370 ;
        RECT 184.580 25.080 184.980 25.880 ;
        RECT 185.845 25.820 186.400 26.150 ;
        RECT 185.845 25.710 186.295 25.820 ;
        RECT 185.170 25.540 186.295 25.710 ;
        RECT 186.570 25.650 186.850 26.320 ;
        RECT 185.170 25.080 185.450 25.540 ;
        RECT 185.970 24.910 186.295 25.370 ;
        RECT 186.465 25.080 186.850 25.650 ;
        RECT 188.605 25.455 188.945 26.285 ;
        RECT 190.425 25.775 190.775 27.025 ;
        RECT 194.125 25.455 194.465 26.285 ;
        RECT 195.945 25.775 196.295 27.025 ;
        RECT 198.060 26.370 200.650 27.460 ;
        RECT 198.060 25.680 199.270 26.200 ;
        RECT 199.440 25.850 200.650 26.370 ;
        RECT 200.820 26.295 201.110 27.460 ;
        RECT 201.280 27.025 206.625 27.460 ;
        RECT 206.800 27.025 212.145 27.460 ;
        RECT 212.320 27.025 217.665 27.460 ;
        RECT 217.840 27.025 223.185 27.460 ;
        RECT 187.020 24.910 192.365 25.455 ;
        RECT 192.540 24.910 197.885 25.455 ;
        RECT 198.060 24.910 200.650 25.680 ;
        RECT 200.820 24.910 201.110 25.635 ;
        RECT 202.865 25.455 203.205 26.285 ;
        RECT 204.685 25.775 205.035 27.025 ;
        RECT 208.385 25.455 208.725 26.285 ;
        RECT 210.205 25.775 210.555 27.025 ;
        RECT 213.905 25.455 214.245 26.285 ;
        RECT 215.725 25.775 216.075 27.025 ;
        RECT 219.425 25.455 219.765 26.285 ;
        RECT 221.245 25.775 221.595 27.025 ;
        RECT 223.360 26.370 225.950 27.460 ;
        RECT 223.360 25.680 224.570 26.200 ;
        RECT 224.740 25.850 225.950 26.370 ;
        RECT 226.580 26.295 226.870 27.460 ;
        RECT 227.040 27.025 232.385 27.460 ;
        RECT 232.560 27.025 237.905 27.460 ;
        RECT 238.080 27.025 243.425 27.460 ;
        RECT 243.600 27.025 248.945 27.460 ;
        RECT 201.280 24.910 206.625 25.455 ;
        RECT 206.800 24.910 212.145 25.455 ;
        RECT 212.320 24.910 217.665 25.455 ;
        RECT 217.840 24.910 223.185 25.455 ;
        RECT 223.360 24.910 225.950 25.680 ;
        RECT 226.580 24.910 226.870 25.635 ;
        RECT 228.625 25.455 228.965 26.285 ;
        RECT 230.445 25.775 230.795 27.025 ;
        RECT 234.145 25.455 234.485 26.285 ;
        RECT 235.965 25.775 236.315 27.025 ;
        RECT 239.665 25.455 240.005 26.285 ;
        RECT 241.485 25.775 241.835 27.025 ;
        RECT 245.185 25.455 245.525 26.285 ;
        RECT 247.005 25.775 247.355 27.025 ;
        RECT 249.120 26.370 251.710 27.460 ;
        RECT 249.120 25.680 250.330 26.200 ;
        RECT 250.500 25.850 251.710 26.370 ;
        RECT 252.340 26.295 252.630 27.460 ;
        RECT 252.800 27.025 258.145 27.460 ;
        RECT 258.320 27.025 263.665 27.460 ;
        RECT 263.840 27.025 269.185 27.460 ;
        RECT 269.360 27.025 274.705 27.460 ;
        RECT 227.040 24.910 232.385 25.455 ;
        RECT 232.560 24.910 237.905 25.455 ;
        RECT 238.080 24.910 243.425 25.455 ;
        RECT 243.600 24.910 248.945 25.455 ;
        RECT 249.120 24.910 251.710 25.680 ;
        RECT 252.340 24.910 252.630 25.635 ;
        RECT 254.385 25.455 254.725 26.285 ;
        RECT 256.205 25.775 256.555 27.025 ;
        RECT 259.905 25.455 260.245 26.285 ;
        RECT 261.725 25.775 262.075 27.025 ;
        RECT 265.425 25.455 265.765 26.285 ;
        RECT 267.245 25.775 267.595 27.025 ;
        RECT 270.945 25.455 271.285 26.285 ;
        RECT 272.765 25.775 273.115 27.025 ;
        RECT 274.880 26.370 277.470 27.460 ;
        RECT 274.880 25.680 276.090 26.200 ;
        RECT 276.260 25.850 277.470 26.370 ;
        RECT 278.100 26.295 278.390 27.460 ;
        RECT 278.560 27.025 283.905 27.460 ;
        RECT 284.080 27.025 289.425 27.460 ;
        RECT 289.600 27.025 294.945 27.460 ;
        RECT 295.120 27.025 300.465 27.460 ;
        RECT 252.800 24.910 258.145 25.455 ;
        RECT 258.320 24.910 263.665 25.455 ;
        RECT 263.840 24.910 269.185 25.455 ;
        RECT 269.360 24.910 274.705 25.455 ;
        RECT 274.880 24.910 277.470 25.680 ;
        RECT 278.100 24.910 278.390 25.635 ;
        RECT 280.145 25.455 280.485 26.285 ;
        RECT 281.965 25.775 282.315 27.025 ;
        RECT 285.665 25.455 286.005 26.285 ;
        RECT 287.485 25.775 287.835 27.025 ;
        RECT 291.185 25.455 291.525 26.285 ;
        RECT 293.005 25.775 293.355 27.025 ;
        RECT 296.705 25.455 297.045 26.285 ;
        RECT 298.525 25.775 298.875 27.025 ;
        RECT 300.640 26.370 303.230 27.460 ;
        RECT 300.640 25.680 301.850 26.200 ;
        RECT 302.020 25.850 303.230 26.370 ;
        RECT 303.860 26.295 304.150 27.460 ;
        RECT 304.320 27.025 309.665 27.460 ;
        RECT 278.560 24.910 283.905 25.455 ;
        RECT 284.080 24.910 289.425 25.455 ;
        RECT 289.600 24.910 294.945 25.455 ;
        RECT 295.120 24.910 300.465 25.455 ;
        RECT 300.640 24.910 303.230 25.680 ;
        RECT 303.860 24.910 304.150 25.635 ;
        RECT 305.905 25.455 306.245 26.285 ;
        RECT 307.725 25.775 308.075 27.025 ;
        RECT 309.840 26.370 311.050 27.460 ;
        RECT 309.840 25.830 310.360 26.370 ;
        RECT 310.530 25.660 311.050 26.200 ;
        RECT 304.320 24.910 309.665 25.455 ;
        RECT 309.840 24.910 311.050 25.660 ;
        RECT 162.095 24.740 311.135 24.910 ;
        RECT 162.180 23.990 163.390 24.740 ;
        RECT 163.560 24.195 168.905 24.740 ;
        RECT 169.080 24.195 174.425 24.740 ;
        RECT 174.600 24.195 179.945 24.740 ;
        RECT 180.120 24.195 185.465 24.740 ;
        RECT 162.180 23.450 162.700 23.990 ;
        RECT 162.870 23.280 163.390 23.820 ;
        RECT 165.145 23.365 165.485 24.195 ;
        RECT 162.180 22.190 163.390 23.280 ;
        RECT 166.965 22.625 167.315 23.875 ;
        RECT 170.665 23.365 171.005 24.195 ;
        RECT 172.485 22.625 172.835 23.875 ;
        RECT 176.185 23.365 176.525 24.195 ;
        RECT 178.005 22.625 178.355 23.875 ;
        RECT 181.705 23.365 182.045 24.195 ;
        RECT 185.640 23.970 187.310 24.740 ;
        RECT 187.940 24.015 188.230 24.740 ;
        RECT 188.400 24.195 193.745 24.740 ;
        RECT 193.920 24.195 199.265 24.740 ;
        RECT 199.440 24.195 204.785 24.740 ;
        RECT 204.960 24.195 210.305 24.740 ;
        RECT 183.525 22.625 183.875 23.875 ;
        RECT 185.640 23.450 186.390 23.970 ;
        RECT 186.560 23.280 187.310 23.800 ;
        RECT 189.985 23.365 190.325 24.195 ;
        RECT 163.560 22.190 168.905 22.625 ;
        RECT 169.080 22.190 174.425 22.625 ;
        RECT 174.600 22.190 179.945 22.625 ;
        RECT 180.120 22.190 185.465 22.625 ;
        RECT 185.640 22.190 187.310 23.280 ;
        RECT 187.940 22.190 188.230 23.355 ;
        RECT 191.805 22.625 192.155 23.875 ;
        RECT 195.505 23.365 195.845 24.195 ;
        RECT 197.325 22.625 197.675 23.875 ;
        RECT 201.025 23.365 201.365 24.195 ;
        RECT 202.845 22.625 203.195 23.875 ;
        RECT 206.545 23.365 206.885 24.195 ;
        RECT 210.480 23.970 213.070 24.740 ;
        RECT 213.700 24.015 213.990 24.740 ;
        RECT 214.160 24.195 219.505 24.740 ;
        RECT 219.680 24.195 225.025 24.740 ;
        RECT 225.200 24.195 230.545 24.740 ;
        RECT 230.720 24.195 236.065 24.740 ;
        RECT 208.365 22.625 208.715 23.875 ;
        RECT 210.480 23.450 211.690 23.970 ;
        RECT 211.860 23.280 213.070 23.800 ;
        RECT 215.745 23.365 216.085 24.195 ;
        RECT 188.400 22.190 193.745 22.625 ;
        RECT 193.920 22.190 199.265 22.625 ;
        RECT 199.440 22.190 204.785 22.625 ;
        RECT 204.960 22.190 210.305 22.625 ;
        RECT 210.480 22.190 213.070 23.280 ;
        RECT 213.700 22.190 213.990 23.355 ;
        RECT 217.565 22.625 217.915 23.875 ;
        RECT 221.265 23.365 221.605 24.195 ;
        RECT 223.085 22.625 223.435 23.875 ;
        RECT 226.785 23.365 227.125 24.195 ;
        RECT 228.605 22.625 228.955 23.875 ;
        RECT 232.305 23.365 232.645 24.195 ;
        RECT 236.240 23.970 238.830 24.740 ;
        RECT 239.460 24.015 239.750 24.740 ;
        RECT 239.920 24.195 245.265 24.740 ;
        RECT 245.440 24.195 250.785 24.740 ;
        RECT 250.960 24.195 256.305 24.740 ;
        RECT 256.480 24.195 261.825 24.740 ;
        RECT 234.125 22.625 234.475 23.875 ;
        RECT 236.240 23.450 237.450 23.970 ;
        RECT 237.620 23.280 238.830 23.800 ;
        RECT 241.505 23.365 241.845 24.195 ;
        RECT 214.160 22.190 219.505 22.625 ;
        RECT 219.680 22.190 225.025 22.625 ;
        RECT 225.200 22.190 230.545 22.625 ;
        RECT 230.720 22.190 236.065 22.625 ;
        RECT 236.240 22.190 238.830 23.280 ;
        RECT 239.460 22.190 239.750 23.355 ;
        RECT 243.325 22.625 243.675 23.875 ;
        RECT 247.025 23.365 247.365 24.195 ;
        RECT 248.845 22.625 249.195 23.875 ;
        RECT 252.545 23.365 252.885 24.195 ;
        RECT 254.365 22.625 254.715 23.875 ;
        RECT 258.065 23.365 258.405 24.195 ;
        RECT 262.000 23.970 264.590 24.740 ;
        RECT 265.220 24.015 265.510 24.740 ;
        RECT 265.680 24.195 271.025 24.740 ;
        RECT 271.200 24.195 276.545 24.740 ;
        RECT 276.720 24.195 282.065 24.740 ;
        RECT 282.240 24.195 287.585 24.740 ;
        RECT 259.885 22.625 260.235 23.875 ;
        RECT 262.000 23.450 263.210 23.970 ;
        RECT 263.380 23.280 264.590 23.800 ;
        RECT 267.265 23.365 267.605 24.195 ;
        RECT 239.920 22.190 245.265 22.625 ;
        RECT 245.440 22.190 250.785 22.625 ;
        RECT 250.960 22.190 256.305 22.625 ;
        RECT 256.480 22.190 261.825 22.625 ;
        RECT 262.000 22.190 264.590 23.280 ;
        RECT 265.220 22.190 265.510 23.355 ;
        RECT 269.085 22.625 269.435 23.875 ;
        RECT 272.785 23.365 273.125 24.195 ;
        RECT 274.605 22.625 274.955 23.875 ;
        RECT 278.305 23.365 278.645 24.195 ;
        RECT 280.125 22.625 280.475 23.875 ;
        RECT 283.825 23.365 284.165 24.195 ;
        RECT 287.760 23.970 290.350 24.740 ;
        RECT 290.980 24.015 291.270 24.740 ;
        RECT 291.440 24.195 296.785 24.740 ;
        RECT 296.960 24.195 302.305 24.740 ;
        RECT 302.480 24.195 307.825 24.740 ;
        RECT 285.645 22.625 285.995 23.875 ;
        RECT 287.760 23.450 288.970 23.970 ;
        RECT 289.140 23.280 290.350 23.800 ;
        RECT 293.025 23.365 293.365 24.195 ;
        RECT 265.680 22.190 271.025 22.625 ;
        RECT 271.200 22.190 276.545 22.625 ;
        RECT 276.720 22.190 282.065 22.625 ;
        RECT 282.240 22.190 287.585 22.625 ;
        RECT 287.760 22.190 290.350 23.280 ;
        RECT 290.980 22.190 291.270 23.355 ;
        RECT 294.845 22.625 295.195 23.875 ;
        RECT 298.545 23.365 298.885 24.195 ;
        RECT 300.365 22.625 300.715 23.875 ;
        RECT 304.065 23.365 304.405 24.195 ;
        RECT 308.000 23.970 309.670 24.740 ;
        RECT 309.840 23.990 311.050 24.740 ;
        RECT 305.885 22.625 306.235 23.875 ;
        RECT 308.000 23.450 308.750 23.970 ;
        RECT 308.920 23.280 309.670 23.800 ;
        RECT 291.440 22.190 296.785 22.625 ;
        RECT 296.960 22.190 302.305 22.625 ;
        RECT 302.480 22.190 307.825 22.625 ;
        RECT 308.000 22.190 309.670 23.280 ;
        RECT 309.840 23.280 310.360 23.820 ;
        RECT 310.530 23.450 311.050 23.990 ;
        RECT 309.840 22.190 311.050 23.280 ;
        RECT 162.095 22.020 311.135 22.190 ;
        RECT 162.180 20.930 163.390 22.020 ;
        RECT 163.560 21.585 168.905 22.020 ;
        RECT 169.080 21.585 174.425 22.020 ;
        RECT 162.180 20.220 162.700 20.760 ;
        RECT 162.870 20.390 163.390 20.930 ;
        RECT 162.180 19.470 163.390 20.220 ;
        RECT 165.145 20.015 165.485 20.845 ;
        RECT 166.965 20.335 167.315 21.585 ;
        RECT 170.665 20.015 171.005 20.845 ;
        RECT 172.485 20.335 172.835 21.585 ;
        RECT 175.060 20.855 175.350 22.020 ;
        RECT 175.520 21.585 180.865 22.020 ;
        RECT 181.040 21.585 186.385 22.020 ;
        RECT 186.560 21.585 191.905 22.020 ;
        RECT 192.080 21.585 197.425 22.020 ;
        RECT 163.560 19.470 168.905 20.015 ;
        RECT 169.080 19.470 174.425 20.015 ;
        RECT 175.060 19.470 175.350 20.195 ;
        RECT 177.105 20.015 177.445 20.845 ;
        RECT 178.925 20.335 179.275 21.585 ;
        RECT 182.625 20.015 182.965 20.845 ;
        RECT 184.445 20.335 184.795 21.585 ;
        RECT 188.145 20.015 188.485 20.845 ;
        RECT 189.965 20.335 190.315 21.585 ;
        RECT 193.665 20.015 194.005 20.845 ;
        RECT 195.485 20.335 195.835 21.585 ;
        RECT 197.600 20.930 200.190 22.020 ;
        RECT 197.600 20.240 198.810 20.760 ;
        RECT 198.980 20.410 200.190 20.930 ;
        RECT 200.820 20.855 201.110 22.020 ;
        RECT 201.280 21.585 206.625 22.020 ;
        RECT 206.800 21.585 212.145 22.020 ;
        RECT 212.320 21.585 217.665 22.020 ;
        RECT 217.840 21.585 223.185 22.020 ;
        RECT 175.520 19.470 180.865 20.015 ;
        RECT 181.040 19.470 186.385 20.015 ;
        RECT 186.560 19.470 191.905 20.015 ;
        RECT 192.080 19.470 197.425 20.015 ;
        RECT 197.600 19.470 200.190 20.240 ;
        RECT 200.820 19.470 201.110 20.195 ;
        RECT 202.865 20.015 203.205 20.845 ;
        RECT 204.685 20.335 205.035 21.585 ;
        RECT 208.385 20.015 208.725 20.845 ;
        RECT 210.205 20.335 210.555 21.585 ;
        RECT 213.905 20.015 214.245 20.845 ;
        RECT 215.725 20.335 216.075 21.585 ;
        RECT 219.425 20.015 219.765 20.845 ;
        RECT 221.245 20.335 221.595 21.585 ;
        RECT 223.360 20.930 225.950 22.020 ;
        RECT 223.360 20.240 224.570 20.760 ;
        RECT 224.740 20.410 225.950 20.930 ;
        RECT 226.580 20.855 226.870 22.020 ;
        RECT 227.040 21.585 232.385 22.020 ;
        RECT 232.560 21.585 237.905 22.020 ;
        RECT 238.080 21.585 243.425 22.020 ;
        RECT 243.600 21.585 248.945 22.020 ;
        RECT 201.280 19.470 206.625 20.015 ;
        RECT 206.800 19.470 212.145 20.015 ;
        RECT 212.320 19.470 217.665 20.015 ;
        RECT 217.840 19.470 223.185 20.015 ;
        RECT 223.360 19.470 225.950 20.240 ;
        RECT 226.580 19.470 226.870 20.195 ;
        RECT 228.625 20.015 228.965 20.845 ;
        RECT 230.445 20.335 230.795 21.585 ;
        RECT 234.145 20.015 234.485 20.845 ;
        RECT 235.965 20.335 236.315 21.585 ;
        RECT 239.665 20.015 240.005 20.845 ;
        RECT 241.485 20.335 241.835 21.585 ;
        RECT 245.185 20.015 245.525 20.845 ;
        RECT 247.005 20.335 247.355 21.585 ;
        RECT 249.120 20.930 251.710 22.020 ;
        RECT 249.120 20.240 250.330 20.760 ;
        RECT 250.500 20.410 251.710 20.930 ;
        RECT 252.340 20.855 252.630 22.020 ;
        RECT 252.800 21.585 258.145 22.020 ;
        RECT 258.320 21.585 263.665 22.020 ;
        RECT 263.840 21.585 269.185 22.020 ;
        RECT 269.360 21.585 274.705 22.020 ;
        RECT 227.040 19.470 232.385 20.015 ;
        RECT 232.560 19.470 237.905 20.015 ;
        RECT 238.080 19.470 243.425 20.015 ;
        RECT 243.600 19.470 248.945 20.015 ;
        RECT 249.120 19.470 251.710 20.240 ;
        RECT 252.340 19.470 252.630 20.195 ;
        RECT 254.385 20.015 254.725 20.845 ;
        RECT 256.205 20.335 256.555 21.585 ;
        RECT 259.905 20.015 260.245 20.845 ;
        RECT 261.725 20.335 262.075 21.585 ;
        RECT 265.425 20.015 265.765 20.845 ;
        RECT 267.245 20.335 267.595 21.585 ;
        RECT 270.945 20.015 271.285 20.845 ;
        RECT 272.765 20.335 273.115 21.585 ;
        RECT 274.880 20.930 277.470 22.020 ;
        RECT 274.880 20.240 276.090 20.760 ;
        RECT 276.260 20.410 277.470 20.930 ;
        RECT 278.100 20.855 278.390 22.020 ;
        RECT 278.560 21.585 283.905 22.020 ;
        RECT 284.080 21.585 289.425 22.020 ;
        RECT 289.600 21.585 294.945 22.020 ;
        RECT 295.120 21.585 300.465 22.020 ;
        RECT 252.800 19.470 258.145 20.015 ;
        RECT 258.320 19.470 263.665 20.015 ;
        RECT 263.840 19.470 269.185 20.015 ;
        RECT 269.360 19.470 274.705 20.015 ;
        RECT 274.880 19.470 277.470 20.240 ;
        RECT 278.100 19.470 278.390 20.195 ;
        RECT 280.145 20.015 280.485 20.845 ;
        RECT 281.965 20.335 282.315 21.585 ;
        RECT 285.665 20.015 286.005 20.845 ;
        RECT 287.485 20.335 287.835 21.585 ;
        RECT 291.185 20.015 291.525 20.845 ;
        RECT 293.005 20.335 293.355 21.585 ;
        RECT 296.705 20.015 297.045 20.845 ;
        RECT 298.525 20.335 298.875 21.585 ;
        RECT 300.640 20.930 303.230 22.020 ;
        RECT 300.640 20.240 301.850 20.760 ;
        RECT 302.020 20.410 303.230 20.930 ;
        RECT 303.860 20.855 304.150 22.020 ;
        RECT 304.320 21.585 309.665 22.020 ;
        RECT 278.560 19.470 283.905 20.015 ;
        RECT 284.080 19.470 289.425 20.015 ;
        RECT 289.600 19.470 294.945 20.015 ;
        RECT 295.120 19.470 300.465 20.015 ;
        RECT 300.640 19.470 303.230 20.240 ;
        RECT 303.860 19.470 304.150 20.195 ;
        RECT 305.905 20.015 306.245 20.845 ;
        RECT 307.725 20.335 308.075 21.585 ;
        RECT 309.840 20.930 311.050 22.020 ;
        RECT 309.840 20.390 310.360 20.930 ;
        RECT 310.530 20.220 311.050 20.760 ;
        RECT 304.320 19.470 309.665 20.015 ;
        RECT 309.840 19.470 311.050 20.220 ;
        RECT 162.095 19.300 311.135 19.470 ;
        RECT 162.180 18.550 163.390 19.300 ;
        RECT 163.560 18.755 168.905 19.300 ;
        RECT 169.080 18.755 174.425 19.300 ;
        RECT 174.600 18.755 179.945 19.300 ;
        RECT 180.120 18.755 185.465 19.300 ;
        RECT 162.180 18.010 162.700 18.550 ;
        RECT 162.870 17.840 163.390 18.380 ;
        RECT 165.145 17.925 165.485 18.755 ;
        RECT 162.180 16.750 163.390 17.840 ;
        RECT 166.965 17.185 167.315 18.435 ;
        RECT 170.665 17.925 171.005 18.755 ;
        RECT 172.485 17.185 172.835 18.435 ;
        RECT 176.185 17.925 176.525 18.755 ;
        RECT 178.005 17.185 178.355 18.435 ;
        RECT 181.705 17.925 182.045 18.755 ;
        RECT 185.640 18.530 187.310 19.300 ;
        RECT 187.940 18.575 188.230 19.300 ;
        RECT 188.400 18.755 193.745 19.300 ;
        RECT 193.920 18.755 199.265 19.300 ;
        RECT 199.440 18.755 204.785 19.300 ;
        RECT 204.960 18.755 210.305 19.300 ;
        RECT 183.525 17.185 183.875 18.435 ;
        RECT 185.640 18.010 186.390 18.530 ;
        RECT 186.560 17.840 187.310 18.360 ;
        RECT 189.985 17.925 190.325 18.755 ;
        RECT 163.560 16.750 168.905 17.185 ;
        RECT 169.080 16.750 174.425 17.185 ;
        RECT 174.600 16.750 179.945 17.185 ;
        RECT 180.120 16.750 185.465 17.185 ;
        RECT 185.640 16.750 187.310 17.840 ;
        RECT 187.940 16.750 188.230 17.915 ;
        RECT 191.805 17.185 192.155 18.435 ;
        RECT 195.505 17.925 195.845 18.755 ;
        RECT 197.325 17.185 197.675 18.435 ;
        RECT 201.025 17.925 201.365 18.755 ;
        RECT 202.845 17.185 203.195 18.435 ;
        RECT 206.545 17.925 206.885 18.755 ;
        RECT 210.480 18.530 213.070 19.300 ;
        RECT 213.700 18.575 213.990 19.300 ;
        RECT 214.160 18.755 219.505 19.300 ;
        RECT 219.680 18.755 225.025 19.300 ;
        RECT 225.200 18.755 230.545 19.300 ;
        RECT 230.720 18.755 236.065 19.300 ;
        RECT 208.365 17.185 208.715 18.435 ;
        RECT 210.480 18.010 211.690 18.530 ;
        RECT 211.860 17.840 213.070 18.360 ;
        RECT 215.745 17.925 216.085 18.755 ;
        RECT 188.400 16.750 193.745 17.185 ;
        RECT 193.920 16.750 199.265 17.185 ;
        RECT 199.440 16.750 204.785 17.185 ;
        RECT 204.960 16.750 210.305 17.185 ;
        RECT 210.480 16.750 213.070 17.840 ;
        RECT 213.700 16.750 213.990 17.915 ;
        RECT 217.565 17.185 217.915 18.435 ;
        RECT 221.265 17.925 221.605 18.755 ;
        RECT 223.085 17.185 223.435 18.435 ;
        RECT 226.785 17.925 227.125 18.755 ;
        RECT 228.605 17.185 228.955 18.435 ;
        RECT 232.305 17.925 232.645 18.755 ;
        RECT 236.240 18.530 238.830 19.300 ;
        RECT 239.460 18.575 239.750 19.300 ;
        RECT 239.920 18.755 245.265 19.300 ;
        RECT 245.440 18.755 250.785 19.300 ;
        RECT 250.960 18.755 256.305 19.300 ;
        RECT 256.480 18.755 261.825 19.300 ;
        RECT 234.125 17.185 234.475 18.435 ;
        RECT 236.240 18.010 237.450 18.530 ;
        RECT 237.620 17.840 238.830 18.360 ;
        RECT 241.505 17.925 241.845 18.755 ;
        RECT 214.160 16.750 219.505 17.185 ;
        RECT 219.680 16.750 225.025 17.185 ;
        RECT 225.200 16.750 230.545 17.185 ;
        RECT 230.720 16.750 236.065 17.185 ;
        RECT 236.240 16.750 238.830 17.840 ;
        RECT 239.460 16.750 239.750 17.915 ;
        RECT 243.325 17.185 243.675 18.435 ;
        RECT 247.025 17.925 247.365 18.755 ;
        RECT 248.845 17.185 249.195 18.435 ;
        RECT 252.545 17.925 252.885 18.755 ;
        RECT 254.365 17.185 254.715 18.435 ;
        RECT 258.065 17.925 258.405 18.755 ;
        RECT 262.000 18.530 264.590 19.300 ;
        RECT 265.220 18.575 265.510 19.300 ;
        RECT 265.680 18.755 271.025 19.300 ;
        RECT 271.200 18.755 276.545 19.300 ;
        RECT 276.720 18.755 282.065 19.300 ;
        RECT 282.240 18.755 287.585 19.300 ;
        RECT 259.885 17.185 260.235 18.435 ;
        RECT 262.000 18.010 263.210 18.530 ;
        RECT 263.380 17.840 264.590 18.360 ;
        RECT 267.265 17.925 267.605 18.755 ;
        RECT 239.920 16.750 245.265 17.185 ;
        RECT 245.440 16.750 250.785 17.185 ;
        RECT 250.960 16.750 256.305 17.185 ;
        RECT 256.480 16.750 261.825 17.185 ;
        RECT 262.000 16.750 264.590 17.840 ;
        RECT 265.220 16.750 265.510 17.915 ;
        RECT 269.085 17.185 269.435 18.435 ;
        RECT 272.785 17.925 273.125 18.755 ;
        RECT 274.605 17.185 274.955 18.435 ;
        RECT 278.305 17.925 278.645 18.755 ;
        RECT 280.125 17.185 280.475 18.435 ;
        RECT 283.825 17.925 284.165 18.755 ;
        RECT 287.760 18.530 290.350 19.300 ;
        RECT 290.980 18.575 291.270 19.300 ;
        RECT 291.440 18.755 296.785 19.300 ;
        RECT 296.960 18.755 302.305 19.300 ;
        RECT 302.480 18.755 307.825 19.300 ;
        RECT 285.645 17.185 285.995 18.435 ;
        RECT 287.760 18.010 288.970 18.530 ;
        RECT 289.140 17.840 290.350 18.360 ;
        RECT 293.025 17.925 293.365 18.755 ;
        RECT 265.680 16.750 271.025 17.185 ;
        RECT 271.200 16.750 276.545 17.185 ;
        RECT 276.720 16.750 282.065 17.185 ;
        RECT 282.240 16.750 287.585 17.185 ;
        RECT 287.760 16.750 290.350 17.840 ;
        RECT 290.980 16.750 291.270 17.915 ;
        RECT 294.845 17.185 295.195 18.435 ;
        RECT 298.545 17.925 298.885 18.755 ;
        RECT 300.365 17.185 300.715 18.435 ;
        RECT 304.065 17.925 304.405 18.755 ;
        RECT 308.000 18.530 309.670 19.300 ;
        RECT 309.840 18.550 311.050 19.300 ;
        RECT 305.885 17.185 306.235 18.435 ;
        RECT 308.000 18.010 308.750 18.530 ;
        RECT 308.920 17.840 309.670 18.360 ;
        RECT 291.440 16.750 296.785 17.185 ;
        RECT 296.960 16.750 302.305 17.185 ;
        RECT 302.480 16.750 307.825 17.185 ;
        RECT 308.000 16.750 309.670 17.840 ;
        RECT 309.840 17.840 310.360 18.380 ;
        RECT 310.530 18.010 311.050 18.550 ;
        RECT 309.840 16.750 311.050 17.840 ;
        RECT 162.095 16.580 311.135 16.750 ;
        RECT 162.180 15.490 163.390 16.580 ;
        RECT 163.560 16.145 168.905 16.580 ;
        RECT 169.080 16.145 174.425 16.580 ;
        RECT 162.180 14.780 162.700 15.320 ;
        RECT 162.870 14.950 163.390 15.490 ;
        RECT 162.180 14.030 163.390 14.780 ;
        RECT 165.145 14.575 165.485 15.405 ;
        RECT 166.965 14.895 167.315 16.145 ;
        RECT 170.665 14.575 171.005 15.405 ;
        RECT 172.485 14.895 172.835 16.145 ;
        RECT 175.060 15.415 175.350 16.580 ;
        RECT 175.520 16.145 180.865 16.580 ;
        RECT 181.040 16.145 186.385 16.580 ;
        RECT 163.560 14.030 168.905 14.575 ;
        RECT 169.080 14.030 174.425 14.575 ;
        RECT 175.060 14.030 175.350 14.755 ;
        RECT 177.105 14.575 177.445 15.405 ;
        RECT 178.925 14.895 179.275 16.145 ;
        RECT 182.625 14.575 182.965 15.405 ;
        RECT 184.445 14.895 184.795 16.145 ;
        RECT 186.560 15.490 187.770 16.580 ;
        RECT 186.560 14.780 187.080 15.320 ;
        RECT 187.250 14.950 187.770 15.490 ;
        RECT 187.940 15.415 188.230 16.580 ;
        RECT 188.400 16.145 193.745 16.580 ;
        RECT 193.920 16.145 199.265 16.580 ;
        RECT 175.520 14.030 180.865 14.575 ;
        RECT 181.040 14.030 186.385 14.575 ;
        RECT 186.560 14.030 187.770 14.780 ;
        RECT 187.940 14.030 188.230 14.755 ;
        RECT 189.985 14.575 190.325 15.405 ;
        RECT 191.805 14.895 192.155 16.145 ;
        RECT 195.505 14.575 195.845 15.405 ;
        RECT 197.325 14.895 197.675 16.145 ;
        RECT 199.440 15.490 200.650 16.580 ;
        RECT 199.440 14.780 199.960 15.320 ;
        RECT 200.130 14.950 200.650 15.490 ;
        RECT 200.820 15.415 201.110 16.580 ;
        RECT 201.280 16.145 206.625 16.580 ;
        RECT 206.800 16.145 212.145 16.580 ;
        RECT 188.400 14.030 193.745 14.575 ;
        RECT 193.920 14.030 199.265 14.575 ;
        RECT 199.440 14.030 200.650 14.780 ;
        RECT 200.820 14.030 201.110 14.755 ;
        RECT 202.865 14.575 203.205 15.405 ;
        RECT 204.685 14.895 205.035 16.145 ;
        RECT 208.385 14.575 208.725 15.405 ;
        RECT 210.205 14.895 210.555 16.145 ;
        RECT 212.320 15.490 213.530 16.580 ;
        RECT 212.320 14.780 212.840 15.320 ;
        RECT 213.010 14.950 213.530 15.490 ;
        RECT 213.700 15.415 213.990 16.580 ;
        RECT 214.160 16.145 219.505 16.580 ;
        RECT 219.680 16.145 225.025 16.580 ;
        RECT 201.280 14.030 206.625 14.575 ;
        RECT 206.800 14.030 212.145 14.575 ;
        RECT 212.320 14.030 213.530 14.780 ;
        RECT 213.700 14.030 213.990 14.755 ;
        RECT 215.745 14.575 216.085 15.405 ;
        RECT 217.565 14.895 217.915 16.145 ;
        RECT 221.265 14.575 221.605 15.405 ;
        RECT 223.085 14.895 223.435 16.145 ;
        RECT 225.200 15.490 226.410 16.580 ;
        RECT 225.200 14.780 225.720 15.320 ;
        RECT 225.890 14.950 226.410 15.490 ;
        RECT 226.580 15.415 226.870 16.580 ;
        RECT 227.040 16.145 232.385 16.580 ;
        RECT 232.560 16.145 237.905 16.580 ;
        RECT 214.160 14.030 219.505 14.575 ;
        RECT 219.680 14.030 225.025 14.575 ;
        RECT 225.200 14.030 226.410 14.780 ;
        RECT 226.580 14.030 226.870 14.755 ;
        RECT 228.625 14.575 228.965 15.405 ;
        RECT 230.445 14.895 230.795 16.145 ;
        RECT 234.145 14.575 234.485 15.405 ;
        RECT 235.965 14.895 236.315 16.145 ;
        RECT 238.080 15.490 239.290 16.580 ;
        RECT 238.080 14.780 238.600 15.320 ;
        RECT 238.770 14.950 239.290 15.490 ;
        RECT 239.460 15.415 239.750 16.580 ;
        RECT 239.920 16.145 245.265 16.580 ;
        RECT 245.440 16.145 250.785 16.580 ;
        RECT 227.040 14.030 232.385 14.575 ;
        RECT 232.560 14.030 237.905 14.575 ;
        RECT 238.080 14.030 239.290 14.780 ;
        RECT 239.460 14.030 239.750 14.755 ;
        RECT 241.505 14.575 241.845 15.405 ;
        RECT 243.325 14.895 243.675 16.145 ;
        RECT 247.025 14.575 247.365 15.405 ;
        RECT 248.845 14.895 249.195 16.145 ;
        RECT 250.960 15.490 252.170 16.580 ;
        RECT 250.960 14.780 251.480 15.320 ;
        RECT 251.650 14.950 252.170 15.490 ;
        RECT 252.340 15.415 252.630 16.580 ;
        RECT 252.800 16.145 258.145 16.580 ;
        RECT 258.320 16.145 263.665 16.580 ;
        RECT 239.920 14.030 245.265 14.575 ;
        RECT 245.440 14.030 250.785 14.575 ;
        RECT 250.960 14.030 252.170 14.780 ;
        RECT 252.340 14.030 252.630 14.755 ;
        RECT 254.385 14.575 254.725 15.405 ;
        RECT 256.205 14.895 256.555 16.145 ;
        RECT 259.905 14.575 260.245 15.405 ;
        RECT 261.725 14.895 262.075 16.145 ;
        RECT 263.840 15.490 265.050 16.580 ;
        RECT 263.840 14.780 264.360 15.320 ;
        RECT 264.530 14.950 265.050 15.490 ;
        RECT 265.220 15.415 265.510 16.580 ;
        RECT 265.680 16.145 271.025 16.580 ;
        RECT 271.200 16.145 276.545 16.580 ;
        RECT 252.800 14.030 258.145 14.575 ;
        RECT 258.320 14.030 263.665 14.575 ;
        RECT 263.840 14.030 265.050 14.780 ;
        RECT 265.220 14.030 265.510 14.755 ;
        RECT 267.265 14.575 267.605 15.405 ;
        RECT 269.085 14.895 269.435 16.145 ;
        RECT 272.785 14.575 273.125 15.405 ;
        RECT 274.605 14.895 274.955 16.145 ;
        RECT 276.720 15.490 277.930 16.580 ;
        RECT 276.720 14.780 277.240 15.320 ;
        RECT 277.410 14.950 277.930 15.490 ;
        RECT 278.100 15.415 278.390 16.580 ;
        RECT 278.560 16.145 283.905 16.580 ;
        RECT 284.080 16.145 289.425 16.580 ;
        RECT 265.680 14.030 271.025 14.575 ;
        RECT 271.200 14.030 276.545 14.575 ;
        RECT 276.720 14.030 277.930 14.780 ;
        RECT 278.100 14.030 278.390 14.755 ;
        RECT 280.145 14.575 280.485 15.405 ;
        RECT 281.965 14.895 282.315 16.145 ;
        RECT 285.665 14.575 286.005 15.405 ;
        RECT 287.485 14.895 287.835 16.145 ;
        RECT 289.600 15.490 290.810 16.580 ;
        RECT 289.600 14.780 290.120 15.320 ;
        RECT 290.290 14.950 290.810 15.490 ;
        RECT 290.980 15.415 291.270 16.580 ;
        RECT 291.440 16.145 296.785 16.580 ;
        RECT 296.960 16.145 302.305 16.580 ;
        RECT 278.560 14.030 283.905 14.575 ;
        RECT 284.080 14.030 289.425 14.575 ;
        RECT 289.600 14.030 290.810 14.780 ;
        RECT 290.980 14.030 291.270 14.755 ;
        RECT 293.025 14.575 293.365 15.405 ;
        RECT 294.845 14.895 295.195 16.145 ;
        RECT 298.545 14.575 298.885 15.405 ;
        RECT 300.365 14.895 300.715 16.145 ;
        RECT 302.480 15.490 303.690 16.580 ;
        RECT 302.480 14.780 303.000 15.320 ;
        RECT 303.170 14.950 303.690 15.490 ;
        RECT 303.860 15.415 304.150 16.580 ;
        RECT 304.320 16.145 309.665 16.580 ;
        RECT 291.440 14.030 296.785 14.575 ;
        RECT 296.960 14.030 302.305 14.575 ;
        RECT 302.480 14.030 303.690 14.780 ;
        RECT 303.860 14.030 304.150 14.755 ;
        RECT 305.905 14.575 306.245 15.405 ;
        RECT 307.725 14.895 308.075 16.145 ;
        RECT 309.840 15.490 311.050 16.580 ;
        RECT 309.840 14.950 310.360 15.490 ;
        RECT 310.530 14.780 311.050 15.320 ;
        RECT 304.320 14.030 309.665 14.575 ;
        RECT 309.840 14.030 311.050 14.780 ;
        RECT 162.095 13.860 311.135 14.030 ;
        RECT 4.300 4.300 155.700 4.700 ;
      LAYER met1 ;
        RECT 45.390 225.410 246.965 225.710 ;
        RECT 45.390 224.810 45.690 225.410 ;
        RECT 59.190 224.810 233.315 225.110 ;
        RECT 246.665 225.010 246.965 225.410 ;
        RECT 62.000 224.210 223.655 224.510 ;
        RECT 233.015 224.410 233.315 224.810 ;
        RECT 223.355 223.810 223.655 224.210 ;
        RECT 4.100 216.515 102.825 222.630 ;
        RECT 106.340 220.315 153.245 220.715 ;
        RECT 106.340 217.515 108.920 220.315 ;
        RECT 109.605 219.705 110.565 219.935 ;
        RECT 110.895 219.705 111.855 220.055 ;
        RECT 109.325 219.255 109.555 219.500 ;
        RECT 110.615 219.255 110.845 219.500 ;
        RECT 111.905 219.255 112.135 219.500 ;
        RECT 109.290 217.755 109.590 219.255 ;
        RECT 110.580 217.755 110.880 219.255 ;
        RECT 111.870 217.755 112.170 219.255 ;
        RECT 4.100 212.490 63.455 216.515 ;
        RECT 64.175 215.825 80.135 216.055 ;
        RECT 81.805 215.825 97.765 216.055 ;
        RECT 63.895 214.620 64.125 215.620 ;
        RECT 80.185 214.620 81.755 215.620 ;
        RECT 97.815 214.620 98.045 215.620 ;
        RECT 64.175 214.185 80.135 214.415 ;
        RECT 81.805 214.185 97.765 214.415 ;
        RECT 77.595 213.035 78.595 213.270 ;
        RECT 83.345 213.035 84.345 213.270 ;
        RECT 64.175 212.805 80.135 213.035 ;
        RECT 81.805 212.805 97.765 213.035 ;
        RECT 4.100 211.660 56.570 212.490 ;
        RECT 4.100 191.850 9.525 211.660 ;
        RECT 10.245 210.970 18.205 211.200 ;
        RECT 18.535 210.970 26.495 211.200 ;
        RECT 28.165 210.970 36.125 211.200 ;
        RECT 36.455 210.970 44.415 211.200 ;
        RECT 9.965 210.465 10.195 210.765 ;
        RECT 9.925 209.065 10.225 210.465 ;
        RECT 9.965 202.765 10.195 209.065 ;
        RECT 18.255 207.465 18.485 210.765 ;
        RECT 18.215 206.065 18.515 207.465 ;
        RECT 18.255 202.765 18.485 206.065 ;
        RECT 26.545 204.465 26.775 210.765 ;
        RECT 27.885 204.465 28.115 210.765 ;
        RECT 36.175 207.465 36.405 210.765 ;
        RECT 44.465 210.465 44.695 210.765 ;
        RECT 44.425 209.065 44.725 210.465 ;
        RECT 45.135 210.150 56.570 211.660 ;
        RECT 36.165 206.065 36.465 207.465 ;
        RECT 26.505 203.065 26.805 204.465 ;
        RECT 27.845 203.065 28.145 204.465 ;
        RECT 26.505 202.560 28.145 203.065 ;
        RECT 36.175 202.765 36.405 206.065 ;
        RECT 44.465 202.765 44.695 209.065 ;
        RECT 45.135 207.460 50.745 210.150 ;
        RECT 54.835 209.565 56.570 210.150 ;
        RECT 51.315 207.460 51.905 209.565 ;
        RECT 52.485 207.460 54.245 209.565 ;
        RECT 54.825 207.460 56.570 209.565 ;
        RECT 10.245 202.330 18.205 202.560 ;
        RECT 18.535 202.330 36.125 202.560 ;
        RECT 36.455 202.330 44.415 202.560 ;
        RECT 10.245 201.180 44.415 202.330 ;
        RECT 10.245 200.950 18.205 201.180 ;
        RECT 18.535 200.950 36.125 201.180 ;
        RECT 36.455 200.950 44.415 201.180 ;
        RECT 9.965 194.445 10.195 200.745 ;
        RECT 18.255 197.445 18.485 200.745 ;
        RECT 26.505 200.445 28.145 200.950 ;
        RECT 26.505 199.045 26.805 200.445 ;
        RECT 27.845 199.045 28.145 200.445 ;
        RECT 18.215 196.045 18.515 197.445 ;
        RECT 9.925 193.045 10.225 194.445 ;
        RECT 9.965 192.745 10.195 193.045 ;
        RECT 18.255 192.745 18.485 196.045 ;
        RECT 26.545 192.745 26.775 199.045 ;
        RECT 27.885 192.745 28.115 199.045 ;
        RECT 36.175 197.445 36.405 200.745 ;
        RECT 36.165 196.045 36.465 197.445 ;
        RECT 36.175 192.745 36.405 196.045 ;
        RECT 44.465 194.445 44.695 200.745 ;
        RECT 44.425 193.045 44.725 194.445 ;
        RECT 44.465 192.745 44.695 193.045 ;
        RECT 10.245 192.310 18.205 192.540 ;
        RECT 18.535 192.310 26.495 192.540 ;
        RECT 28.165 192.310 36.125 192.540 ;
        RECT 36.455 192.310 44.415 192.540 ;
        RECT 45.135 191.850 49.450 207.460 ;
        RECT 4.100 190.670 49.450 191.850 ;
        RECT 4.100 180.880 9.525 190.670 ;
        RECT 9.965 189.980 12.205 190.210 ;
        RECT 12.535 189.980 14.495 190.210 ;
        RECT 9.965 184.050 10.195 189.980 ;
        RECT 12.535 189.775 13.090 189.980 ;
        RECT 12.255 189.350 13.090 189.775 ;
        RECT 9.930 182.650 10.230 184.050 ;
        RECT 9.965 181.570 10.195 182.650 ;
        RECT 12.255 181.775 12.485 189.350 ;
        RECT 14.545 188.900 14.775 189.775 ;
        RECT 14.510 187.500 14.810 188.900 ;
        RECT 14.545 181.775 14.775 187.500 ;
        RECT 9.965 181.340 12.205 181.570 ;
        RECT 12.535 181.340 14.495 181.570 ;
        RECT 15.215 180.880 16.545 190.670 ;
        RECT 45.135 190.570 49.450 190.670 ;
        RECT 56.110 190.570 56.570 207.460 ;
        RECT 17.265 189.980 19.225 190.210 ;
        RECT 19.555 189.980 21.515 190.210 ;
        RECT 21.845 189.980 23.805 190.210 ;
        RECT 24.135 189.980 26.095 190.210 ;
        RECT 26.425 189.980 28.385 190.210 ;
        RECT 28.715 189.980 30.675 190.210 ;
        RECT 31.005 189.980 32.965 190.210 ;
        RECT 33.295 189.980 35.255 190.210 ;
        RECT 35.585 189.980 37.545 190.210 ;
        RECT 37.875 189.980 39.835 190.210 ;
        RECT 40.165 189.980 42.125 190.210 ;
        RECT 42.455 189.980 44.415 190.210 ;
        RECT 16.985 189.645 17.215 189.775 ;
        RECT 16.950 188.245 17.250 189.645 ;
        RECT 16.985 181.775 17.215 188.245 ;
        RECT 19.275 186.555 19.505 189.775 ;
        RECT 21.565 189.645 21.795 189.775 ;
        RECT 21.530 188.245 21.830 189.645 ;
        RECT 19.240 184.995 19.540 186.555 ;
        RECT 19.275 181.775 19.505 184.995 ;
        RECT 21.565 181.775 21.795 188.245 ;
        RECT 23.855 186.555 24.085 189.775 ;
        RECT 26.145 189.645 26.375 189.775 ;
        RECT 26.110 188.245 26.410 189.645 ;
        RECT 23.820 184.995 24.120 186.555 ;
        RECT 23.855 181.775 24.085 184.995 ;
        RECT 26.145 181.775 26.375 188.245 ;
        RECT 28.435 186.555 28.665 189.775 ;
        RECT 30.725 189.645 30.955 189.775 ;
        RECT 30.690 188.245 30.990 189.645 ;
        RECT 28.400 184.995 28.700 186.555 ;
        RECT 28.435 181.775 28.665 184.995 ;
        RECT 30.725 181.775 30.955 188.245 ;
        RECT 33.015 186.555 33.245 189.775 ;
        RECT 35.305 189.645 35.535 189.775 ;
        RECT 35.270 188.245 35.570 189.645 ;
        RECT 32.980 184.995 33.280 186.555 ;
        RECT 33.015 181.775 33.245 184.995 ;
        RECT 35.305 181.775 35.535 188.245 ;
        RECT 37.595 186.555 37.825 189.775 ;
        RECT 39.885 189.645 40.115 189.775 ;
        RECT 39.850 188.245 40.150 189.645 ;
        RECT 37.560 184.995 37.860 186.555 ;
        RECT 37.595 181.775 37.825 184.995 ;
        RECT 39.885 181.775 40.115 188.245 ;
        RECT 42.175 186.555 42.405 189.775 ;
        RECT 44.465 189.645 44.695 189.775 ;
        RECT 44.430 188.245 44.730 189.645 ;
        RECT 42.140 184.995 42.440 186.555 ;
        RECT 42.175 181.775 42.405 184.995 ;
        RECT 44.465 181.775 44.695 188.245 ;
        RECT 45.135 187.880 50.745 190.570 ;
        RECT 51.315 188.465 53.075 190.570 ;
        RECT 53.655 188.465 54.245 190.570 ;
        RECT 54.825 188.465 56.570 190.570 ;
        RECT 54.835 187.880 56.570 188.465 ;
        RECT 45.135 187.650 56.570 187.880 ;
        RECT 17.465 181.570 19.025 181.605 ;
        RECT 19.755 181.570 21.315 181.605 ;
        RECT 22.045 181.570 23.605 181.605 ;
        RECT 24.335 181.570 25.895 181.605 ;
        RECT 26.625 181.570 28.185 181.605 ;
        RECT 28.915 181.570 30.475 181.605 ;
        RECT 31.205 181.570 32.765 181.605 ;
        RECT 33.495 181.570 35.055 181.605 ;
        RECT 35.785 181.570 37.345 181.605 ;
        RECT 38.075 181.570 39.635 181.605 ;
        RECT 40.365 181.570 41.925 181.605 ;
        RECT 42.655 181.570 44.215 181.605 ;
        RECT 17.265 181.340 44.415 181.570 ;
        RECT 17.465 181.305 19.025 181.340 ;
        RECT 19.755 181.305 21.315 181.340 ;
        RECT 22.045 181.305 23.605 181.340 ;
        RECT 24.335 181.305 25.895 181.340 ;
        RECT 26.625 181.305 28.185 181.340 ;
        RECT 28.915 181.305 30.475 181.340 ;
        RECT 31.205 181.305 32.765 181.340 ;
        RECT 33.495 181.305 35.055 181.340 ;
        RECT 35.785 181.305 37.345 181.340 ;
        RECT 38.075 181.305 39.635 181.340 ;
        RECT 40.365 181.305 41.925 181.340 ;
        RECT 42.655 181.305 44.215 181.340 ;
        RECT 45.135 180.880 46.085 187.650 ;
        RECT 4.100 180.050 46.085 180.880 ;
        RECT 4.100 127.485 4.900 180.050 ;
        RECT 5.910 178.420 53.180 179.250 ;
        RECT 5.910 168.720 9.530 178.420 ;
        RECT 17.400 177.960 18.800 178.130 ;
        RECT 19.690 177.960 21.090 178.130 ;
        RECT 26.560 177.960 27.960 178.130 ;
        RECT 28.850 177.960 30.250 178.130 ;
        RECT 35.720 177.960 37.120 178.130 ;
        RECT 38.010 177.960 39.410 178.130 ;
        RECT 44.880 177.960 46.280 178.130 ;
        RECT 47.170 177.960 48.570 178.130 ;
        RECT 49.460 177.960 50.860 178.130 ;
        RECT 10.250 177.730 12.210 177.960 ;
        RECT 12.540 177.730 14.500 177.960 ;
        RECT 14.830 177.730 16.790 177.960 ;
        RECT 17.120 177.730 19.080 177.960 ;
        RECT 19.410 177.730 21.370 177.960 ;
        RECT 21.700 177.730 23.660 177.960 ;
        RECT 23.990 177.730 25.950 177.960 ;
        RECT 26.280 177.730 28.240 177.960 ;
        RECT 28.570 177.730 30.530 177.960 ;
        RECT 30.860 177.730 32.820 177.960 ;
        RECT 33.150 177.730 35.110 177.960 ;
        RECT 35.440 177.730 37.400 177.960 ;
        RECT 37.730 177.730 39.690 177.960 ;
        RECT 40.020 177.730 41.980 177.960 ;
        RECT 42.310 177.730 44.270 177.960 ;
        RECT 44.600 177.730 46.560 177.960 ;
        RECT 46.890 177.730 48.850 177.960 ;
        RECT 49.180 177.730 51.140 177.960 ;
        RECT 9.970 174.270 10.200 177.570 ;
        RECT 12.260 174.270 12.490 177.570 ;
        RECT 14.550 176.670 14.780 177.570 ;
        RECT 14.465 175.270 14.865 176.670 ;
        RECT 9.885 172.870 10.285 174.270 ;
        RECT 12.175 172.870 12.575 174.270 ;
        RECT 9.970 169.570 10.200 172.870 ;
        RECT 12.260 169.570 12.490 172.870 ;
        RECT 14.550 169.570 14.780 175.270 ;
        RECT 16.840 174.270 17.070 177.570 ;
        RECT 16.755 172.870 17.155 174.270 ;
        RECT 16.840 169.570 17.070 172.870 ;
        RECT 19.130 171.870 19.360 177.570 ;
        RECT 21.420 174.270 21.650 177.570 ;
        RECT 23.710 176.670 23.940 177.570 ;
        RECT 23.625 175.270 24.025 176.670 ;
        RECT 21.335 172.870 21.735 174.270 ;
        RECT 19.045 170.470 19.445 171.870 ;
        RECT 19.130 169.570 19.360 170.470 ;
        RECT 21.420 169.570 21.650 172.870 ;
        RECT 23.710 169.570 23.940 175.270 ;
        RECT 26.000 174.270 26.230 177.570 ;
        RECT 25.915 172.870 26.315 174.270 ;
        RECT 26.000 169.570 26.230 172.870 ;
        RECT 28.290 171.870 28.520 177.570 ;
        RECT 30.580 174.270 30.810 177.570 ;
        RECT 32.870 176.670 33.100 177.570 ;
        RECT 32.785 175.270 33.185 176.670 ;
        RECT 30.495 172.870 30.895 174.270 ;
        RECT 28.205 170.470 28.605 171.870 ;
        RECT 28.290 169.570 28.520 170.470 ;
        RECT 30.580 169.570 30.810 172.870 ;
        RECT 32.870 169.570 33.100 175.270 ;
        RECT 35.160 174.270 35.390 177.570 ;
        RECT 35.075 172.870 35.475 174.270 ;
        RECT 35.160 169.570 35.390 172.870 ;
        RECT 37.450 171.870 37.680 177.570 ;
        RECT 39.740 174.270 39.970 177.570 ;
        RECT 42.030 176.670 42.260 177.570 ;
        RECT 41.945 175.270 42.345 176.670 ;
        RECT 39.655 172.870 40.055 174.270 ;
        RECT 37.365 170.470 37.765 171.870 ;
        RECT 37.450 169.570 37.680 170.470 ;
        RECT 39.740 169.570 39.970 172.870 ;
        RECT 42.030 169.570 42.260 175.270 ;
        RECT 44.320 174.270 44.550 177.570 ;
        RECT 44.235 172.870 44.635 174.270 ;
        RECT 44.320 169.570 44.550 172.870 ;
        RECT 46.610 171.870 46.840 177.570 ;
        RECT 48.900 174.270 49.130 177.570 ;
        RECT 51.190 174.270 51.420 177.570 ;
        RECT 48.815 172.870 49.215 174.270 ;
        RECT 51.105 172.870 51.505 174.270 ;
        RECT 46.525 170.470 46.925 171.870 ;
        RECT 46.610 169.570 46.840 170.470 ;
        RECT 48.900 169.570 49.130 172.870 ;
        RECT 51.190 169.570 51.420 172.870 ;
        RECT 10.250 169.180 12.210 169.410 ;
        RECT 12.540 169.180 14.500 169.410 ;
        RECT 14.830 169.180 16.790 169.410 ;
        RECT 17.120 169.180 19.080 169.410 ;
        RECT 19.410 169.180 21.370 169.410 ;
        RECT 21.700 169.180 23.660 169.410 ;
        RECT 23.990 169.180 25.950 169.410 ;
        RECT 26.280 169.180 28.240 169.410 ;
        RECT 28.570 169.180 30.530 169.410 ;
        RECT 30.860 169.180 32.820 169.410 ;
        RECT 33.150 169.180 35.110 169.410 ;
        RECT 35.440 169.180 37.400 169.410 ;
        RECT 37.730 169.180 39.690 169.410 ;
        RECT 40.020 169.180 41.980 169.410 ;
        RECT 42.310 169.180 44.270 169.410 ;
        RECT 44.600 169.180 46.560 169.410 ;
        RECT 46.890 169.180 48.850 169.410 ;
        RECT 49.180 169.180 51.140 169.410 ;
        RECT 10.530 169.010 11.930 169.180 ;
        RECT 12.820 169.010 14.220 169.180 ;
        RECT 15.110 169.010 16.510 169.180 ;
        RECT 21.980 169.010 23.380 169.180 ;
        RECT 24.270 169.010 25.670 169.180 ;
        RECT 31.140 169.010 32.540 169.180 ;
        RECT 33.430 169.010 34.830 169.180 ;
        RECT 40.300 169.010 41.700 169.180 ;
        RECT 42.590 169.010 43.990 169.180 ;
        RECT 51.860 168.720 53.180 178.420 ;
        RECT 5.910 167.830 53.180 168.720 ;
        RECT 5.910 148.290 9.530 167.830 ;
        RECT 10.310 167.140 12.270 167.370 ;
        RECT 12.600 167.140 14.560 167.370 ;
        RECT 16.350 167.140 18.310 167.370 ;
        RECT 18.640 167.140 20.600 167.370 ;
        RECT 22.390 167.140 24.350 167.370 ;
        RECT 24.680 167.140 26.640 167.370 ;
        RECT 28.430 167.140 30.390 167.370 ;
        RECT 30.720 167.140 32.680 167.370 ;
        RECT 34.470 167.140 36.430 167.370 ;
        RECT 36.760 167.140 38.720 167.370 ;
        RECT 40.510 167.140 42.470 167.370 ;
        RECT 42.800 167.140 44.760 167.370 ;
        RECT 46.550 167.140 48.510 167.370 ;
        RECT 48.840 167.140 50.800 167.370 ;
        RECT 10.030 161.265 10.260 166.980 ;
        RECT 12.320 161.265 12.550 166.980 ;
        RECT 14.610 161.265 14.840 166.980 ;
        RECT 16.070 161.265 16.300 166.980 ;
        RECT 18.360 166.565 18.590 166.980 ;
        RECT 18.325 165.865 18.625 166.565 ;
        RECT 9.995 159.865 10.295 161.265 ;
        RECT 12.285 159.865 12.585 161.265 ;
        RECT 14.575 159.865 14.875 161.265 ;
        RECT 16.035 159.865 16.335 161.265 ;
        RECT 10.030 158.820 10.260 159.865 ;
        RECT 12.320 158.820 12.550 159.865 ;
        RECT 14.610 158.820 14.840 159.865 ;
        RECT 16.070 158.980 16.300 159.865 ;
        RECT 18.360 158.980 18.590 165.865 ;
        RECT 20.650 161.265 20.880 166.980 ;
        RECT 22.110 161.265 22.340 166.980 ;
        RECT 24.400 166.565 24.630 166.980 ;
        RECT 24.365 165.865 24.665 166.565 ;
        RECT 20.615 159.865 20.915 161.265 ;
        RECT 22.075 159.865 22.375 161.265 ;
        RECT 20.650 158.980 20.880 159.865 ;
        RECT 22.110 158.980 22.340 159.865 ;
        RECT 24.400 158.980 24.630 165.865 ;
        RECT 26.690 161.265 26.920 166.980 ;
        RECT 28.150 161.265 28.380 166.980 ;
        RECT 30.440 162.965 30.670 166.980 ;
        RECT 30.405 162.265 30.705 162.965 ;
        RECT 26.655 159.865 26.955 161.265 ;
        RECT 28.115 159.865 28.415 161.265 ;
        RECT 26.690 158.980 26.920 159.865 ;
        RECT 28.150 158.980 28.380 159.865 ;
        RECT 30.440 158.980 30.670 162.265 ;
        RECT 32.730 161.265 32.960 166.980 ;
        RECT 34.190 161.265 34.420 166.980 ;
        RECT 36.480 166.565 36.710 166.980 ;
        RECT 36.445 165.865 36.745 166.565 ;
        RECT 32.695 159.865 32.995 161.265 ;
        RECT 34.155 159.865 34.455 161.265 ;
        RECT 32.730 158.980 32.960 159.865 ;
        RECT 34.190 158.980 34.420 159.865 ;
        RECT 36.480 158.980 36.710 165.865 ;
        RECT 38.770 161.265 39.000 166.980 ;
        RECT 40.230 161.265 40.460 166.980 ;
        RECT 42.520 166.565 42.750 166.980 ;
        RECT 42.485 165.865 42.785 166.565 ;
        RECT 38.735 159.865 39.035 161.265 ;
        RECT 40.195 159.865 40.495 161.265 ;
        RECT 38.770 158.980 39.000 159.865 ;
        RECT 40.230 158.980 40.460 159.865 ;
        RECT 42.520 158.980 42.750 165.865 ;
        RECT 44.810 161.265 45.040 166.980 ;
        RECT 46.270 161.265 46.500 166.980 ;
        RECT 48.560 161.265 48.790 166.980 ;
        RECT 50.850 161.265 51.080 166.980 ;
        RECT 44.775 159.865 45.075 161.265 ;
        RECT 46.235 159.865 46.535 161.265 ;
        RECT 48.525 159.865 48.825 161.265 ;
        RECT 50.815 159.865 51.115 161.265 ;
        RECT 44.810 158.980 45.040 159.865 ;
        RECT 46.270 158.820 46.500 159.865 ;
        RECT 48.560 158.820 48.790 159.865 ;
        RECT 50.850 158.820 51.080 159.865 ;
        RECT 10.030 158.590 14.840 158.820 ;
        RECT 10.030 157.210 14.840 157.440 ;
        RECT 16.350 157.210 44.760 158.820 ;
        RECT 46.270 158.590 51.080 158.820 ;
        RECT 46.270 157.210 51.080 157.440 ;
        RECT 10.030 156.165 10.260 157.210 ;
        RECT 12.320 156.165 12.550 157.210 ;
        RECT 14.610 156.165 14.840 157.210 ;
        RECT 16.070 156.165 16.300 157.050 ;
        RECT 9.995 154.765 10.295 156.165 ;
        RECT 12.285 154.765 12.585 156.165 ;
        RECT 14.575 154.765 14.875 156.165 ;
        RECT 16.035 154.765 16.335 156.165 ;
        RECT 10.030 149.050 10.260 154.765 ;
        RECT 12.320 149.050 12.550 154.765 ;
        RECT 14.610 149.050 14.840 154.765 ;
        RECT 16.070 149.050 16.300 154.765 ;
        RECT 18.360 150.165 18.590 157.050 ;
        RECT 20.650 156.165 20.880 157.050 ;
        RECT 22.110 156.165 22.340 157.050 ;
        RECT 20.615 154.765 20.915 156.165 ;
        RECT 22.075 154.765 22.375 156.165 ;
        RECT 18.325 149.465 18.625 150.165 ;
        RECT 18.360 149.050 18.590 149.465 ;
        RECT 20.650 149.050 20.880 154.765 ;
        RECT 22.110 149.050 22.340 154.765 ;
        RECT 24.400 151.965 24.630 157.050 ;
        RECT 26.690 156.165 26.920 157.050 ;
        RECT 28.150 156.165 28.380 157.050 ;
        RECT 26.655 154.765 26.955 156.165 ;
        RECT 28.115 154.765 28.415 156.165 ;
        RECT 24.365 151.265 24.665 151.965 ;
        RECT 24.400 149.050 24.630 151.265 ;
        RECT 26.690 149.050 26.920 154.765 ;
        RECT 28.150 149.050 28.380 154.765 ;
        RECT 30.440 149.050 30.670 157.210 ;
        RECT 32.730 156.165 32.960 157.050 ;
        RECT 32.695 154.765 32.995 156.165 ;
        RECT 32.730 149.050 32.960 154.765 ;
        RECT 34.190 149.050 34.420 157.210 ;
        RECT 36.480 149.050 36.710 157.210 ;
        RECT 38.770 149.050 39.000 157.210 ;
        RECT 40.230 156.165 40.460 157.050 ;
        RECT 40.195 154.765 40.495 156.165 ;
        RECT 40.230 149.050 40.460 154.765 ;
        RECT 42.520 150.165 42.750 157.050 ;
        RECT 44.810 156.165 45.040 157.050 ;
        RECT 46.270 156.165 46.500 157.210 ;
        RECT 48.560 156.165 48.790 157.210 ;
        RECT 50.850 156.165 51.080 157.210 ;
        RECT 44.775 154.765 45.075 156.165 ;
        RECT 46.235 154.765 46.535 156.165 ;
        RECT 48.525 154.765 48.825 156.165 ;
        RECT 50.815 154.765 51.115 156.165 ;
        RECT 42.485 149.465 42.785 150.165 ;
        RECT 42.520 149.050 42.750 149.465 ;
        RECT 44.810 149.050 45.040 154.765 ;
        RECT 46.270 149.050 46.500 154.765 ;
        RECT 48.560 149.050 48.790 154.765 ;
        RECT 50.850 149.050 51.080 154.765 ;
        RECT 10.310 148.660 12.270 148.890 ;
        RECT 12.600 148.660 14.560 148.890 ;
        RECT 16.350 148.660 18.310 148.890 ;
        RECT 18.640 148.660 20.600 148.890 ;
        RECT 22.390 148.660 24.350 148.890 ;
        RECT 24.680 148.660 26.640 148.890 ;
        RECT 28.430 148.660 30.390 148.890 ;
        RECT 30.720 148.660 32.680 148.890 ;
        RECT 34.470 148.660 36.430 148.890 ;
        RECT 36.760 148.660 38.720 148.890 ;
        RECT 40.510 148.660 42.470 148.890 ;
        RECT 42.800 148.660 44.760 148.890 ;
        RECT 46.550 148.660 48.510 148.890 ;
        RECT 48.840 148.660 50.800 148.890 ;
        RECT 51.580 148.290 53.180 167.830 ;
        RECT 5.910 143.745 53.180 148.290 ;
        RECT 62.865 171.445 63.455 212.490 ;
        RECT 63.895 211.600 64.595 212.600 ;
        RECT 77.595 212.570 78.595 212.805 ;
        RECT 77.595 211.395 78.595 211.630 ;
        RECT 80.185 211.600 81.755 212.600 ;
        RECT 83.345 212.570 84.345 212.805 ;
        RECT 83.345 211.395 84.345 211.630 ;
        RECT 97.345 211.600 98.045 212.600 ;
        RECT 64.175 211.165 80.135 211.395 ;
        RECT 81.805 211.165 97.765 211.395 ;
        RECT 77.595 210.930 78.595 211.165 ;
        RECT 83.345 210.930 84.345 211.165 ;
        RECT 77.595 210.015 78.595 210.250 ;
        RECT 83.345 210.015 84.345 210.250 ;
        RECT 64.175 209.785 80.135 210.015 ;
        RECT 81.805 209.785 97.765 210.015 ;
        RECT 63.895 208.580 64.595 209.580 ;
        RECT 77.595 209.550 78.595 209.785 ;
        RECT 77.595 208.375 78.595 208.610 ;
        RECT 80.185 208.580 81.755 209.580 ;
        RECT 83.345 209.550 84.345 209.785 ;
        RECT 83.345 208.375 84.345 208.610 ;
        RECT 97.345 208.580 98.045 209.580 ;
        RECT 64.175 208.145 80.135 208.375 ;
        RECT 81.805 208.145 97.765 208.375 ;
        RECT 77.595 207.910 78.595 208.145 ;
        RECT 83.345 207.910 84.345 208.145 ;
        RECT 77.595 206.995 78.595 207.230 ;
        RECT 83.345 206.995 84.345 207.230 ;
        RECT 64.175 206.765 80.135 206.995 ;
        RECT 81.805 206.765 97.765 206.995 ;
        RECT 63.895 205.560 64.595 206.560 ;
        RECT 77.595 206.530 78.595 206.765 ;
        RECT 77.595 205.355 78.595 205.590 ;
        RECT 80.185 205.560 81.755 206.560 ;
        RECT 83.345 206.530 84.345 206.765 ;
        RECT 83.345 205.355 84.345 205.590 ;
        RECT 97.345 205.560 98.045 206.560 ;
        RECT 64.175 205.125 80.135 205.355 ;
        RECT 81.805 205.125 97.765 205.355 ;
        RECT 77.595 204.890 78.595 205.125 ;
        RECT 83.345 204.890 84.345 205.125 ;
        RECT 77.595 203.975 78.595 204.210 ;
        RECT 83.345 203.975 84.345 204.210 ;
        RECT 64.175 203.745 80.135 203.975 ;
        RECT 81.805 203.745 97.765 203.975 ;
        RECT 63.895 202.540 75.695 203.540 ;
        RECT 77.595 203.510 78.595 203.745 ;
        RECT 77.595 202.335 78.595 202.570 ;
        RECT 80.185 202.540 81.755 203.540 ;
        RECT 83.345 203.510 84.345 203.745 ;
        RECT 83.345 202.335 84.345 202.570 ;
        RECT 86.245 202.540 98.045 203.540 ;
        RECT 64.175 202.105 80.135 202.335 ;
        RECT 81.805 202.105 97.765 202.335 ;
        RECT 77.595 201.870 78.595 202.105 ;
        RECT 83.345 201.870 84.345 202.105 ;
        RECT 77.595 200.955 78.595 201.190 ;
        RECT 83.345 200.955 84.345 201.190 ;
        RECT 64.175 200.725 80.135 200.955 ;
        RECT 81.805 200.725 97.765 200.955 ;
        RECT 63.895 199.520 70.195 200.520 ;
        RECT 77.595 200.490 78.595 200.725 ;
        RECT 77.595 199.315 78.595 199.550 ;
        RECT 80.185 199.520 81.755 200.520 ;
        RECT 83.345 200.490 84.345 200.725 ;
        RECT 83.345 199.315 84.345 199.550 ;
        RECT 91.745 199.520 98.045 200.520 ;
        RECT 64.175 199.085 80.135 199.315 ;
        RECT 81.805 199.085 97.765 199.315 ;
        RECT 77.595 198.850 78.595 199.085 ;
        RECT 83.345 198.850 84.345 199.085 ;
        RECT 77.595 197.935 78.595 198.170 ;
        RECT 83.345 197.935 84.345 198.170 ;
        RECT 64.175 197.705 80.135 197.935 ;
        RECT 81.805 197.705 97.765 197.935 ;
        RECT 63.895 196.500 67.445 197.500 ;
        RECT 77.595 197.470 78.595 197.705 ;
        RECT 77.595 196.295 78.595 196.530 ;
        RECT 80.185 196.500 81.755 197.500 ;
        RECT 83.345 197.470 84.345 197.705 ;
        RECT 83.345 196.295 84.345 196.530 ;
        RECT 94.495 196.500 98.045 197.500 ;
        RECT 64.175 196.065 80.135 196.295 ;
        RECT 81.805 196.065 97.765 196.295 ;
        RECT 77.595 195.830 78.595 196.065 ;
        RECT 83.345 195.830 84.345 196.065 ;
        RECT 77.595 194.915 78.595 195.150 ;
        RECT 83.345 194.915 84.345 195.150 ;
        RECT 64.175 194.685 80.135 194.915 ;
        RECT 81.805 194.685 97.765 194.915 ;
        RECT 63.895 193.480 72.945 194.480 ;
        RECT 77.595 194.450 78.595 194.685 ;
        RECT 77.595 193.275 78.595 193.510 ;
        RECT 80.185 193.480 81.755 194.480 ;
        RECT 83.345 194.450 84.345 194.685 ;
        RECT 83.345 193.275 84.345 193.510 ;
        RECT 88.995 193.480 98.045 194.480 ;
        RECT 64.175 193.045 80.135 193.275 ;
        RECT 81.805 193.045 97.765 193.275 ;
        RECT 77.595 192.810 78.595 193.045 ;
        RECT 83.345 192.810 84.345 193.045 ;
        RECT 77.595 191.895 78.595 192.130 ;
        RECT 83.345 191.895 84.345 192.130 ;
        RECT 64.175 191.665 80.135 191.895 ;
        RECT 81.805 191.665 97.765 191.895 ;
        RECT 63.895 190.460 67.445 191.460 ;
        RECT 77.595 191.430 78.595 191.665 ;
        RECT 77.595 190.255 78.595 190.490 ;
        RECT 80.185 190.460 81.755 191.460 ;
        RECT 83.345 191.430 84.345 191.665 ;
        RECT 83.345 190.255 84.345 190.490 ;
        RECT 94.495 190.460 98.045 191.460 ;
        RECT 64.175 190.025 80.135 190.255 ;
        RECT 81.805 190.025 97.765 190.255 ;
        RECT 77.595 189.790 78.595 190.025 ;
        RECT 83.345 189.790 84.345 190.025 ;
        RECT 77.595 188.875 78.595 189.110 ;
        RECT 83.345 188.875 84.345 189.110 ;
        RECT 64.175 188.645 80.135 188.875 ;
        RECT 81.805 188.645 97.765 188.875 ;
        RECT 63.895 187.440 70.195 188.440 ;
        RECT 77.595 188.410 78.595 188.645 ;
        RECT 77.595 187.235 78.595 187.470 ;
        RECT 80.185 187.440 81.755 188.440 ;
        RECT 83.345 188.410 84.345 188.645 ;
        RECT 83.345 187.235 84.345 187.470 ;
        RECT 91.745 187.440 98.045 188.440 ;
        RECT 64.175 187.005 80.135 187.235 ;
        RECT 81.805 187.005 97.765 187.235 ;
        RECT 77.595 186.770 78.595 187.005 ;
        RECT 83.345 186.770 84.345 187.005 ;
        RECT 77.595 185.855 78.595 186.090 ;
        RECT 83.345 185.855 84.345 186.090 ;
        RECT 64.175 185.625 80.135 185.855 ;
        RECT 81.805 185.625 97.765 185.855 ;
        RECT 63.895 184.420 75.695 185.420 ;
        RECT 77.595 185.390 78.595 185.625 ;
        RECT 77.595 184.215 78.595 184.450 ;
        RECT 80.185 184.420 81.755 185.420 ;
        RECT 83.345 185.390 84.345 185.625 ;
        RECT 83.345 184.215 84.345 184.450 ;
        RECT 86.245 184.420 98.045 185.420 ;
        RECT 64.175 183.985 80.135 184.215 ;
        RECT 81.805 183.985 97.765 184.215 ;
        RECT 77.595 183.750 78.595 183.985 ;
        RECT 83.345 183.750 84.345 183.985 ;
        RECT 77.595 182.835 78.595 183.070 ;
        RECT 83.345 182.835 84.345 183.070 ;
        RECT 64.175 182.605 80.135 182.835 ;
        RECT 81.805 182.605 97.765 182.835 ;
        RECT 98.485 182.710 102.825 216.515 ;
        RECT 108.520 216.690 108.920 217.515 ;
        RECT 109.325 217.500 109.555 217.755 ;
        RECT 110.615 217.500 110.845 217.755 ;
        RECT 111.905 217.500 112.135 217.755 ;
        RECT 109.605 216.945 110.565 217.295 ;
        RECT 110.895 217.065 111.855 217.295 ;
        RECT 112.545 216.690 112.950 220.315 ;
        RECT 113.635 219.705 114.595 219.935 ;
        RECT 114.925 219.705 115.885 220.055 ;
        RECT 113.355 219.255 113.585 219.500 ;
        RECT 114.645 219.255 114.875 219.500 ;
        RECT 115.935 219.255 116.165 219.500 ;
        RECT 113.320 217.755 113.620 219.255 ;
        RECT 114.610 217.755 114.910 219.255 ;
        RECT 115.900 217.755 116.200 219.255 ;
        RECT 113.355 217.500 113.585 217.755 ;
        RECT 114.645 217.500 114.875 217.755 ;
        RECT 115.935 217.500 116.165 217.755 ;
        RECT 113.635 216.945 114.595 217.295 ;
        RECT 114.925 217.065 115.885 217.295 ;
        RECT 116.575 216.690 116.980 220.315 ;
        RECT 117.665 219.705 118.625 219.935 ;
        RECT 118.955 219.705 119.915 220.055 ;
        RECT 117.385 219.255 117.615 219.500 ;
        RECT 118.675 219.255 118.905 219.500 ;
        RECT 119.965 219.255 120.195 219.500 ;
        RECT 117.350 217.755 117.650 219.255 ;
        RECT 118.640 217.755 118.940 219.255 ;
        RECT 119.930 217.755 120.230 219.255 ;
        RECT 117.385 217.500 117.615 217.755 ;
        RECT 118.675 217.500 118.905 217.755 ;
        RECT 119.965 217.500 120.195 217.755 ;
        RECT 117.665 216.945 118.625 217.295 ;
        RECT 118.955 217.065 119.915 217.295 ;
        RECT 120.605 216.690 121.010 220.315 ;
        RECT 121.695 219.705 122.655 219.935 ;
        RECT 122.985 219.705 123.945 220.055 ;
        RECT 121.415 219.255 121.645 219.500 ;
        RECT 122.705 219.255 122.935 219.500 ;
        RECT 123.995 219.255 124.225 219.500 ;
        RECT 121.380 217.755 121.680 219.255 ;
        RECT 122.670 217.755 122.970 219.255 ;
        RECT 123.960 217.755 124.260 219.255 ;
        RECT 121.415 217.500 121.645 217.755 ;
        RECT 122.705 217.500 122.935 217.755 ;
        RECT 123.995 217.500 124.225 217.755 ;
        RECT 121.695 216.945 122.655 217.295 ;
        RECT 122.985 217.065 123.945 217.295 ;
        RECT 124.635 216.690 125.040 220.315 ;
        RECT 125.725 219.705 126.685 219.935 ;
        RECT 127.015 219.705 127.975 220.055 ;
        RECT 125.445 219.255 125.675 219.500 ;
        RECT 126.735 219.255 126.965 219.500 ;
        RECT 128.025 219.255 128.255 219.500 ;
        RECT 125.410 217.755 125.710 219.255 ;
        RECT 126.700 217.755 127.000 219.255 ;
        RECT 127.990 217.755 128.290 219.255 ;
        RECT 125.445 217.500 125.675 217.755 ;
        RECT 126.735 217.500 126.965 217.755 ;
        RECT 128.025 217.500 128.255 217.755 ;
        RECT 125.725 216.945 126.685 217.295 ;
        RECT 127.015 217.065 127.975 217.295 ;
        RECT 128.665 216.690 129.070 220.315 ;
        RECT 129.755 219.705 130.715 219.935 ;
        RECT 131.045 219.705 132.005 220.055 ;
        RECT 129.475 219.255 129.705 219.500 ;
        RECT 130.765 219.255 130.995 219.500 ;
        RECT 132.055 219.255 132.285 219.500 ;
        RECT 129.440 217.755 129.740 219.255 ;
        RECT 130.730 217.755 131.030 219.255 ;
        RECT 132.020 217.755 132.320 219.255 ;
        RECT 129.475 217.500 129.705 217.755 ;
        RECT 130.765 217.500 130.995 217.755 ;
        RECT 132.055 217.500 132.285 217.755 ;
        RECT 129.755 216.945 130.715 217.295 ;
        RECT 131.045 217.065 132.005 217.295 ;
        RECT 132.695 216.690 133.100 220.315 ;
        RECT 133.785 219.705 134.745 219.935 ;
        RECT 135.075 219.705 136.035 220.055 ;
        RECT 133.505 219.255 133.735 219.500 ;
        RECT 134.795 219.255 135.025 219.500 ;
        RECT 136.085 219.255 136.315 219.500 ;
        RECT 133.470 217.755 133.770 219.255 ;
        RECT 134.760 217.755 135.060 219.255 ;
        RECT 136.050 217.755 136.350 219.255 ;
        RECT 133.505 217.500 133.735 217.755 ;
        RECT 134.795 217.500 135.025 217.755 ;
        RECT 136.085 217.500 136.315 217.755 ;
        RECT 133.785 216.945 134.745 217.295 ;
        RECT 135.075 217.065 136.035 217.295 ;
        RECT 136.725 216.690 137.130 220.315 ;
        RECT 137.815 219.705 138.775 219.935 ;
        RECT 139.105 219.705 140.065 220.055 ;
        RECT 137.535 219.255 137.765 219.500 ;
        RECT 138.825 219.255 139.055 219.500 ;
        RECT 140.115 219.255 140.345 219.500 ;
        RECT 137.500 217.755 137.800 219.255 ;
        RECT 138.790 217.755 139.090 219.255 ;
        RECT 140.080 217.755 140.380 219.255 ;
        RECT 137.535 217.500 137.765 217.755 ;
        RECT 138.825 217.500 139.055 217.755 ;
        RECT 140.115 217.500 140.345 217.755 ;
        RECT 137.815 216.945 138.775 217.295 ;
        RECT 139.105 217.065 140.065 217.295 ;
        RECT 140.755 216.690 141.160 220.315 ;
        RECT 141.845 219.705 142.805 219.935 ;
        RECT 143.135 219.705 144.095 220.055 ;
        RECT 141.565 219.255 141.795 219.500 ;
        RECT 142.855 219.255 143.085 219.500 ;
        RECT 144.145 219.255 144.375 219.500 ;
        RECT 141.530 217.755 141.830 219.255 ;
        RECT 142.820 217.755 143.120 219.255 ;
        RECT 144.110 217.755 144.410 219.255 ;
        RECT 141.565 217.500 141.795 217.755 ;
        RECT 142.855 217.500 143.085 217.755 ;
        RECT 144.145 217.500 144.375 217.755 ;
        RECT 141.845 216.945 142.805 217.295 ;
        RECT 143.135 217.065 144.095 217.295 ;
        RECT 144.785 216.690 145.190 220.315 ;
        RECT 145.875 219.705 146.835 219.935 ;
        RECT 147.165 219.705 148.125 220.055 ;
        RECT 145.595 219.255 145.825 219.500 ;
        RECT 146.885 219.255 147.115 219.500 ;
        RECT 148.175 219.255 148.405 219.500 ;
        RECT 145.560 217.755 145.860 219.255 ;
        RECT 146.850 217.755 147.150 219.255 ;
        RECT 148.140 217.755 148.440 219.255 ;
        RECT 145.595 217.500 145.825 217.755 ;
        RECT 146.885 217.500 147.115 217.755 ;
        RECT 148.175 217.500 148.405 217.755 ;
        RECT 145.875 216.945 146.835 217.295 ;
        RECT 147.165 217.065 148.125 217.295 ;
        RECT 148.815 216.690 149.220 220.315 ;
        RECT 149.905 219.705 150.865 219.935 ;
        RECT 151.195 219.705 152.155 220.055 ;
        RECT 149.625 219.255 149.855 219.500 ;
        RECT 150.915 219.255 151.145 219.500 ;
        RECT 152.205 219.255 152.435 219.500 ;
        RECT 149.590 217.755 149.890 219.255 ;
        RECT 150.880 217.755 151.180 219.255 ;
        RECT 152.170 217.755 152.470 219.255 ;
        RECT 149.625 217.500 149.855 217.755 ;
        RECT 150.915 217.500 151.145 217.755 ;
        RECT 152.205 217.500 152.435 217.755 ;
        RECT 149.905 216.945 150.865 217.295 ;
        RECT 151.195 217.065 152.155 217.295 ;
        RECT 152.845 216.690 153.245 220.315 ;
        RECT 108.520 216.290 153.245 216.690 ;
        RECT 106.415 213.340 153.245 213.740 ;
        RECT 106.415 210.540 108.915 213.340 ;
        RECT 109.605 212.735 110.565 212.965 ;
        RECT 110.895 212.735 111.855 212.965 ;
        RECT 108.515 203.720 108.915 210.540 ;
        RECT 109.325 205.495 109.555 212.530 ;
        RECT 110.615 211.190 110.845 212.530 ;
        RECT 110.580 209.690 110.880 211.190 ;
        RECT 109.290 204.795 109.590 205.495 ;
        RECT 109.325 204.530 109.555 204.795 ;
        RECT 110.615 204.530 110.845 209.690 ;
        RECT 111.905 206.705 112.135 212.530 ;
        RECT 111.870 206.005 112.170 206.705 ;
        RECT 111.905 204.530 112.135 206.005 ;
        RECT 109.605 203.995 110.565 204.325 ;
        RECT 110.895 203.995 111.855 204.325 ;
        RECT 112.545 203.720 112.945 213.340 ;
        RECT 113.635 212.735 114.595 212.965 ;
        RECT 114.925 212.735 115.885 212.965 ;
        RECT 113.355 205.495 113.585 212.530 ;
        RECT 114.645 211.190 114.875 212.530 ;
        RECT 114.610 209.690 114.910 211.190 ;
        RECT 113.320 204.795 113.620 205.495 ;
        RECT 113.355 204.530 113.585 204.795 ;
        RECT 114.645 204.530 114.875 209.690 ;
        RECT 115.935 206.705 116.165 212.530 ;
        RECT 115.900 206.005 116.200 206.705 ;
        RECT 115.935 204.530 116.165 206.005 ;
        RECT 113.635 203.995 114.595 204.325 ;
        RECT 114.925 203.995 115.885 204.325 ;
        RECT 116.575 203.720 116.975 213.340 ;
        RECT 117.665 212.735 118.625 212.965 ;
        RECT 118.955 212.735 119.915 212.965 ;
        RECT 117.385 205.495 117.615 212.530 ;
        RECT 118.675 211.190 118.905 212.530 ;
        RECT 118.640 209.690 118.940 211.190 ;
        RECT 117.350 204.795 117.650 205.495 ;
        RECT 117.385 204.530 117.615 204.795 ;
        RECT 118.675 204.530 118.905 209.690 ;
        RECT 119.965 206.705 120.195 212.530 ;
        RECT 119.930 206.005 120.230 206.705 ;
        RECT 119.965 204.530 120.195 206.005 ;
        RECT 117.665 203.995 118.625 204.325 ;
        RECT 118.955 203.995 119.915 204.325 ;
        RECT 120.605 203.720 121.005 213.340 ;
        RECT 121.695 212.735 122.655 212.965 ;
        RECT 122.985 212.735 123.945 212.965 ;
        RECT 121.415 205.495 121.645 212.530 ;
        RECT 122.705 211.190 122.935 212.530 ;
        RECT 122.670 209.690 122.970 211.190 ;
        RECT 121.380 204.795 121.680 205.495 ;
        RECT 121.415 204.530 121.645 204.795 ;
        RECT 122.705 204.530 122.935 209.690 ;
        RECT 123.995 206.705 124.225 212.530 ;
        RECT 123.960 206.005 124.260 206.705 ;
        RECT 123.995 204.530 124.225 206.005 ;
        RECT 121.695 203.995 122.655 204.325 ;
        RECT 122.985 203.995 123.945 204.325 ;
        RECT 124.635 203.720 125.035 213.340 ;
        RECT 125.725 212.735 126.685 212.965 ;
        RECT 127.015 212.735 127.975 212.965 ;
        RECT 125.445 205.495 125.675 212.530 ;
        RECT 126.735 211.190 126.965 212.530 ;
        RECT 126.700 209.690 127.000 211.190 ;
        RECT 125.410 204.795 125.710 205.495 ;
        RECT 125.445 204.530 125.675 204.795 ;
        RECT 126.735 204.530 126.965 209.690 ;
        RECT 128.025 206.705 128.255 212.530 ;
        RECT 127.990 206.005 128.290 206.705 ;
        RECT 128.025 204.530 128.255 206.005 ;
        RECT 125.725 203.995 126.685 204.325 ;
        RECT 127.015 203.995 127.975 204.325 ;
        RECT 128.665 203.720 129.065 213.340 ;
        RECT 129.755 212.735 130.715 212.965 ;
        RECT 131.045 212.735 132.005 212.965 ;
        RECT 129.475 205.495 129.705 212.530 ;
        RECT 130.765 211.190 130.995 212.530 ;
        RECT 130.730 209.690 131.030 211.190 ;
        RECT 129.440 204.795 129.740 205.495 ;
        RECT 129.475 204.530 129.705 204.795 ;
        RECT 130.765 204.530 130.995 209.690 ;
        RECT 132.055 206.705 132.285 212.530 ;
        RECT 132.020 206.005 132.320 206.705 ;
        RECT 132.055 204.530 132.285 206.005 ;
        RECT 129.755 203.995 130.715 204.325 ;
        RECT 131.045 203.995 132.005 204.325 ;
        RECT 132.695 203.720 133.095 213.340 ;
        RECT 133.785 212.735 134.745 212.965 ;
        RECT 135.075 212.735 136.035 212.965 ;
        RECT 133.505 205.495 133.735 212.530 ;
        RECT 134.795 211.190 135.025 212.530 ;
        RECT 134.760 209.690 135.060 211.190 ;
        RECT 133.470 204.795 133.770 205.495 ;
        RECT 133.505 204.530 133.735 204.795 ;
        RECT 134.795 204.530 135.025 209.690 ;
        RECT 136.085 206.705 136.315 212.530 ;
        RECT 136.050 206.005 136.350 206.705 ;
        RECT 136.085 204.530 136.315 206.005 ;
        RECT 133.785 203.995 134.745 204.325 ;
        RECT 135.075 203.995 136.035 204.325 ;
        RECT 136.725 203.720 137.125 213.340 ;
        RECT 137.815 212.735 138.775 212.965 ;
        RECT 139.105 212.735 140.065 212.965 ;
        RECT 137.535 205.495 137.765 212.530 ;
        RECT 138.825 211.190 139.055 212.530 ;
        RECT 138.790 209.690 139.090 211.190 ;
        RECT 137.500 204.795 137.800 205.495 ;
        RECT 137.535 204.530 137.765 204.795 ;
        RECT 138.825 204.530 139.055 209.690 ;
        RECT 140.115 206.705 140.345 212.530 ;
        RECT 140.080 206.005 140.380 206.705 ;
        RECT 140.115 204.530 140.345 206.005 ;
        RECT 137.815 203.995 138.775 204.325 ;
        RECT 139.105 203.995 140.065 204.325 ;
        RECT 140.755 203.720 141.155 213.340 ;
        RECT 141.845 212.735 142.805 212.965 ;
        RECT 143.135 212.735 144.095 212.965 ;
        RECT 141.565 205.495 141.795 212.530 ;
        RECT 142.855 211.190 143.085 212.530 ;
        RECT 142.820 209.690 143.120 211.190 ;
        RECT 141.530 204.795 141.830 205.495 ;
        RECT 141.565 204.530 141.795 204.795 ;
        RECT 142.855 204.530 143.085 209.690 ;
        RECT 144.145 206.705 144.375 212.530 ;
        RECT 144.110 206.005 144.410 206.705 ;
        RECT 144.145 204.530 144.375 206.005 ;
        RECT 141.845 203.995 142.805 204.325 ;
        RECT 143.135 203.995 144.095 204.325 ;
        RECT 144.785 203.720 145.185 213.340 ;
        RECT 145.875 212.735 146.835 212.965 ;
        RECT 147.165 212.735 148.125 212.965 ;
        RECT 145.595 205.495 145.825 212.530 ;
        RECT 146.885 211.190 147.115 212.530 ;
        RECT 146.850 209.690 147.150 211.190 ;
        RECT 145.560 204.795 145.860 205.495 ;
        RECT 145.595 204.530 145.825 204.795 ;
        RECT 146.885 204.530 147.115 209.690 ;
        RECT 148.175 206.705 148.405 212.530 ;
        RECT 148.140 206.005 148.440 206.705 ;
        RECT 148.175 204.530 148.405 206.005 ;
        RECT 145.875 203.995 146.835 204.325 ;
        RECT 147.165 203.995 148.125 204.325 ;
        RECT 148.815 203.720 149.215 213.340 ;
        RECT 149.905 212.735 150.865 212.965 ;
        RECT 151.195 212.735 152.155 212.965 ;
        RECT 149.625 205.495 149.855 212.530 ;
        RECT 150.915 211.190 151.145 212.530 ;
        RECT 150.880 209.690 151.180 211.190 ;
        RECT 149.590 204.795 149.890 205.495 ;
        RECT 149.625 204.530 149.855 204.795 ;
        RECT 150.915 204.530 151.145 209.690 ;
        RECT 152.205 206.705 152.435 212.530 ;
        RECT 152.170 206.005 152.470 206.705 ;
        RECT 152.205 204.530 152.435 206.005 ;
        RECT 149.905 203.995 150.865 204.325 ;
        RECT 151.195 203.995 152.155 204.325 ;
        RECT 152.845 203.720 153.245 213.340 ;
        RECT 108.515 203.320 153.245 203.720 ;
        RECT 162.095 201.250 236.155 201.730 ;
        RECT 165.385 201.050 165.705 201.110 ;
        RECT 166.320 201.050 166.610 201.095 ;
        RECT 108.515 200.625 153.245 201.025 ;
        RECT 165.385 200.910 166.610 201.050 ;
        RECT 165.385 200.850 165.705 200.910 ;
        RECT 166.320 200.865 166.610 200.910 ;
        RECT 175.045 201.050 175.365 201.110 ;
        RECT 176.440 201.050 176.730 201.095 ;
        RECT 175.045 200.910 176.730 201.050 ;
        RECT 175.045 200.850 175.365 200.910 ;
        RECT 176.440 200.865 176.730 200.910 ;
        RECT 184.705 201.050 185.025 201.110 ;
        RECT 186.100 201.050 186.390 201.095 ;
        RECT 184.705 200.910 186.390 201.050 ;
        RECT 184.705 200.850 185.025 200.910 ;
        RECT 186.100 200.865 186.390 200.910 ;
        RECT 194.365 201.050 194.685 201.110 ;
        RECT 195.760 201.050 196.050 201.095 ;
        RECT 194.365 200.910 196.050 201.050 ;
        RECT 194.365 200.850 194.685 200.910 ;
        RECT 195.760 200.865 196.050 200.910 ;
        RECT 204.025 201.050 204.345 201.110 ;
        RECT 205.420 201.050 205.710 201.095 ;
        RECT 204.025 200.910 205.710 201.050 ;
        RECT 204.025 200.850 204.345 200.910 ;
        RECT 205.420 200.865 205.710 200.910 ;
        RECT 213.685 201.050 214.005 201.110 ;
        RECT 215.080 201.050 215.370 201.095 ;
        RECT 213.685 200.910 215.370 201.050 ;
        RECT 213.685 200.850 214.005 200.910 ;
        RECT 215.080 200.865 215.370 200.910 ;
        RECT 223.345 201.050 223.665 201.110 ;
        RECT 224.740 201.050 225.030 201.095 ;
        RECT 223.345 200.910 225.030 201.050 ;
        RECT 223.345 200.850 223.665 200.910 ;
        RECT 224.740 200.865 225.030 200.910 ;
        RECT 233.005 201.050 233.325 201.110 ;
        RECT 233.940 201.050 234.230 201.095 ;
        RECT 233.005 200.910 234.230 201.050 ;
        RECT 233.005 200.850 233.325 200.910 ;
        RECT 233.940 200.865 234.230 200.910 ;
        RECT 108.515 195.095 108.915 200.625 ;
        RECT 109.735 200.250 110.435 200.320 ;
        RECT 111.025 200.250 111.725 200.320 ;
        RECT 109.605 200.020 110.565 200.250 ;
        RECT 110.895 200.020 111.855 200.250 ;
        RECT 109.325 199.635 109.555 199.860 ;
        RECT 109.290 198.935 109.590 199.635 ;
        RECT 110.615 198.955 110.845 199.860 ;
        RECT 111.905 199.635 112.135 199.860 ;
        RECT 109.325 195.860 109.555 198.935 ;
        RECT 110.580 196.855 110.880 198.955 ;
        RECT 111.870 198.935 112.170 199.635 ;
        RECT 110.615 195.860 110.845 196.855 ;
        RECT 111.905 195.860 112.135 198.935 ;
        RECT 109.605 195.470 110.565 195.700 ;
        RECT 110.895 195.470 111.855 195.700 ;
        RECT 112.545 195.095 112.945 200.625 ;
        RECT 113.765 200.250 114.465 200.320 ;
        RECT 115.055 200.250 115.755 200.320 ;
        RECT 113.635 200.020 114.595 200.250 ;
        RECT 114.925 200.020 115.885 200.250 ;
        RECT 113.355 199.635 113.585 199.860 ;
        RECT 113.320 198.935 113.620 199.635 ;
        RECT 114.645 198.955 114.875 199.860 ;
        RECT 115.935 199.635 116.165 199.860 ;
        RECT 113.355 195.860 113.585 198.935 ;
        RECT 114.610 196.855 114.910 198.955 ;
        RECT 115.900 198.935 116.200 199.635 ;
        RECT 114.645 195.860 114.875 196.855 ;
        RECT 115.935 195.860 116.165 198.935 ;
        RECT 113.635 195.470 114.595 195.700 ;
        RECT 114.925 195.470 115.885 195.700 ;
        RECT 116.575 195.095 116.975 200.625 ;
        RECT 117.795 200.250 118.495 200.320 ;
        RECT 119.085 200.250 119.785 200.320 ;
        RECT 117.665 200.020 118.625 200.250 ;
        RECT 118.955 200.020 119.915 200.250 ;
        RECT 117.385 199.635 117.615 199.860 ;
        RECT 117.350 198.935 117.650 199.635 ;
        RECT 118.675 198.955 118.905 199.860 ;
        RECT 119.965 199.635 120.195 199.860 ;
        RECT 117.385 195.860 117.615 198.935 ;
        RECT 118.640 196.855 118.940 198.955 ;
        RECT 119.930 198.935 120.230 199.635 ;
        RECT 118.675 195.860 118.905 196.855 ;
        RECT 119.965 195.860 120.195 198.935 ;
        RECT 117.665 195.470 118.625 195.700 ;
        RECT 118.955 195.470 119.915 195.700 ;
        RECT 120.605 195.095 121.005 200.625 ;
        RECT 121.825 200.250 122.525 200.320 ;
        RECT 123.115 200.250 123.815 200.320 ;
        RECT 121.695 200.020 122.655 200.250 ;
        RECT 122.985 200.020 123.945 200.250 ;
        RECT 121.415 199.635 121.645 199.860 ;
        RECT 121.380 198.935 121.680 199.635 ;
        RECT 122.705 198.955 122.935 199.860 ;
        RECT 123.995 199.635 124.225 199.860 ;
        RECT 121.415 195.860 121.645 198.935 ;
        RECT 122.670 196.855 122.970 198.955 ;
        RECT 123.960 198.935 124.260 199.635 ;
        RECT 122.705 195.860 122.935 196.855 ;
        RECT 123.995 195.860 124.225 198.935 ;
        RECT 121.695 195.470 122.655 195.700 ;
        RECT 122.985 195.470 123.945 195.700 ;
        RECT 124.635 195.095 125.035 200.625 ;
        RECT 125.855 200.250 126.555 200.320 ;
        RECT 127.145 200.250 127.845 200.320 ;
        RECT 125.725 200.020 126.685 200.250 ;
        RECT 127.015 200.020 127.975 200.250 ;
        RECT 125.445 199.635 125.675 199.860 ;
        RECT 125.410 198.935 125.710 199.635 ;
        RECT 126.735 198.955 126.965 199.860 ;
        RECT 128.025 199.635 128.255 199.860 ;
        RECT 125.445 195.860 125.675 198.935 ;
        RECT 126.700 196.855 127.000 198.955 ;
        RECT 127.990 198.935 128.290 199.635 ;
        RECT 126.735 195.860 126.965 196.855 ;
        RECT 128.025 195.860 128.255 198.935 ;
        RECT 125.725 195.470 126.685 195.700 ;
        RECT 127.015 195.470 127.975 195.700 ;
        RECT 128.665 195.095 129.065 200.625 ;
        RECT 129.885 200.250 130.585 200.320 ;
        RECT 131.175 200.250 131.875 200.320 ;
        RECT 129.755 200.020 130.715 200.250 ;
        RECT 131.045 200.020 132.005 200.250 ;
        RECT 129.475 199.635 129.705 199.860 ;
        RECT 129.440 198.935 129.740 199.635 ;
        RECT 130.765 198.955 130.995 199.860 ;
        RECT 132.055 199.635 132.285 199.860 ;
        RECT 129.475 195.860 129.705 198.935 ;
        RECT 130.730 196.855 131.030 198.955 ;
        RECT 132.020 198.935 132.320 199.635 ;
        RECT 130.765 195.860 130.995 196.855 ;
        RECT 132.055 195.860 132.285 198.935 ;
        RECT 129.755 195.470 130.715 195.700 ;
        RECT 131.045 195.470 132.005 195.700 ;
        RECT 132.695 195.095 133.095 200.625 ;
        RECT 133.915 200.250 134.615 200.320 ;
        RECT 135.205 200.250 135.905 200.320 ;
        RECT 133.785 200.020 134.745 200.250 ;
        RECT 135.075 200.020 136.035 200.250 ;
        RECT 133.505 199.635 133.735 199.860 ;
        RECT 133.470 198.935 133.770 199.635 ;
        RECT 134.795 198.955 135.025 199.860 ;
        RECT 136.085 199.635 136.315 199.860 ;
        RECT 133.505 195.860 133.735 198.935 ;
        RECT 134.760 196.855 135.060 198.955 ;
        RECT 136.050 198.935 136.350 199.635 ;
        RECT 134.795 195.860 135.025 196.855 ;
        RECT 136.085 195.860 136.315 198.935 ;
        RECT 133.785 195.470 134.745 195.700 ;
        RECT 135.075 195.470 136.035 195.700 ;
        RECT 136.725 195.095 137.125 200.625 ;
        RECT 137.945 200.250 138.645 200.320 ;
        RECT 139.235 200.250 139.935 200.320 ;
        RECT 137.815 200.020 138.775 200.250 ;
        RECT 139.105 200.020 140.065 200.250 ;
        RECT 137.535 199.635 137.765 199.860 ;
        RECT 137.500 198.935 137.800 199.635 ;
        RECT 138.825 198.955 139.055 199.860 ;
        RECT 140.115 199.635 140.345 199.860 ;
        RECT 137.535 195.860 137.765 198.935 ;
        RECT 138.790 196.855 139.090 198.955 ;
        RECT 140.080 198.935 140.380 199.635 ;
        RECT 138.825 195.860 139.055 196.855 ;
        RECT 140.115 195.860 140.345 198.935 ;
        RECT 137.815 195.470 138.775 195.700 ;
        RECT 139.105 195.470 140.065 195.700 ;
        RECT 140.755 195.095 141.155 200.625 ;
        RECT 141.975 200.250 142.675 200.320 ;
        RECT 143.265 200.250 143.965 200.320 ;
        RECT 141.845 200.020 142.805 200.250 ;
        RECT 143.135 200.020 144.095 200.250 ;
        RECT 141.565 199.635 141.795 199.860 ;
        RECT 141.530 198.935 141.830 199.635 ;
        RECT 142.855 198.955 143.085 199.860 ;
        RECT 144.145 199.635 144.375 199.860 ;
        RECT 141.565 195.860 141.795 198.935 ;
        RECT 142.820 196.855 143.120 198.955 ;
        RECT 144.110 198.935 144.410 199.635 ;
        RECT 142.855 195.860 143.085 196.855 ;
        RECT 144.145 195.860 144.375 198.935 ;
        RECT 141.845 195.470 142.805 195.700 ;
        RECT 143.135 195.470 144.095 195.700 ;
        RECT 144.785 195.095 145.185 200.625 ;
        RECT 146.005 200.250 146.705 200.320 ;
        RECT 147.295 200.250 147.995 200.320 ;
        RECT 145.875 200.020 146.835 200.250 ;
        RECT 147.165 200.020 148.125 200.250 ;
        RECT 145.595 199.635 145.825 199.860 ;
        RECT 145.560 198.935 145.860 199.635 ;
        RECT 146.885 198.955 147.115 199.860 ;
        RECT 148.175 199.635 148.405 199.860 ;
        RECT 145.595 195.860 145.825 198.935 ;
        RECT 146.850 196.855 147.150 198.955 ;
        RECT 148.140 198.935 148.440 199.635 ;
        RECT 146.885 195.860 147.115 196.855 ;
        RECT 148.175 195.860 148.405 198.935 ;
        RECT 145.875 195.470 146.835 195.700 ;
        RECT 147.165 195.470 148.125 195.700 ;
        RECT 148.815 195.095 149.215 200.625 ;
        RECT 150.035 200.250 150.735 200.320 ;
        RECT 151.325 200.250 152.025 200.320 ;
        RECT 149.905 200.020 150.865 200.250 ;
        RECT 151.195 200.020 152.155 200.250 ;
        RECT 149.625 199.635 149.855 199.860 ;
        RECT 149.590 198.935 149.890 199.635 ;
        RECT 150.915 198.955 151.145 199.860 ;
        RECT 152.205 199.635 152.435 199.860 ;
        RECT 149.625 195.860 149.855 198.935 ;
        RECT 150.880 196.855 151.180 198.955 ;
        RECT 152.170 198.935 152.470 199.635 ;
        RECT 150.915 195.860 151.145 196.855 ;
        RECT 152.205 195.860 152.435 198.935 ;
        RECT 149.905 195.470 150.865 195.700 ;
        RECT 151.195 195.470 152.155 195.700 ;
        RECT 152.845 195.095 153.245 200.625 ;
        RECT 167.225 199.830 167.545 200.090 ;
        RECT 175.505 199.830 175.825 200.090 ;
        RECT 185.165 199.830 185.485 200.090 ;
        RECT 194.825 199.830 195.145 200.090 ;
        RECT 204.485 199.830 204.805 200.090 ;
        RECT 214.145 199.830 214.465 200.090 ;
        RECT 223.805 199.830 224.125 200.090 ;
        RECT 233.005 199.830 233.325 200.090 ;
        RECT 164.005 199.490 164.325 199.750 ;
        RECT 164.940 199.690 165.230 199.735 ;
        RECT 175.045 199.690 175.365 199.750 ;
        RECT 164.940 199.550 175.365 199.690 ;
        RECT 164.940 199.505 165.230 199.550 ;
        RECT 175.045 199.490 175.365 199.550 ;
        RECT 162.095 198.530 236.155 199.010 ;
        RECT 162.095 195.810 236.155 196.290 ;
        RECT 108.515 194.695 153.245 195.095 ;
        RECT 175.045 194.930 175.365 194.990 ;
        RECT 199.425 194.930 199.745 194.990 ;
        RECT 175.045 194.790 199.745 194.930 ;
        RECT 175.045 194.730 175.365 194.790 ;
        RECT 199.425 194.730 199.745 194.790 ;
        RECT 108.515 185.165 108.915 194.695 ;
        RECT 109.605 194.320 110.305 194.390 ;
        RECT 111.155 194.320 111.855 194.390 ;
        RECT 109.605 194.090 110.565 194.320 ;
        RECT 110.895 194.090 111.855 194.320 ;
        RECT 109.325 192.835 109.555 193.930 ;
        RECT 109.290 191.335 109.590 192.835 ;
        RECT 109.325 185.930 109.555 191.335 ;
        RECT 110.615 189.090 110.845 193.930 ;
        RECT 111.905 192.835 112.135 193.930 ;
        RECT 111.870 191.335 112.170 192.835 ;
        RECT 110.580 187.590 110.880 189.090 ;
        RECT 110.615 185.930 110.845 187.590 ;
        RECT 111.905 185.930 112.135 191.335 ;
        RECT 109.605 185.540 110.565 185.770 ;
        RECT 110.895 185.540 111.855 185.770 ;
        RECT 112.545 185.165 112.945 194.695 ;
        RECT 113.635 194.320 114.335 194.390 ;
        RECT 115.185 194.320 115.885 194.390 ;
        RECT 113.635 194.090 114.595 194.320 ;
        RECT 114.925 194.090 115.885 194.320 ;
        RECT 113.355 192.835 113.585 193.930 ;
        RECT 113.320 191.335 113.620 192.835 ;
        RECT 113.355 185.930 113.585 191.335 ;
        RECT 114.645 189.090 114.875 193.930 ;
        RECT 115.935 192.835 116.165 193.930 ;
        RECT 115.900 191.335 116.200 192.835 ;
        RECT 114.610 187.590 114.910 189.090 ;
        RECT 114.645 185.930 114.875 187.590 ;
        RECT 115.935 185.930 116.165 191.335 ;
        RECT 113.635 185.540 114.595 185.770 ;
        RECT 114.925 185.540 115.885 185.770 ;
        RECT 116.575 185.165 116.975 194.695 ;
        RECT 117.665 194.320 118.365 194.390 ;
        RECT 119.215 194.320 119.915 194.390 ;
        RECT 117.665 194.090 118.625 194.320 ;
        RECT 118.955 194.090 119.915 194.320 ;
        RECT 117.385 192.835 117.615 193.930 ;
        RECT 117.350 191.335 117.650 192.835 ;
        RECT 117.385 185.930 117.615 191.335 ;
        RECT 118.675 189.090 118.905 193.930 ;
        RECT 119.965 192.835 120.195 193.930 ;
        RECT 119.930 191.335 120.230 192.835 ;
        RECT 118.640 187.590 118.940 189.090 ;
        RECT 118.675 185.930 118.905 187.590 ;
        RECT 119.965 185.930 120.195 191.335 ;
        RECT 117.665 185.540 118.625 185.770 ;
        RECT 118.955 185.540 119.915 185.770 ;
        RECT 120.605 185.165 121.005 194.695 ;
        RECT 121.695 194.320 122.395 194.390 ;
        RECT 123.245 194.320 123.945 194.390 ;
        RECT 121.695 194.090 122.655 194.320 ;
        RECT 122.985 194.090 123.945 194.320 ;
        RECT 121.415 192.835 121.645 193.930 ;
        RECT 121.380 191.335 121.680 192.835 ;
        RECT 121.415 185.930 121.645 191.335 ;
        RECT 122.705 189.090 122.935 193.930 ;
        RECT 123.995 192.835 124.225 193.930 ;
        RECT 123.960 191.335 124.260 192.835 ;
        RECT 122.670 187.590 122.970 189.090 ;
        RECT 122.705 185.930 122.935 187.590 ;
        RECT 123.995 185.930 124.225 191.335 ;
        RECT 121.695 185.540 122.655 185.770 ;
        RECT 122.985 185.540 123.945 185.770 ;
        RECT 124.635 185.165 125.035 194.695 ;
        RECT 125.725 194.320 126.425 194.390 ;
        RECT 127.275 194.320 127.975 194.390 ;
        RECT 125.725 194.090 126.685 194.320 ;
        RECT 127.015 194.090 127.975 194.320 ;
        RECT 125.445 192.835 125.675 193.930 ;
        RECT 125.410 191.335 125.710 192.835 ;
        RECT 125.445 185.930 125.675 191.335 ;
        RECT 126.735 189.090 126.965 193.930 ;
        RECT 128.025 192.835 128.255 193.930 ;
        RECT 127.990 191.335 128.290 192.835 ;
        RECT 126.700 187.590 127.000 189.090 ;
        RECT 126.735 185.930 126.965 187.590 ;
        RECT 128.025 185.930 128.255 191.335 ;
        RECT 125.725 185.540 126.685 185.770 ;
        RECT 127.015 185.540 127.975 185.770 ;
        RECT 128.665 185.165 129.065 194.695 ;
        RECT 129.755 194.320 130.455 194.390 ;
        RECT 131.305 194.320 132.005 194.390 ;
        RECT 129.755 194.090 130.715 194.320 ;
        RECT 131.045 194.090 132.005 194.320 ;
        RECT 129.475 192.835 129.705 193.930 ;
        RECT 129.440 191.335 129.740 192.835 ;
        RECT 129.475 185.930 129.705 191.335 ;
        RECT 130.765 189.090 130.995 193.930 ;
        RECT 132.055 192.835 132.285 193.930 ;
        RECT 132.020 191.335 132.320 192.835 ;
        RECT 130.730 187.590 131.030 189.090 ;
        RECT 130.765 185.930 130.995 187.590 ;
        RECT 132.055 185.930 132.285 191.335 ;
        RECT 129.755 185.540 130.715 185.770 ;
        RECT 131.045 185.540 132.005 185.770 ;
        RECT 132.695 185.165 133.095 194.695 ;
        RECT 133.785 194.320 134.485 194.390 ;
        RECT 135.335 194.320 136.035 194.390 ;
        RECT 133.785 194.090 134.745 194.320 ;
        RECT 135.075 194.090 136.035 194.320 ;
        RECT 133.505 192.835 133.735 193.930 ;
        RECT 133.470 191.335 133.770 192.835 ;
        RECT 133.505 185.930 133.735 191.335 ;
        RECT 134.795 189.090 135.025 193.930 ;
        RECT 136.085 192.835 136.315 193.930 ;
        RECT 136.050 191.335 136.350 192.835 ;
        RECT 134.760 187.590 135.060 189.090 ;
        RECT 134.795 185.930 135.025 187.590 ;
        RECT 136.085 185.930 136.315 191.335 ;
        RECT 133.785 185.540 134.745 185.770 ;
        RECT 135.075 185.540 136.035 185.770 ;
        RECT 136.725 185.165 137.125 194.695 ;
        RECT 137.815 194.320 138.515 194.390 ;
        RECT 139.365 194.320 140.065 194.390 ;
        RECT 137.815 194.090 138.775 194.320 ;
        RECT 139.105 194.090 140.065 194.320 ;
        RECT 137.535 192.835 137.765 193.930 ;
        RECT 137.500 191.335 137.800 192.835 ;
        RECT 137.535 185.930 137.765 191.335 ;
        RECT 138.825 189.090 139.055 193.930 ;
        RECT 140.115 192.835 140.345 193.930 ;
        RECT 140.080 191.335 140.380 192.835 ;
        RECT 138.790 187.590 139.090 189.090 ;
        RECT 138.825 185.930 139.055 187.590 ;
        RECT 140.115 185.930 140.345 191.335 ;
        RECT 137.815 185.540 138.775 185.770 ;
        RECT 139.105 185.540 140.065 185.770 ;
        RECT 140.755 185.165 141.155 194.695 ;
        RECT 141.845 194.320 142.545 194.390 ;
        RECT 143.395 194.320 144.095 194.390 ;
        RECT 141.845 194.090 142.805 194.320 ;
        RECT 143.135 194.090 144.095 194.320 ;
        RECT 141.565 192.835 141.795 193.930 ;
        RECT 141.530 191.335 141.830 192.835 ;
        RECT 141.565 185.930 141.795 191.335 ;
        RECT 142.855 189.090 143.085 193.930 ;
        RECT 144.145 192.835 144.375 193.930 ;
        RECT 144.110 191.335 144.410 192.835 ;
        RECT 142.820 187.590 143.120 189.090 ;
        RECT 142.855 185.930 143.085 187.590 ;
        RECT 144.145 185.930 144.375 191.335 ;
        RECT 141.845 185.540 142.805 185.770 ;
        RECT 143.135 185.540 144.095 185.770 ;
        RECT 144.785 185.165 145.185 194.695 ;
        RECT 145.875 194.320 146.575 194.390 ;
        RECT 147.425 194.320 148.125 194.390 ;
        RECT 145.875 194.090 146.835 194.320 ;
        RECT 147.165 194.090 148.125 194.320 ;
        RECT 145.595 192.835 145.825 193.930 ;
        RECT 145.560 191.335 145.860 192.835 ;
        RECT 145.595 185.930 145.825 191.335 ;
        RECT 146.885 189.090 147.115 193.930 ;
        RECT 148.175 192.835 148.405 193.930 ;
        RECT 148.140 191.335 148.440 192.835 ;
        RECT 146.850 187.590 147.150 189.090 ;
        RECT 146.885 185.930 147.115 187.590 ;
        RECT 148.175 185.930 148.405 191.335 ;
        RECT 145.875 185.540 146.835 185.770 ;
        RECT 147.165 185.540 148.125 185.770 ;
        RECT 148.815 185.165 149.215 194.695 ;
        RECT 149.905 194.320 150.605 194.390 ;
        RECT 151.455 194.320 152.155 194.390 ;
        RECT 149.905 194.090 150.865 194.320 ;
        RECT 151.195 194.090 152.155 194.320 ;
        RECT 149.625 192.835 149.855 193.930 ;
        RECT 149.590 191.335 149.890 192.835 ;
        RECT 149.625 185.930 149.855 191.335 ;
        RECT 150.915 189.090 151.145 193.930 ;
        RECT 152.205 192.835 152.435 193.930 ;
        RECT 152.170 191.335 152.470 192.835 ;
        RECT 150.880 187.590 151.180 189.090 ;
        RECT 150.915 185.930 151.145 187.590 ;
        RECT 152.205 185.930 152.435 191.335 ;
        RECT 152.845 187.965 153.245 194.695 ;
        RECT 176.440 194.590 176.730 194.635 ;
        RECT 176.885 194.590 177.205 194.650 ;
        RECT 176.440 194.450 177.205 194.590 ;
        RECT 176.440 194.405 176.730 194.450 ;
        RECT 176.885 194.390 177.205 194.450 ;
        RECT 178.725 194.250 179.045 194.310 ;
        RECT 205.405 194.250 205.725 194.310 ;
        RECT 178.725 194.110 205.725 194.250 ;
        RECT 178.725 194.050 179.045 194.110 ;
        RECT 205.405 194.050 205.725 194.110 ;
        RECT 173.205 193.910 173.525 193.970 ;
        RECT 175.980 193.910 176.270 193.955 ;
        RECT 187.005 193.910 187.325 193.970 ;
        RECT 173.205 193.770 187.325 193.910 ;
        RECT 173.205 193.710 173.525 193.770 ;
        RECT 175.980 193.725 176.270 193.770 ;
        RECT 187.005 193.710 187.325 193.770 ;
        RECT 162.095 193.090 236.155 193.570 ;
        RECT 178.725 192.890 179.045 192.950 ;
        RECT 173.065 192.750 179.045 192.890 ;
        RECT 168.145 192.210 168.465 192.270 ;
        RECT 170.920 192.210 171.210 192.255 ;
        RECT 168.145 192.070 171.210 192.210 ;
        RECT 168.145 192.010 168.465 192.070 ;
        RECT 170.920 192.025 171.210 192.070 ;
        RECT 172.300 192.210 172.590 192.255 ;
        RECT 173.065 192.210 173.205 192.750 ;
        RECT 178.725 192.690 179.045 192.750 ;
        RECT 184.720 192.890 185.010 192.935 ;
        RECT 185.165 192.890 185.485 192.950 ;
        RECT 184.720 192.750 185.485 192.890 ;
        RECT 184.720 192.705 185.010 192.750 ;
        RECT 185.165 192.690 185.485 192.750 ;
        RECT 194.380 192.890 194.670 192.935 ;
        RECT 194.825 192.890 195.145 192.950 ;
        RECT 194.380 192.750 195.145 192.890 ;
        RECT 194.380 192.705 194.670 192.750 ;
        RECT 194.825 192.690 195.145 192.750 ;
        RECT 204.485 192.690 204.805 192.950 ;
        RECT 177.360 192.550 177.650 192.595 ;
        RECT 189.765 192.550 190.085 192.610 ;
        RECT 174.675 192.410 190.085 192.550 ;
        RECT 174.675 192.255 174.815 192.410 ;
        RECT 177.360 192.365 177.650 192.410 ;
        RECT 189.765 192.350 190.085 192.410 ;
        RECT 172.300 192.070 173.205 192.210 ;
        RECT 172.300 192.025 172.590 192.070 ;
        RECT 174.600 192.025 174.890 192.255 ;
        RECT 175.045 192.210 175.365 192.270 ;
        RECT 175.520 192.210 175.810 192.255 ;
        RECT 175.045 192.070 175.810 192.210 ;
        RECT 175.045 192.010 175.365 192.070 ;
        RECT 175.520 192.025 175.810 192.070 ;
        RECT 175.965 192.210 176.285 192.270 ;
        RECT 177.820 192.210 178.110 192.255 ;
        RECT 175.965 192.070 178.110 192.210 ;
        RECT 175.965 192.010 176.285 192.070 ;
        RECT 177.820 192.025 178.110 192.070 ;
        RECT 180.580 192.025 180.870 192.255 ;
        RECT 182.865 192.210 183.185 192.270 ;
        RECT 185.640 192.210 185.930 192.255 ;
        RECT 182.865 192.070 185.930 192.210 ;
        RECT 176.425 191.870 176.745 191.930 ;
        RECT 180.655 191.870 180.795 192.025 ;
        RECT 182.865 192.010 183.185 192.070 ;
        RECT 185.640 192.025 185.930 192.070 ;
        RECT 187.005 192.010 187.325 192.270 ;
        RECT 189.305 192.210 189.625 192.270 ;
        RECT 195.300 192.210 195.590 192.255 ;
        RECT 189.305 192.070 195.590 192.210 ;
        RECT 189.305 192.010 189.625 192.070 ;
        RECT 195.300 192.025 195.590 192.070 ;
        RECT 198.505 192.210 198.825 192.270 ;
        RECT 203.580 192.210 203.870 192.255 ;
        RECT 198.505 192.070 203.870 192.210 ;
        RECT 198.505 192.010 198.825 192.070 ;
        RECT 203.580 192.025 203.870 192.070 ;
        RECT 176.425 191.730 180.795 191.870 ;
        RECT 187.095 191.870 187.235 192.010 ;
        RECT 196.680 191.870 196.970 191.915 ;
        RECT 202.200 191.870 202.490 191.915 ;
        RECT 211.385 191.870 211.705 191.930 ;
        RECT 187.095 191.730 211.705 191.870 ;
        RECT 176.425 191.670 176.745 191.730 ;
        RECT 196.680 191.685 196.970 191.730 ;
        RECT 202.200 191.685 202.490 191.730 ;
        RECT 211.385 191.670 211.705 191.730 ;
        RECT 171.365 191.330 171.685 191.590 ;
        RECT 166.305 191.190 166.625 191.250 ;
        RECT 170.000 191.190 170.290 191.235 ;
        RECT 166.305 191.050 170.290 191.190 ;
        RECT 166.305 190.990 166.625 191.050 ;
        RECT 170.000 191.005 170.290 191.050 ;
        RECT 171.825 191.190 172.145 191.250 ;
        RECT 173.680 191.190 173.970 191.235 ;
        RECT 171.825 191.050 173.970 191.190 ;
        RECT 171.825 190.990 172.145 191.050 ;
        RECT 173.680 191.005 173.970 191.050 ;
        RECT 179.645 190.990 179.965 191.250 ;
        RECT 186.545 190.990 186.865 191.250 ;
        RECT 196.205 190.990 196.525 191.250 ;
        RECT 202.645 190.990 202.965 191.250 ;
        RECT 162.095 190.370 236.155 190.850 ;
        RECT 164.480 190.170 164.770 190.215 ;
        RECT 175.965 190.170 176.285 190.230 ;
        RECT 164.480 190.030 176.285 190.170 ;
        RECT 164.480 189.985 164.770 190.030 ;
        RECT 175.965 189.970 176.285 190.030 ;
        RECT 178.740 190.170 179.030 190.215 ;
        RECT 178.740 190.030 189.075 190.170 ;
        RECT 178.740 189.985 179.030 190.030 ;
        RECT 169.080 189.645 169.370 189.875 ;
        RECT 169.540 189.830 169.830 189.875 ;
        RECT 169.540 189.690 173.895 189.830 ;
        RECT 169.540 189.645 169.830 189.690 ;
        RECT 169.155 189.490 169.295 189.645 ;
        RECT 173.755 189.490 173.895 189.690 ;
        RECT 182.865 189.630 183.185 189.890 ;
        RECT 188.385 189.830 188.705 189.890 ;
        RECT 186.175 189.690 188.705 189.830 ;
        RECT 188.935 189.830 189.075 190.030 ;
        RECT 189.305 189.970 189.625 190.230 ;
        RECT 189.765 190.170 190.085 190.230 ;
        RECT 213.700 190.170 213.990 190.215 ;
        RECT 214.145 190.170 214.465 190.230 ;
        RECT 189.765 190.030 199.195 190.170 ;
        RECT 189.765 189.970 190.085 190.030 ;
        RECT 197.585 189.830 197.905 189.890 ;
        RECT 188.935 189.690 197.905 189.830 ;
        RECT 169.155 189.350 172.515 189.490 ;
        RECT 163.545 188.950 163.865 189.210 ;
        RECT 164.005 189.150 164.325 189.210 ;
        RECT 166.780 189.150 167.070 189.195 ;
        RECT 164.005 189.010 167.070 189.150 ;
        RECT 164.005 188.950 164.325 189.010 ;
        RECT 166.780 188.965 167.070 189.010 ;
        RECT 168.160 189.150 168.450 189.195 ;
        RECT 169.985 189.150 170.305 189.210 ;
        RECT 168.160 189.010 170.305 189.150 ;
        RECT 168.160 188.965 168.450 189.010 ;
        RECT 169.985 188.950 170.305 189.010 ;
        RECT 171.380 189.150 171.670 189.195 ;
        RECT 171.825 189.150 172.145 189.210 ;
        RECT 172.375 189.195 172.515 189.350 ;
        RECT 173.755 189.350 180.340 189.490 ;
        RECT 171.380 189.010 172.145 189.150 ;
        RECT 171.380 188.965 171.670 189.010 ;
        RECT 171.825 188.950 172.145 189.010 ;
        RECT 172.300 188.965 172.590 189.195 ;
        RECT 172.745 189.150 173.065 189.210 ;
        RECT 173.755 189.195 173.895 189.350 ;
        RECT 173.680 189.150 173.970 189.195 ;
        RECT 172.745 189.010 173.970 189.150 ;
        RECT 172.745 188.950 173.065 189.010 ;
        RECT 173.680 188.965 173.970 189.010 ;
        RECT 174.585 188.950 174.905 189.210 ;
        RECT 175.520 189.150 175.810 189.195 ;
        RECT 175.965 189.150 176.285 189.210 ;
        RECT 177.895 189.195 178.035 189.350 ;
        RECT 175.520 189.010 176.285 189.150 ;
        RECT 175.520 188.965 175.810 189.010 ;
        RECT 175.965 188.950 176.285 189.010 ;
        RECT 176.440 188.965 176.730 189.195 ;
        RECT 177.820 188.965 178.110 189.195 ;
        RECT 179.185 189.150 179.505 189.210 ;
        RECT 180.200 189.195 180.340 189.350 ;
        RECT 179.660 189.150 179.950 189.195 ;
        RECT 179.185 189.010 179.950 189.150 ;
        RECT 170.460 188.625 170.750 188.855 ;
        RECT 170.905 188.810 171.225 188.870 ;
        RECT 176.515 188.810 176.655 188.965 ;
        RECT 179.185 188.950 179.505 189.010 ;
        RECT 179.660 188.965 179.950 189.010 ;
        RECT 180.125 188.965 180.415 189.195 ;
        RECT 170.905 188.670 176.655 188.810 ;
        RECT 179.735 188.810 179.875 188.965 ;
        RECT 181.025 188.950 181.345 189.210 ;
        RECT 181.485 188.950 181.805 189.210 ;
        RECT 182.190 189.150 182.480 189.195 ;
        RECT 182.865 189.150 183.185 189.210 ;
        RECT 182.190 189.010 183.185 189.150 ;
        RECT 182.190 188.965 182.480 189.010 ;
        RECT 182.865 188.950 183.185 189.010 ;
        RECT 183.325 188.950 183.645 189.210 ;
        RECT 184.110 189.150 184.400 189.195 ;
        RECT 184.705 189.150 185.025 189.210 ;
        RECT 186.175 189.195 186.315 189.690 ;
        RECT 188.385 189.630 188.705 189.690 ;
        RECT 197.585 189.630 197.905 189.690 ;
        RECT 187.005 189.490 187.325 189.550 ;
        RECT 191.605 189.490 191.925 189.550 ;
        RECT 199.055 189.535 199.195 190.030 ;
        RECT 213.700 190.030 214.465 190.170 ;
        RECT 213.700 189.985 213.990 190.030 ;
        RECT 214.145 189.970 214.465 190.030 ;
        RECT 222.900 190.170 223.190 190.215 ;
        RECT 223.805 190.170 224.125 190.230 ;
        RECT 222.900 190.030 224.125 190.170 ;
        RECT 222.900 189.985 223.190 190.030 ;
        RECT 223.805 189.970 224.125 190.030 ;
        RECT 224.740 190.170 225.030 190.215 ;
        RECT 229.325 190.170 229.645 190.230 ;
        RECT 224.740 190.030 229.645 190.170 ;
        RECT 224.740 189.985 225.030 190.030 ;
        RECT 229.325 189.970 229.645 190.030 ;
        RECT 211.860 189.830 212.150 189.875 ;
        RECT 226.565 189.830 226.885 189.890 ;
        RECT 211.860 189.690 226.885 189.830 ;
        RECT 211.860 189.645 212.150 189.690 ;
        RECT 226.565 189.630 226.885 189.690 ;
        RECT 227.960 189.830 228.250 189.875 ;
        RECT 228.405 189.830 228.725 189.890 ;
        RECT 227.960 189.690 228.725 189.830 ;
        RECT 227.960 189.645 228.250 189.690 ;
        RECT 228.405 189.630 228.725 189.690 ;
        RECT 198.980 189.490 199.270 189.535 ;
        RECT 207.705 189.490 208.025 189.550 ;
        RECT 187.005 189.350 190.920 189.490 ;
        RECT 187.005 189.290 187.325 189.350 ;
        RECT 184.110 189.010 185.025 189.150 ;
        RECT 184.110 188.965 184.400 189.010 ;
        RECT 184.705 188.950 185.025 189.010 ;
        RECT 186.100 188.965 186.390 189.195 ;
        RECT 186.545 189.150 186.865 189.210 ;
        RECT 188.845 189.195 189.165 189.210 ;
        RECT 190.780 189.195 190.920 189.350 ;
        RECT 191.605 189.350 197.815 189.490 ;
        RECT 191.605 189.290 191.925 189.350 ;
        RECT 197.675 189.195 197.815 189.350 ;
        RECT 198.980 189.350 208.025 189.490 ;
        RECT 198.980 189.305 199.270 189.350 ;
        RECT 207.705 189.290 208.025 189.350 ;
        RECT 211.385 189.490 211.705 189.550 ;
        RECT 225.200 189.490 225.490 189.535 ;
        RECT 229.785 189.490 230.105 189.550 ;
        RECT 211.385 189.350 230.105 189.490 ;
        RECT 211.385 189.290 211.705 189.350 ;
        RECT 225.200 189.305 225.490 189.350 ;
        RECT 229.785 189.290 230.105 189.350 ;
        RECT 186.545 189.010 187.060 189.150 ;
        RECT 186.175 188.810 186.315 188.965 ;
        RECT 186.545 188.950 186.865 189.010 ;
        RECT 188.630 188.965 189.165 189.195 ;
        RECT 190.240 188.965 190.530 189.195 ;
        RECT 190.705 188.965 190.995 189.195 ;
        RECT 197.600 188.965 197.890 189.195 ;
        RECT 212.780 188.965 213.070 189.195 ;
        RECT 220.125 189.150 220.445 189.210 ;
        RECT 223.820 189.150 224.110 189.195 ;
        RECT 220.125 189.010 224.110 189.150 ;
        RECT 188.845 188.950 189.165 188.965 ;
        RECT 179.735 188.670 186.315 188.810 ;
        RECT 167.700 188.470 167.990 188.515 ;
        RECT 169.065 188.470 169.385 188.530 ;
        RECT 167.700 188.330 169.385 188.470 ;
        RECT 170.535 188.470 170.675 188.625 ;
        RECT 170.905 188.610 171.225 188.670 ;
        RECT 187.465 188.610 187.785 188.870 ;
        RECT 187.940 188.625 188.230 188.855 ;
        RECT 190.315 188.810 190.455 188.965 ;
        RECT 191.605 188.810 191.925 188.870 ;
        RECT 190.315 188.670 191.925 188.810 ;
        RECT 171.365 188.470 171.685 188.530 ;
        RECT 177.345 188.470 177.665 188.530 ;
        RECT 170.535 188.330 177.665 188.470 ;
        RECT 167.700 188.285 167.990 188.330 ;
        RECT 169.065 188.270 169.385 188.330 ;
        RECT 171.365 188.270 171.685 188.330 ;
        RECT 177.345 188.270 177.665 188.330 ;
        RECT 181.025 188.470 181.345 188.530 ;
        RECT 183.785 188.470 184.105 188.530 ;
        RECT 181.025 188.330 184.105 188.470 ;
        RECT 181.025 188.270 181.345 188.330 ;
        RECT 183.785 188.270 184.105 188.330 ;
        RECT 185.180 188.470 185.470 188.515 ;
        RECT 188.015 188.470 188.155 188.625 ;
        RECT 191.605 188.610 191.925 188.670 ;
        RECT 192.080 188.810 192.370 188.855 ;
        RECT 197.125 188.810 197.445 188.870 ;
        RECT 192.080 188.670 197.445 188.810 ;
        RECT 192.080 188.625 192.370 188.670 ;
        RECT 197.125 188.610 197.445 188.670 ;
        RECT 208.165 188.810 208.485 188.870 ;
        RECT 212.855 188.810 212.995 188.965 ;
        RECT 220.125 188.950 220.445 189.010 ;
        RECT 223.820 188.965 224.110 189.010 ;
        RECT 225.645 189.150 225.965 189.210 ;
        RECT 227.040 189.150 227.330 189.195 ;
        RECT 225.645 189.010 227.330 189.150 ;
        RECT 225.645 188.950 225.965 189.010 ;
        RECT 227.040 188.965 227.330 189.010 ;
        RECT 229.340 188.965 229.630 189.195 ;
        RECT 208.165 188.670 212.995 188.810 ;
        RECT 226.105 188.810 226.425 188.870 ;
        RECT 229.415 188.810 229.555 188.965 ;
        RECT 230.705 188.950 231.025 189.210 ;
        RECT 226.105 188.670 229.555 188.810 ;
        RECT 208.165 188.610 208.485 188.670 ;
        RECT 226.105 188.610 226.425 188.670 ;
        RECT 185.180 188.330 188.155 188.470 ;
        RECT 195.760 188.470 196.050 188.515 ;
        RECT 196.665 188.470 196.985 188.530 ;
        RECT 195.760 188.330 196.985 188.470 ;
        RECT 185.180 188.285 185.470 188.330 ;
        RECT 195.760 188.285 196.050 188.330 ;
        RECT 196.665 188.270 196.985 188.330 ;
        RECT 198.045 188.270 198.365 188.530 ;
        RECT 222.885 188.470 223.205 188.530 ;
        RECT 228.420 188.470 228.710 188.515 ;
        RECT 222.885 188.330 228.710 188.470 ;
        RECT 222.885 188.270 223.205 188.330 ;
        RECT 228.420 188.285 228.710 188.330 ;
        RECT 228.865 188.470 229.185 188.530 ;
        RECT 229.800 188.470 230.090 188.515 ;
        RECT 228.865 188.330 230.090 188.470 ;
        RECT 228.865 188.270 229.185 188.330 ;
        RECT 229.800 188.285 230.090 188.330 ;
        RECT 149.905 185.540 150.865 185.770 ;
        RECT 151.195 185.540 152.155 185.770 ;
        RECT 152.845 185.165 155.165 187.965 ;
        RECT 162.095 187.650 236.155 188.130 ;
        RECT 165.860 187.265 166.150 187.495 ;
        RECT 167.225 187.450 167.545 187.510 ;
        RECT 167.700 187.450 167.990 187.495 ;
        RECT 173.205 187.450 173.525 187.510 ;
        RECT 167.225 187.310 167.990 187.450 ;
        RECT 165.935 187.110 166.075 187.265 ;
        RECT 167.225 187.250 167.545 187.310 ;
        RECT 167.700 187.265 167.990 187.310 ;
        RECT 170.075 187.310 173.525 187.450 ;
        RECT 169.525 187.110 169.845 187.170 ;
        RECT 165.935 186.970 169.845 187.110 ;
        RECT 169.525 186.910 169.845 186.970 ;
        RECT 163.085 186.770 163.405 186.830 ;
        RECT 163.560 186.770 163.850 186.815 ;
        RECT 163.085 186.630 163.850 186.770 ;
        RECT 163.085 186.570 163.405 186.630 ;
        RECT 163.560 186.585 163.850 186.630 ;
        RECT 164.940 186.770 165.230 186.815 ;
        RECT 165.385 186.770 165.705 186.830 ;
        RECT 164.940 186.630 165.705 186.770 ;
        RECT 164.940 186.585 165.230 186.630 ;
        RECT 165.385 186.570 165.705 186.630 ;
        RECT 166.320 186.585 166.610 186.815 ;
        RECT 166.765 186.770 167.085 186.830 ;
        RECT 170.075 186.815 170.215 187.310 ;
        RECT 173.205 187.250 173.525 187.310 ;
        RECT 175.060 187.450 175.350 187.495 ;
        RECT 175.505 187.450 175.825 187.510 ;
        RECT 175.060 187.310 175.825 187.450 ;
        RECT 175.060 187.265 175.350 187.310 ;
        RECT 175.505 187.250 175.825 187.310 ;
        RECT 180.565 187.250 180.885 187.510 ;
        RECT 181.960 187.450 182.250 187.495 ;
        RECT 183.325 187.450 183.645 187.510 ;
        RECT 181.960 187.310 183.645 187.450 ;
        RECT 181.960 187.265 182.250 187.310 ;
        RECT 183.325 187.250 183.645 187.310 ;
        RECT 186.545 187.250 186.865 187.510 ;
        RECT 187.480 187.450 187.770 187.495 ;
        RECT 190.685 187.450 191.005 187.510 ;
        RECT 187.480 187.310 191.005 187.450 ;
        RECT 187.480 187.265 187.770 187.310 ;
        RECT 190.685 187.250 191.005 187.310 ;
        RECT 191.260 187.310 195.975 187.450 ;
        RECT 170.905 187.110 171.225 187.170 ;
        RECT 170.535 186.970 171.225 187.110 ;
        RECT 170.535 186.815 170.675 186.970 ;
        RECT 170.905 186.910 171.225 186.970 ;
        RECT 168.620 186.770 168.910 186.815 ;
        RECT 166.765 186.630 168.910 186.770 ;
        RECT 166.395 186.430 166.535 186.585 ;
        RECT 166.765 186.570 167.085 186.630 ;
        RECT 168.620 186.585 168.910 186.630 ;
        RECT 170.000 186.585 170.290 186.815 ;
        RECT 170.460 186.585 170.750 186.815 ;
        RECT 171.380 186.585 171.670 186.815 ;
        RECT 169.525 186.430 169.845 186.490 ;
        RECT 166.395 186.290 169.845 186.430 ;
        RECT 169.525 186.230 169.845 186.290 ;
        RECT 164.480 186.090 164.770 186.135 ;
        RECT 171.455 186.090 171.595 186.585 ;
        RECT 172.745 186.570 173.065 186.830 ;
        RECT 164.480 185.950 171.595 186.090 ;
        RECT 173.295 186.090 173.435 187.250 ;
        RECT 173.680 187.110 173.970 187.155 ;
        RECT 186.635 187.110 186.775 187.250 ;
        RECT 189.305 187.110 189.625 187.170 ;
        RECT 191.260 187.110 191.400 187.310 ;
        RECT 173.680 186.970 182.175 187.110 ;
        RECT 186.635 186.970 191.400 187.110 ;
        RECT 191.620 187.110 191.910 187.155 ;
        RECT 193.445 187.110 193.765 187.170 ;
        RECT 191.620 186.970 193.765 187.110 ;
        RECT 173.680 186.925 173.970 186.970 ;
        RECT 182.035 186.830 182.175 186.970 ;
        RECT 189.305 186.910 189.625 186.970 ;
        RECT 174.585 186.770 174.905 186.830 ;
        RECT 175.980 186.770 176.270 186.815 ;
        RECT 174.585 186.630 176.270 186.770 ;
        RECT 174.585 186.570 174.905 186.630 ;
        RECT 175.980 186.585 176.270 186.630 ;
        RECT 176.885 186.570 177.205 186.830 ;
        RECT 177.360 186.770 177.650 186.815 ;
        RECT 177.805 186.770 178.125 186.830 ;
        RECT 177.360 186.630 178.125 186.770 ;
        RECT 177.360 186.585 177.650 186.630 ;
        RECT 177.805 186.570 178.125 186.630 ;
        RECT 178.740 186.585 179.030 186.815 ;
        RECT 179.205 186.585 179.495 186.815 ;
        RECT 180.105 186.770 180.425 186.830 ;
        RECT 181.040 186.770 181.330 186.815 ;
        RECT 180.105 186.630 181.330 186.770 ;
        RECT 174.125 186.430 174.445 186.490 ;
        RECT 178.815 186.430 178.955 186.585 ;
        RECT 174.125 186.290 178.955 186.430 ;
        RECT 174.125 186.230 174.445 186.290 ;
        RECT 177.805 186.090 178.125 186.150 ;
        RECT 173.295 185.950 178.125 186.090 ;
        RECT 164.480 185.905 164.770 185.950 ;
        RECT 177.805 185.890 178.125 185.950 ;
        RECT 167.240 185.750 167.530 185.795 ;
        RECT 168.145 185.750 168.465 185.810 ;
        RECT 167.240 185.610 168.465 185.750 ;
        RECT 167.240 185.565 167.530 185.610 ;
        RECT 168.145 185.550 168.465 185.610 ;
        RECT 169.540 185.750 169.830 185.795 ;
        RECT 171.825 185.750 172.145 185.810 ;
        RECT 169.540 185.610 172.145 185.750 ;
        RECT 169.540 185.565 169.830 185.610 ;
        RECT 171.825 185.550 172.145 185.610 ;
        RECT 175.965 185.750 176.285 185.810 ;
        RECT 179.275 185.750 179.415 186.585 ;
        RECT 180.105 186.570 180.425 186.630 ;
        RECT 181.040 186.585 181.330 186.630 ;
        RECT 181.945 186.570 182.265 186.830 ;
        RECT 182.420 186.770 182.710 186.815 ;
        RECT 182.865 186.770 183.185 186.830 ;
        RECT 182.420 186.630 183.185 186.770 ;
        RECT 182.420 186.585 182.710 186.630 ;
        RECT 182.865 186.570 183.185 186.630 ;
        RECT 183.800 186.770 184.090 186.815 ;
        RECT 186.085 186.770 186.405 186.830 ;
        RECT 183.800 186.630 186.405 186.770 ;
        RECT 183.800 186.585 184.090 186.630 ;
        RECT 181.485 186.430 181.805 186.490 ;
        RECT 183.875 186.430 184.015 186.585 ;
        RECT 186.085 186.570 186.405 186.630 ;
        RECT 186.560 186.770 186.850 186.815 ;
        RECT 188.385 186.770 188.705 186.830 ;
        RECT 186.560 186.630 188.705 186.770 ;
        RECT 186.560 186.585 186.850 186.630 ;
        RECT 188.385 186.570 188.705 186.630 ;
        RECT 188.860 186.770 189.150 186.815 ;
        RECT 189.765 186.770 190.085 186.830 ;
        RECT 190.780 186.815 190.920 186.970 ;
        RECT 191.620 186.925 191.910 186.970 ;
        RECT 193.445 186.910 193.765 186.970 ;
        RECT 188.860 186.630 190.085 186.770 ;
        RECT 188.860 186.585 189.150 186.630 ;
        RECT 189.765 186.570 190.085 186.630 ;
        RECT 190.240 186.585 190.530 186.815 ;
        RECT 190.705 186.585 190.995 186.815 ;
        RECT 190.315 186.430 190.455 186.585 ;
        RECT 192.065 186.570 192.385 186.830 ;
        RECT 192.525 186.815 192.845 186.830 ;
        RECT 192.525 186.585 192.855 186.815 ;
        RECT 192.525 186.570 192.845 186.585 ;
        RECT 194.825 186.570 195.145 186.830 ;
        RECT 195.285 186.570 195.605 186.830 ;
        RECT 195.835 186.815 195.975 187.310 ;
        RECT 198.505 187.250 198.825 187.510 ;
        RECT 208.165 187.250 208.485 187.510 ;
        RECT 209.085 187.450 209.405 187.510 ;
        RECT 218.300 187.450 218.590 187.495 ;
        RECT 209.085 187.310 218.590 187.450 ;
        RECT 209.085 187.250 209.405 187.310 ;
        RECT 218.300 187.265 218.590 187.310 ;
        RECT 221.965 187.450 222.285 187.510 ;
        RECT 221.965 187.310 228.635 187.450 ;
        RECT 221.965 187.250 222.285 187.310 ;
        RECT 196.665 186.910 196.985 187.170 ;
        RECT 197.125 186.910 197.445 187.170 ;
        RECT 208.255 187.110 208.395 187.250 ;
        RECT 200.435 186.970 208.395 187.110 ;
        RECT 221.525 187.110 221.815 187.155 ;
        RECT 227.045 187.110 227.335 187.155 ;
        RECT 227.965 187.110 228.255 187.155 ;
        RECT 221.525 186.970 228.255 187.110 ;
        RECT 228.495 187.110 228.635 187.310 ;
        RECT 229.325 187.250 229.645 187.510 ;
        RECT 232.100 187.450 232.390 187.495 ;
        RECT 233.005 187.450 233.325 187.510 ;
        RECT 232.100 187.310 233.325 187.450 ;
        RECT 232.100 187.265 232.390 187.310 ;
        RECT 233.005 187.250 233.325 187.310 ;
        RECT 228.495 186.970 232.775 187.110 ;
        RECT 197.585 186.815 197.905 186.830 ;
        RECT 195.765 186.585 196.055 186.815 ;
        RECT 197.585 186.770 197.915 186.815 ;
        RECT 197.585 186.630 198.100 186.770 ;
        RECT 197.585 186.585 197.915 186.630 ;
        RECT 199.900 186.585 200.190 186.815 ;
        RECT 197.585 186.570 197.905 186.585 ;
        RECT 194.365 186.430 194.685 186.490 ;
        RECT 181.485 186.290 184.015 186.430 ;
        RECT 188.935 186.290 190.455 186.430 ;
        RECT 193.995 186.290 194.685 186.430 ;
        RECT 181.485 186.230 181.805 186.290 ;
        RECT 188.935 186.150 189.075 186.290 ;
        RECT 188.845 185.890 189.165 186.150 ;
        RECT 193.995 186.135 194.135 186.290 ;
        RECT 194.365 186.230 194.685 186.290 ;
        RECT 196.665 186.430 196.985 186.490 ;
        RECT 199.975 186.430 200.115 186.585 ;
        RECT 196.665 186.290 200.115 186.430 ;
        RECT 196.665 186.230 196.985 186.290 ;
        RECT 193.920 185.905 194.210 186.135 ;
        RECT 195.745 186.090 196.065 186.150 ;
        RECT 200.435 186.090 200.575 186.970 ;
        RECT 221.525 186.925 221.815 186.970 ;
        RECT 227.045 186.925 227.335 186.970 ;
        RECT 227.965 186.925 228.255 186.970 ;
        RECT 206.785 186.770 207.105 186.830 ;
        RECT 208.180 186.770 208.470 186.815 ;
        RECT 206.785 186.630 208.470 186.770 ;
        RECT 206.785 186.570 207.105 186.630 ;
        RECT 208.180 186.585 208.470 186.630 ;
        RECT 208.625 186.690 208.945 186.830 ;
        RECT 210.925 186.770 211.245 186.830 ;
        RECT 211.400 186.770 211.690 186.815 ;
        RECT 209.560 186.690 209.850 186.735 ;
        RECT 208.625 186.570 209.850 186.690 ;
        RECT 208.805 186.550 209.850 186.570 ;
        RECT 209.560 186.505 209.850 186.550 ;
        RECT 210.020 186.690 210.310 186.735 ;
        RECT 210.020 186.550 210.695 186.690 ;
        RECT 210.925 186.630 211.690 186.770 ;
        RECT 210.925 186.570 211.245 186.630 ;
        RECT 211.400 186.585 211.690 186.630 ;
        RECT 211.845 186.770 212.165 186.830 ;
        RECT 214.160 186.770 214.450 186.815 ;
        RECT 211.845 186.630 214.450 186.770 ;
        RECT 211.845 186.570 212.165 186.630 ;
        RECT 214.160 186.585 214.450 186.630 ;
        RECT 215.540 186.585 215.830 186.815 ;
        RECT 216.445 186.770 216.765 186.830 ;
        RECT 217.840 186.770 218.130 186.815 ;
        RECT 216.445 186.630 218.130 186.770 ;
        RECT 210.020 186.505 210.310 186.550 ;
        RECT 210.555 186.150 210.695 186.550 ;
        RECT 212.765 186.430 213.085 186.490 ;
        RECT 215.615 186.430 215.755 186.585 ;
        RECT 216.445 186.570 216.765 186.630 ;
        RECT 217.840 186.585 218.130 186.630 ;
        RECT 219.220 186.585 219.510 186.815 ;
        RECT 219.665 186.770 219.985 186.830 ;
        RECT 221.060 186.770 221.350 186.815 ;
        RECT 219.665 186.630 221.350 186.770 ;
        RECT 212.765 186.290 215.755 186.430 ;
        RECT 216.905 186.430 217.225 186.490 ;
        RECT 219.295 186.430 219.435 186.585 ;
        RECT 219.665 186.570 219.985 186.630 ;
        RECT 221.060 186.585 221.350 186.630 ;
        RECT 222.445 186.770 222.735 186.815 ;
        RECT 224.285 186.770 224.575 186.815 ;
        RECT 222.445 186.630 224.575 186.770 ;
        RECT 222.445 186.585 222.735 186.630 ;
        RECT 224.285 186.585 224.575 186.630 ;
        RECT 226.630 186.770 226.920 186.815 ;
        RECT 228.470 186.770 228.760 186.815 ;
        RECT 226.630 186.630 228.760 186.770 ;
        RECT 226.630 186.585 226.920 186.630 ;
        RECT 228.470 186.585 228.760 186.630 ;
        RECT 229.785 186.570 230.105 186.830 ;
        RECT 231.165 186.570 231.485 186.830 ;
        RECT 225.645 186.475 225.965 186.490 ;
        RECT 216.905 186.290 219.435 186.430 ;
        RECT 212.765 186.230 213.085 186.290 ;
        RECT 216.905 186.230 217.225 186.290 ;
        RECT 220.140 186.245 220.430 186.475 ;
        RECT 224.740 186.430 225.030 186.475 ;
        RECT 223.895 186.290 225.030 186.430 ;
        RECT 195.745 185.950 200.575 186.090 ;
        RECT 204.945 186.090 205.265 186.150 ;
        RECT 207.705 186.090 208.025 186.150 ;
        RECT 204.945 185.950 208.025 186.090 ;
        RECT 195.745 185.890 196.065 185.950 ;
        RECT 204.945 185.890 205.265 185.950 ;
        RECT 207.705 185.890 208.025 185.950 ;
        RECT 210.465 185.890 210.785 186.150 ;
        RECT 210.940 186.090 211.230 186.135 ;
        RECT 214.145 186.090 214.465 186.150 ;
        RECT 210.940 185.950 214.465 186.090 ;
        RECT 210.940 185.905 211.230 185.950 ;
        RECT 214.145 185.890 214.465 185.950 ;
        RECT 216.460 186.090 216.750 186.135 ;
        RECT 220.215 186.090 220.355 186.245 ;
        RECT 216.460 185.950 220.355 186.090 ;
        RECT 221.045 186.090 221.365 186.150 ;
        RECT 223.360 186.090 223.650 186.135 ;
        RECT 221.045 185.950 223.650 186.090 ;
        RECT 216.460 185.905 216.750 185.950 ;
        RECT 221.045 185.890 221.365 185.950 ;
        RECT 223.360 185.905 223.650 185.950 ;
        RECT 175.965 185.610 179.415 185.750 ;
        RECT 175.965 185.550 176.285 185.610 ;
        RECT 183.325 185.550 183.645 185.810 ;
        RECT 184.705 185.750 185.025 185.810 ;
        RECT 186.545 185.750 186.865 185.810 ;
        RECT 184.705 185.610 186.865 185.750 ;
        RECT 184.705 185.550 185.025 185.610 ;
        RECT 186.545 185.550 186.865 185.610 ;
        RECT 189.780 185.750 190.070 185.795 ;
        RECT 191.605 185.750 191.925 185.810 ;
        RECT 189.780 185.610 191.925 185.750 ;
        RECT 189.780 185.565 190.070 185.610 ;
        RECT 191.605 185.550 191.925 185.610 ;
        RECT 193.460 185.750 193.750 185.795 ;
        RECT 197.585 185.750 197.905 185.810 ;
        RECT 193.460 185.610 197.905 185.750 ;
        RECT 193.460 185.565 193.750 185.610 ;
        RECT 197.585 185.550 197.905 185.610 ;
        RECT 198.505 185.750 198.825 185.810 ;
        RECT 198.980 185.750 199.270 185.795 ;
        RECT 198.505 185.610 199.270 185.750 ;
        RECT 198.505 185.550 198.825 185.610 ;
        RECT 198.980 185.565 199.270 185.610 ;
        RECT 204.025 185.750 204.345 185.810 ;
        RECT 207.260 185.750 207.550 185.795 ;
        RECT 204.025 185.610 207.550 185.750 ;
        RECT 204.025 185.550 204.345 185.610 ;
        RECT 207.260 185.565 207.550 185.610 ;
        RECT 208.165 185.750 208.485 185.810 ;
        RECT 208.640 185.750 208.930 185.795 ;
        RECT 208.165 185.610 208.930 185.750 ;
        RECT 208.165 185.550 208.485 185.610 ;
        RECT 208.640 185.565 208.930 185.610 ;
        RECT 212.320 185.750 212.610 185.795 ;
        RECT 213.225 185.750 213.545 185.810 ;
        RECT 212.320 185.610 213.545 185.750 ;
        RECT 212.320 185.565 212.610 185.610 ;
        RECT 213.225 185.550 213.545 185.610 ;
        RECT 215.065 185.550 215.385 185.810 ;
        RECT 215.525 185.750 215.845 185.810 ;
        RECT 216.920 185.750 217.210 185.795 ;
        RECT 215.525 185.610 217.210 185.750 ;
        RECT 223.895 185.750 224.035 186.290 ;
        RECT 224.740 186.245 225.030 186.290 ;
        RECT 225.430 186.245 225.965 186.475 ;
        RECT 226.120 186.430 226.410 186.475 ;
        RECT 227.025 186.430 227.345 186.490 ;
        RECT 226.120 186.290 227.345 186.430 ;
        RECT 226.120 186.245 226.410 186.290 ;
        RECT 225.645 186.230 225.965 186.245 ;
        RECT 227.025 186.230 227.345 186.290 ;
        RECT 227.945 186.430 228.265 186.490 ;
        RECT 227.945 186.290 230.935 186.430 ;
        RECT 227.945 186.230 228.265 186.290 ;
        RECT 224.320 186.090 224.610 186.135 ;
        RECT 227.550 186.090 227.840 186.135 ;
        RECT 224.320 185.950 227.840 186.090 ;
        RECT 224.320 185.905 224.610 185.950 ;
        RECT 227.550 185.905 227.840 185.950 ;
        RECT 228.865 185.750 229.185 185.810 ;
        RECT 223.895 185.610 229.185 185.750 ;
        RECT 215.525 185.550 215.845 185.610 ;
        RECT 216.920 185.565 217.210 185.610 ;
        RECT 228.865 185.550 229.185 185.610 ;
        RECT 230.245 185.550 230.565 185.810 ;
        RECT 230.795 185.750 230.935 186.290 ;
        RECT 232.635 186.135 232.775 186.970 ;
        RECT 233.480 186.585 233.770 186.815 ;
        RECT 232.560 185.905 232.850 186.135 ;
        RECT 233.555 185.750 233.695 186.585 ;
        RECT 230.795 185.610 233.695 185.750 ;
        RECT 108.515 184.765 155.165 185.165 ;
        RECT 162.095 184.930 236.155 185.410 ;
        RECT 166.765 184.530 167.085 184.790 ;
        RECT 169.525 184.730 169.845 184.790 ;
        RECT 169.525 184.590 173.205 184.730 ;
        RECT 169.525 184.530 169.845 184.590 ;
        RECT 167.225 184.390 167.545 184.450 ;
        RECT 169.985 184.390 170.305 184.450 ;
        RECT 167.225 184.250 170.305 184.390 ;
        RECT 173.065 184.390 173.205 184.590 ;
        RECT 174.585 184.530 174.905 184.790 ;
        RECT 178.265 184.730 178.585 184.790 ;
        RECT 181.485 184.730 181.805 184.790 ;
        RECT 178.265 184.590 181.805 184.730 ;
        RECT 178.265 184.530 178.585 184.590 ;
        RECT 181.485 184.530 181.805 184.590 ;
        RECT 182.405 184.730 182.725 184.790 ;
        RECT 185.625 184.730 185.945 184.790 ;
        RECT 182.405 184.590 185.945 184.730 ;
        RECT 182.405 184.530 182.725 184.590 ;
        RECT 185.625 184.530 185.945 184.590 ;
        RECT 186.100 184.730 186.390 184.775 ;
        RECT 197.585 184.730 197.905 184.790 ;
        RECT 186.100 184.590 196.895 184.730 ;
        RECT 186.100 184.545 186.390 184.590 ;
        RECT 175.045 184.390 175.365 184.450 ;
        RECT 173.065 184.250 175.365 184.390 ;
        RECT 167.225 184.190 167.545 184.250 ;
        RECT 169.985 184.190 170.305 184.250 ;
        RECT 175.045 184.190 175.365 184.250 ;
        RECT 180.580 184.390 180.870 184.435 ;
        RECT 187.925 184.390 188.245 184.450 ;
        RECT 180.580 184.250 188.245 184.390 ;
        RECT 180.580 184.205 180.870 184.250 ;
        RECT 187.925 184.190 188.245 184.250 ;
        RECT 191.605 184.390 191.925 184.450 ;
        RECT 194.825 184.390 195.145 184.450 ;
        RECT 191.605 184.250 195.145 184.390 ;
        RECT 191.605 184.190 191.925 184.250 ;
        RECT 194.825 184.190 195.145 184.250 ;
        RECT 195.745 184.190 196.065 184.450 ;
        RECT 196.220 184.205 196.510 184.435 ;
        RECT 168.145 184.050 168.465 184.110 ;
        RECT 181.025 184.050 181.345 184.110 ;
        RECT 168.145 183.910 176.655 184.050 ;
        RECT 168.145 183.850 168.465 183.910 ;
        RECT 164.020 183.710 164.310 183.755 ;
        RECT 164.465 183.710 164.785 183.770 ;
        RECT 164.020 183.570 164.785 183.710 ;
        RECT 164.020 183.525 164.310 183.570 ;
        RECT 164.465 183.510 164.785 183.570 ;
        RECT 165.400 183.710 165.690 183.755 ;
        RECT 166.765 183.710 167.085 183.770 ;
        RECT 167.685 183.755 168.005 183.770 ;
        RECT 165.400 183.570 167.085 183.710 ;
        RECT 165.400 183.525 165.690 183.570 ;
        RECT 166.765 183.510 167.085 183.570 ;
        RECT 167.675 183.525 168.005 183.755 ;
        RECT 169.525 183.710 169.845 183.770 ;
        RECT 169.330 183.570 169.845 183.710 ;
        RECT 167.685 183.510 168.005 183.525 ;
        RECT 169.525 183.510 169.845 183.570 ;
        RECT 169.985 183.710 170.305 183.770 ;
        RECT 171.380 183.710 171.670 183.755 ;
        RECT 169.985 183.570 171.670 183.710 ;
        RECT 169.985 183.510 170.305 183.570 ;
        RECT 171.380 183.525 171.670 183.570 ;
        RECT 171.845 183.525 172.135 183.755 ;
        RECT 166.395 183.230 167.915 183.370 ;
        RECT 164.925 182.830 165.245 183.090 ;
        RECT 166.395 183.075 166.535 183.230 ;
        RECT 166.320 182.845 166.610 183.075 ;
        RECT 167.775 183.030 167.915 183.230 ;
        RECT 168.145 183.170 168.465 183.430 ;
        RECT 168.620 183.370 168.910 183.415 ;
        RECT 170.905 183.370 171.225 183.430 ;
        RECT 168.620 183.230 171.225 183.370 ;
        RECT 171.920 183.370 172.060 183.525 ;
        RECT 172.745 183.510 173.065 183.770 ;
        RECT 173.205 183.510 173.525 183.770 ;
        RECT 173.665 183.755 173.985 183.770 ;
        RECT 173.665 183.710 173.995 183.755 ;
        RECT 173.665 183.570 174.180 183.710 ;
        RECT 173.665 183.525 173.995 183.570 ;
        RECT 173.665 183.510 173.985 183.525 ;
        RECT 175.505 183.510 175.825 183.770 ;
        RECT 176.515 183.755 176.655 183.910 ;
        RECT 178.355 183.910 181.345 184.050 ;
        RECT 176.440 183.525 176.730 183.755 ;
        RECT 177.820 183.525 178.110 183.755 ;
        RECT 172.285 183.370 172.605 183.430 ;
        RECT 177.895 183.370 178.035 183.525 ;
        RECT 171.920 183.230 178.035 183.370 ;
        RECT 168.620 183.185 168.910 183.230 ;
        RECT 170.905 183.170 171.225 183.230 ;
        RECT 172.285 183.170 172.605 183.230 ;
        RECT 176.425 183.030 176.745 183.090 ;
        RECT 167.775 182.890 176.745 183.030 ;
        RECT 176.425 182.830 176.745 182.890 ;
        RECT 177.805 183.030 178.125 183.090 ;
        RECT 178.355 183.030 178.495 183.910 ;
        RECT 181.025 183.850 181.345 183.910 ;
        RECT 183.325 184.050 183.645 184.110 ;
        RECT 196.295 184.050 196.435 184.205 ;
        RECT 183.325 183.910 186.775 184.050 ;
        RECT 183.325 183.850 183.645 183.910 ;
        RECT 179.645 183.510 179.965 183.770 ;
        RECT 181.960 183.525 182.250 183.755 ;
        RECT 178.740 183.370 179.030 183.415 ;
        RECT 181.485 183.370 181.805 183.430 ;
        RECT 178.740 183.230 181.805 183.370 ;
        RECT 182.035 183.370 182.175 183.525 ;
        RECT 182.405 183.510 182.725 183.770 ;
        RECT 183.800 183.710 184.090 183.755 ;
        RECT 183.800 183.570 184.935 183.710 ;
        RECT 183.800 183.525 184.090 183.570 ;
        RECT 184.245 183.370 184.565 183.430 ;
        RECT 182.035 183.230 184.565 183.370 ;
        RECT 184.795 183.370 184.935 183.570 ;
        RECT 185.165 183.510 185.485 183.770 ;
        RECT 186.635 183.755 186.775 183.910 ;
        RECT 189.400 183.910 193.220 184.050 ;
        RECT 189.400 183.770 189.540 183.910 ;
        RECT 186.560 183.525 186.850 183.755 ;
        RECT 187.005 183.710 187.325 183.770 ;
        RECT 187.005 183.570 187.520 183.710 ;
        RECT 187.005 183.510 187.325 183.570 ;
        RECT 188.845 183.510 189.165 183.770 ;
        RECT 189.305 183.710 189.625 183.770 ;
        RECT 191.605 183.755 191.925 183.770 ;
        RECT 189.305 183.570 189.820 183.710 ;
        RECT 189.305 183.510 189.625 183.570 ;
        RECT 191.390 183.525 191.925 183.755 ;
        RECT 191.605 183.510 191.925 183.525 ;
        RECT 192.525 183.510 192.845 183.770 ;
        RECT 193.080 183.755 193.220 183.910 ;
        RECT 193.995 183.910 196.435 184.050 ;
        RECT 193.995 183.755 194.135 183.910 ;
        RECT 195.285 183.755 195.605 183.770 ;
        RECT 193.005 183.525 193.295 183.755 ;
        RECT 193.920 183.525 194.210 183.755 ;
        RECT 195.070 183.525 195.605 183.755 ;
        RECT 196.755 183.710 196.895 184.590 ;
        RECT 197.585 184.590 213.455 184.730 ;
        RECT 197.585 184.530 197.905 184.590 ;
        RECT 197.125 184.390 197.445 184.450 ;
        RECT 206.325 184.390 206.645 184.450 ;
        RECT 207.245 184.390 207.565 184.450 ;
        RECT 208.640 184.390 208.930 184.435 ;
        RECT 197.125 184.250 203.795 184.390 ;
        RECT 197.125 184.190 197.445 184.250 ;
        RECT 198.505 183.850 198.825 184.110 ;
        RECT 199.425 184.050 199.745 184.110 ;
        RECT 199.425 183.910 203.335 184.050 ;
        RECT 199.425 183.850 199.745 183.910 ;
        RECT 198.060 183.710 198.350 183.755 ;
        RECT 196.755 183.570 198.350 183.710 ;
        RECT 198.060 183.525 198.350 183.570 ;
        RECT 202.200 183.525 202.490 183.755 ;
        RECT 195.285 183.510 195.605 183.525 ;
        RECT 184.795 183.230 187.235 183.370 ;
        RECT 178.740 183.185 179.030 183.230 ;
        RECT 181.485 183.170 181.805 183.230 ;
        RECT 184.245 183.170 184.565 183.230 ;
        RECT 187.095 183.090 187.235 183.230 ;
        RECT 190.225 183.170 190.545 183.430 ;
        RECT 190.685 183.170 191.005 183.430 ;
        RECT 194.380 183.370 194.670 183.415 ;
        RECT 197.125 183.370 197.445 183.430 ;
        RECT 191.695 183.230 194.670 183.370 ;
        RECT 177.805 182.890 178.495 183.030 ;
        RECT 177.805 182.830 178.125 182.890 ;
        RECT 181.025 182.830 181.345 183.090 ;
        RECT 183.325 182.830 183.645 183.090 ;
        RECT 184.705 182.830 185.025 183.090 ;
        RECT 187.005 182.830 187.325 183.090 ;
        RECT 188.400 183.030 188.690 183.075 ;
        RECT 191.695 183.030 191.835 183.230 ;
        RECT 194.380 183.185 194.670 183.230 ;
        RECT 195.375 183.230 197.445 183.370 ;
        RECT 195.375 183.090 195.515 183.230 ;
        RECT 197.125 183.170 197.445 183.230 ;
        RECT 197.585 183.370 197.905 183.430 ;
        RECT 202.275 183.370 202.415 183.525 ;
        RECT 197.585 183.230 202.415 183.370 ;
        RECT 197.585 183.170 197.905 183.230 ;
        RECT 188.400 182.890 191.835 183.030 ;
        RECT 192.080 183.030 192.370 183.075 ;
        RECT 192.525 183.030 192.845 183.090 ;
        RECT 192.080 182.890 192.845 183.030 ;
        RECT 188.400 182.845 188.690 182.890 ;
        RECT 192.080 182.845 192.370 182.890 ;
        RECT 192.525 182.830 192.845 182.890 ;
        RECT 195.285 182.830 195.605 183.090 ;
        RECT 196.205 183.030 196.525 183.090 ;
        RECT 201.280 183.030 201.570 183.075 ;
        RECT 196.205 182.890 201.570 183.030 ;
        RECT 196.205 182.830 196.525 182.890 ;
        RECT 201.280 182.845 201.570 182.890 ;
        RECT 201.725 183.030 202.045 183.090 ;
        RECT 202.660 183.030 202.950 183.075 ;
        RECT 201.725 182.890 202.950 183.030 ;
        RECT 203.195 183.030 203.335 183.910 ;
        RECT 203.655 183.755 203.795 184.250 ;
        RECT 206.325 184.250 208.930 184.390 ;
        RECT 206.325 184.190 206.645 184.250 ;
        RECT 207.245 184.190 207.565 184.250 ;
        RECT 208.640 184.205 208.930 184.250 ;
        RECT 209.600 184.390 209.890 184.435 ;
        RECT 212.830 184.390 213.120 184.435 ;
        RECT 209.600 184.250 213.120 184.390 ;
        RECT 213.315 184.390 213.455 184.590 ;
        RECT 214.605 184.530 214.925 184.790 ;
        RECT 216.445 184.730 216.765 184.790 ;
        RECT 217.365 184.730 217.685 184.790 ;
        RECT 216.445 184.590 217.685 184.730 ;
        RECT 216.445 184.530 216.765 184.590 ;
        RECT 217.365 184.530 217.685 184.590 ;
        RECT 217.825 184.730 218.145 184.790 ;
        RECT 219.665 184.730 219.985 184.790 ;
        RECT 217.825 184.590 219.985 184.730 ;
        RECT 217.825 184.530 218.145 184.590 ;
        RECT 219.665 184.530 219.985 184.590 ;
        RECT 220.125 184.530 220.445 184.790 ;
        RECT 225.645 184.730 225.965 184.790 ;
        RECT 227.040 184.730 227.330 184.775 ;
        RECT 230.245 184.730 230.565 184.790 ;
        RECT 220.675 184.590 224.955 184.730 ;
        RECT 220.215 184.390 220.355 184.530 ;
        RECT 213.315 184.250 220.355 184.390 ;
        RECT 209.600 184.205 209.890 184.250 ;
        RECT 212.830 184.205 213.120 184.250 ;
        RECT 205.420 184.050 205.710 184.095 ;
        RECT 208.165 184.050 208.485 184.110 ;
        RECT 205.420 183.910 208.485 184.050 ;
        RECT 205.420 183.865 205.710 183.910 ;
        RECT 208.165 183.850 208.485 183.910 ;
        RECT 210.020 184.050 210.310 184.095 ;
        RECT 215.985 184.050 216.305 184.110 ;
        RECT 210.020 183.910 216.305 184.050 ;
        RECT 210.020 183.865 210.310 183.910 ;
        RECT 215.985 183.850 216.305 183.910 ;
        RECT 216.445 184.050 216.765 184.110 ;
        RECT 217.840 184.050 218.130 184.095 ;
        RECT 219.665 184.050 219.985 184.110 ;
        RECT 216.445 183.910 218.130 184.050 ;
        RECT 216.445 183.850 216.765 183.910 ;
        RECT 217.840 183.865 218.130 183.910 ;
        RECT 218.835 183.910 219.985 184.050 ;
        RECT 203.580 183.525 203.870 183.755 ;
        RECT 204.485 183.710 204.805 183.770 ;
        RECT 210.465 183.755 210.785 183.770 ;
        RECT 206.340 183.710 206.630 183.755 ;
        RECT 204.485 183.570 206.630 183.710 ;
        RECT 204.485 183.510 204.805 183.570 ;
        RECT 206.340 183.525 206.630 183.570 ;
        RECT 207.725 183.710 208.015 183.755 ;
        RECT 209.565 183.710 209.855 183.755 ;
        RECT 207.725 183.570 209.855 183.710 ;
        RECT 207.725 183.525 208.015 183.570 ;
        RECT 209.565 183.525 209.855 183.570 ;
        RECT 210.465 183.525 210.895 183.755 ;
        RECT 210.465 183.510 210.785 183.525 ;
        RECT 211.385 183.510 211.705 183.770 ;
        RECT 211.910 183.710 212.200 183.755 ;
        RECT 213.750 183.710 214.040 183.755 ;
        RECT 211.910 183.570 214.040 183.710 ;
        RECT 211.910 183.525 212.200 183.570 ;
        RECT 213.750 183.525 214.040 183.570 ;
        RECT 214.605 183.710 214.925 183.770 ;
        RECT 215.080 183.710 215.370 183.755 ;
        RECT 214.605 183.570 215.370 183.710 ;
        RECT 214.605 183.510 214.925 183.570 ;
        RECT 215.080 183.525 215.370 183.570 ;
        RECT 216.920 183.710 217.210 183.755 ;
        RECT 218.835 183.710 218.975 183.910 ;
        RECT 219.665 183.850 219.985 183.910 ;
        RECT 220.125 183.850 220.445 184.110 ;
        RECT 220.675 184.050 220.815 184.590 ;
        RECT 221.100 184.390 221.390 184.435 ;
        RECT 224.330 184.390 224.620 184.435 ;
        RECT 221.100 184.250 224.620 184.390 ;
        RECT 221.100 184.205 221.390 184.250 ;
        RECT 224.330 184.205 224.620 184.250 ;
        RECT 222.105 184.050 222.395 184.095 ;
        RECT 220.675 183.910 222.395 184.050 ;
        RECT 224.815 184.050 224.955 184.590 ;
        RECT 225.645 184.590 227.330 184.730 ;
        RECT 225.645 184.530 225.965 184.590 ;
        RECT 227.040 184.545 227.330 184.590 ;
        RECT 228.035 184.590 230.565 184.730 ;
        RECT 226.120 184.390 226.410 184.435 ;
        RECT 228.035 184.390 228.175 184.590 ;
        RECT 230.245 184.530 230.565 184.590 ;
        RECT 226.120 184.250 228.175 184.390 ;
        RECT 226.120 184.205 226.410 184.250 ;
        RECT 228.420 184.205 228.710 184.435 ;
        RECT 228.495 184.050 228.635 184.205 ;
        RECT 231.625 184.050 231.945 184.110 ;
        RECT 224.815 183.910 228.635 184.050 ;
        RECT 229.415 183.910 231.945 184.050 ;
        RECT 222.105 183.865 222.395 183.910 ;
        RECT 216.920 183.570 218.975 183.710 ;
        RECT 219.225 183.710 219.515 183.755 ;
        RECT 221.065 183.710 221.355 183.755 ;
        RECT 219.225 183.570 221.355 183.710 ;
        RECT 216.920 183.525 217.210 183.570 ;
        RECT 219.225 183.525 219.515 183.570 ;
        RECT 221.065 183.525 221.355 183.570 ;
        RECT 221.505 183.510 221.825 183.770 ;
        RECT 222.885 183.510 223.205 183.770 ;
        RECT 223.410 183.710 223.700 183.755 ;
        RECT 225.250 183.710 225.540 183.755 ;
        RECT 223.410 183.570 225.540 183.710 ;
        RECT 223.410 183.525 223.700 183.570 ;
        RECT 225.250 183.525 225.540 183.570 ;
        RECT 227.945 183.510 228.265 183.770 ;
        RECT 229.415 183.755 229.555 183.910 ;
        RECT 231.625 183.850 231.945 183.910 ;
        RECT 229.340 183.525 229.630 183.755 ;
        RECT 230.245 183.710 230.565 183.770 ;
        RECT 230.720 183.710 231.010 183.755 ;
        RECT 230.245 183.570 231.010 183.710 ;
        RECT 230.245 183.510 230.565 183.570 ;
        RECT 230.720 183.525 231.010 183.570 ;
        RECT 232.100 183.525 232.390 183.755 ;
        RECT 206.805 183.370 207.095 183.415 ;
        RECT 212.325 183.370 212.615 183.415 ;
        RECT 213.245 183.370 213.535 183.415 ;
        RECT 206.805 183.230 213.535 183.370 ;
        RECT 206.805 183.185 207.095 183.230 ;
        RECT 212.325 183.185 212.615 183.230 ;
        RECT 213.245 183.185 213.535 183.230 ;
        RECT 218.305 183.370 218.595 183.415 ;
        RECT 223.825 183.370 224.115 183.415 ;
        RECT 224.745 183.370 225.035 183.415 ;
        RECT 218.305 183.230 225.035 183.370 ;
        RECT 218.305 183.185 218.595 183.230 ;
        RECT 223.825 183.185 224.115 183.230 ;
        RECT 224.745 183.185 225.035 183.230 ;
        RECT 225.645 183.370 225.965 183.430 ;
        RECT 232.175 183.370 232.315 183.525 ;
        RECT 233.465 183.510 233.785 183.770 ;
        RECT 225.645 183.230 232.315 183.370 ;
        RECT 225.645 183.170 225.965 183.230 ;
        RECT 207.245 183.030 207.565 183.090 ;
        RECT 203.195 182.890 207.565 183.030 ;
        RECT 201.725 182.830 202.045 182.890 ;
        RECT 202.660 182.845 202.950 182.890 ;
        RECT 207.245 182.830 207.565 182.890 ;
        RECT 209.085 183.030 209.405 183.090 ;
        RECT 215.525 183.030 215.845 183.090 ;
        RECT 209.085 182.890 215.845 183.030 ;
        RECT 209.085 182.830 209.405 182.890 ;
        RECT 215.525 182.830 215.845 182.890 ;
        RECT 216.000 183.030 216.290 183.075 ;
        RECT 223.345 183.030 223.665 183.090 ;
        RECT 216.000 182.890 223.665 183.030 ;
        RECT 216.000 182.845 216.290 182.890 ;
        RECT 223.345 182.830 223.665 182.890 ;
        RECT 224.265 183.030 224.585 183.090 ;
        RECT 227.025 183.030 227.345 183.090 ;
        RECT 224.265 182.890 227.345 183.030 ;
        RECT 224.265 182.830 224.585 182.890 ;
        RECT 227.025 182.830 227.345 182.890 ;
        RECT 229.785 182.830 230.105 183.090 ;
        RECT 231.165 182.830 231.485 183.090 ;
        RECT 232.545 182.830 232.865 183.090 ;
        RECT 63.895 181.400 64.595 182.400 ;
        RECT 77.595 182.370 78.595 182.605 ;
        RECT 77.595 181.195 78.595 181.430 ;
        RECT 80.185 181.400 81.755 182.400 ;
        RECT 83.345 182.370 84.345 182.605 ;
        RECT 83.345 181.195 84.345 181.430 ;
        RECT 97.345 181.400 98.045 182.400 ;
        RECT 64.175 180.965 80.135 181.195 ;
        RECT 81.805 180.965 97.765 181.195 ;
        RECT 77.595 180.730 78.595 180.965 ;
        RECT 83.345 180.730 84.345 180.965 ;
        RECT 98.485 180.110 155.900 182.710 ;
        RECT 162.095 182.210 236.155 182.690 ;
        RECT 167.685 181.810 168.005 182.070 ;
        RECT 171.380 182.010 171.670 182.055 ;
        RECT 173.665 182.010 173.985 182.070 ;
        RECT 171.380 181.870 173.985 182.010 ;
        RECT 171.380 181.825 171.670 181.870 ;
        RECT 173.665 181.810 173.985 181.870 ;
        RECT 175.505 182.010 175.825 182.070 ;
        RECT 179.660 182.010 179.950 182.055 ;
        RECT 175.505 181.870 179.950 182.010 ;
        RECT 175.505 181.810 175.825 181.870 ;
        RECT 179.660 181.825 179.950 181.870 ;
        RECT 180.565 182.010 180.885 182.070 ;
        RECT 181.500 182.010 181.790 182.055 ;
        RECT 180.565 181.870 181.790 182.010 ;
        RECT 180.565 181.810 180.885 181.870 ;
        RECT 181.500 181.825 181.790 181.870 ;
        RECT 183.325 182.010 183.645 182.070 ;
        RECT 185.640 182.010 185.930 182.055 ;
        RECT 183.325 181.870 185.930 182.010 ;
        RECT 183.325 181.810 183.645 181.870 ;
        RECT 185.640 181.825 185.930 181.870 ;
        RECT 186.085 181.810 186.405 182.070 ;
        RECT 187.465 182.010 187.785 182.070 ;
        RECT 188.860 182.010 189.150 182.055 ;
        RECT 187.465 181.870 189.150 182.010 ;
        RECT 187.465 181.810 187.785 181.870 ;
        RECT 188.860 181.825 189.150 181.870 ;
        RECT 190.225 182.010 190.545 182.070 ;
        RECT 193.460 182.010 193.750 182.055 ;
        RECT 190.225 181.870 193.750 182.010 ;
        RECT 190.225 181.810 190.545 181.870 ;
        RECT 193.460 181.825 193.750 181.870 ;
        RECT 195.760 182.010 196.050 182.055 ;
        RECT 198.520 182.010 198.810 182.055 ;
        RECT 195.760 181.870 198.810 182.010 ;
        RECT 195.760 181.825 196.050 181.870 ;
        RECT 198.520 181.825 198.810 181.870 ;
        RECT 202.200 182.010 202.490 182.055 ;
        RECT 203.580 182.010 203.870 182.055 ;
        RECT 212.305 182.010 212.625 182.070 ;
        RECT 202.200 181.870 203.335 182.010 ;
        RECT 202.200 181.825 202.490 181.870 ;
        RECT 166.305 181.670 166.625 181.730 ;
        RECT 169.525 181.670 169.845 181.730 ;
        RECT 172.285 181.670 172.605 181.730 ;
        RECT 178.265 181.670 178.585 181.730 ;
        RECT 164.555 181.530 166.625 181.670 ;
        RECT 164.555 181.375 164.695 181.530 ;
        RECT 166.305 181.470 166.625 181.530 ;
        RECT 166.855 181.530 174.355 181.670 ;
        RECT 166.855 181.375 166.995 181.530 ;
        RECT 169.525 181.470 169.845 181.530 ;
        RECT 164.480 181.145 164.770 181.375 ;
        RECT 165.400 181.145 165.690 181.375 ;
        RECT 166.780 181.145 167.070 181.375 ;
        RECT 168.160 181.330 168.450 181.375 ;
        RECT 167.775 181.190 168.450 181.330 ;
        RECT 165.475 180.990 165.615 181.145 ;
        RECT 167.775 180.990 167.915 181.190 ;
        RECT 168.160 181.145 168.450 181.190 ;
        RECT 169.080 181.330 169.370 181.375 ;
        RECT 169.080 181.280 169.750 181.330 ;
        RECT 169.985 181.280 170.305 181.390 ;
        RECT 170.535 181.375 170.675 181.530 ;
        RECT 172.285 181.470 172.605 181.530 ;
        RECT 169.080 181.190 170.305 181.280 ;
        RECT 169.080 181.145 169.370 181.190 ;
        RECT 169.610 181.140 170.305 181.190 ;
        RECT 170.460 181.145 170.750 181.375 ;
        RECT 171.840 181.145 172.130 181.375 ;
        RECT 169.985 181.130 170.305 181.140 ;
        RECT 168.605 180.990 168.925 181.050 ;
        RECT 171.365 180.990 171.685 181.050 ;
        RECT 171.915 180.990 172.055 181.145 ;
        RECT 172.745 181.130 173.065 181.390 ;
        RECT 174.215 181.375 174.355 181.530 ;
        RECT 175.595 181.530 178.585 181.670 ;
        RECT 175.595 181.375 175.735 181.530 ;
        RECT 178.265 181.470 178.585 181.530 ;
        RECT 178.740 181.670 179.030 181.715 ;
        RECT 181.945 181.670 182.265 181.730 ;
        RECT 178.740 181.530 182.265 181.670 ;
        RECT 178.740 181.485 179.030 181.530 ;
        RECT 181.945 181.470 182.265 181.530 ;
        RECT 184.705 181.670 185.025 181.730 ;
        RECT 190.700 181.670 190.990 181.715 ;
        RECT 184.705 181.530 190.990 181.670 ;
        RECT 184.705 181.470 185.025 181.530 ;
        RECT 190.700 181.485 190.990 181.530 ;
        RECT 191.160 181.670 191.450 181.715 ;
        RECT 200.805 181.670 201.125 181.730 ;
        RECT 201.725 181.670 202.045 181.730 ;
        RECT 191.160 181.530 201.125 181.670 ;
        RECT 191.160 181.485 191.450 181.530 ;
        RECT 200.805 181.470 201.125 181.530 ;
        RECT 201.355 181.530 202.045 181.670 ;
        RECT 203.195 181.670 203.335 181.870 ;
        RECT 203.580 181.870 212.625 182.010 ;
        RECT 203.580 181.825 203.870 181.870 ;
        RECT 212.305 181.810 212.625 181.870 ;
        RECT 213.240 182.010 213.530 182.055 ;
        RECT 213.685 182.010 214.005 182.070 ;
        RECT 213.240 181.870 214.005 182.010 ;
        RECT 213.240 181.825 213.530 181.870 ;
        RECT 213.685 181.810 214.005 181.870 ;
        RECT 215.985 182.010 216.305 182.070 ;
        RECT 233.480 182.010 233.770 182.055 ;
        RECT 215.985 181.870 233.770 182.010 ;
        RECT 215.985 181.810 216.305 181.870 ;
        RECT 233.480 181.825 233.770 181.870 ;
        RECT 204.945 181.670 205.265 181.730 ;
        RECT 203.195 181.530 205.265 181.670 ;
        RECT 174.140 181.145 174.430 181.375 ;
        RECT 175.060 181.145 175.350 181.375 ;
        RECT 175.520 181.145 175.810 181.375 ;
        RECT 165.475 180.850 172.055 180.990 ;
        RECT 175.135 180.990 175.275 181.145 ;
        RECT 176.425 181.130 176.745 181.390 ;
        RECT 176.885 181.330 177.205 181.390 ;
        RECT 177.820 181.330 178.110 181.375 ;
        RECT 176.885 181.190 178.110 181.330 ;
        RECT 176.885 181.130 177.205 181.190 ;
        RECT 177.820 181.145 178.110 181.190 ;
        RECT 179.645 181.330 179.965 181.390 ;
        RECT 183.325 181.330 183.645 181.390 ;
        RECT 179.645 181.190 183.645 181.330 ;
        RECT 179.645 181.130 179.965 181.190 ;
        RECT 183.325 181.130 183.645 181.190 ;
        RECT 185.165 181.330 185.485 181.390 ;
        RECT 189.305 181.330 189.625 181.390 ;
        RECT 185.165 181.190 189.625 181.330 ;
        RECT 185.165 181.130 185.485 181.190 ;
        RECT 189.305 181.130 189.625 181.190 ;
        RECT 195.300 181.145 195.590 181.375 ;
        RECT 198.505 181.330 198.825 181.390 ;
        RECT 201.355 181.375 201.495 181.530 ;
        RECT 201.725 181.470 202.045 181.530 ;
        RECT 204.945 181.470 205.265 181.530 ;
        RECT 205.425 181.670 205.715 181.715 ;
        RECT 210.945 181.670 211.235 181.715 ;
        RECT 211.865 181.670 212.155 181.715 ;
        RECT 205.425 181.530 212.155 181.670 ;
        RECT 205.425 181.485 205.715 181.530 ;
        RECT 210.945 181.485 211.235 181.530 ;
        RECT 211.865 181.485 212.155 181.530 ;
        RECT 215.545 181.670 215.835 181.715 ;
        RECT 221.065 181.670 221.355 181.715 ;
        RECT 221.985 181.670 222.275 181.715 ;
        RECT 215.545 181.530 222.275 181.670 ;
        RECT 215.545 181.485 215.835 181.530 ;
        RECT 221.065 181.485 221.355 181.530 ;
        RECT 221.985 181.485 222.275 181.530 ;
        RECT 225.205 181.670 225.495 181.715 ;
        RECT 230.725 181.670 231.015 181.715 ;
        RECT 231.645 181.670 231.935 181.715 ;
        RECT 225.205 181.530 231.935 181.670 ;
        RECT 225.205 181.485 225.495 181.530 ;
        RECT 230.725 181.485 231.015 181.530 ;
        RECT 231.645 181.485 231.935 181.530 ;
        RECT 199.440 181.330 199.730 181.375 ;
        RECT 198.505 181.190 199.730 181.330 ;
        RECT 181.025 180.990 181.345 181.050 ;
        RECT 181.960 180.990 182.250 181.035 ;
        RECT 175.135 180.850 178.035 180.990 ;
        RECT 168.605 180.790 168.925 180.850 ;
        RECT 171.365 180.790 171.685 180.850 ;
        RECT 177.895 180.710 178.035 180.850 ;
        RECT 181.025 180.850 182.250 180.990 ;
        RECT 181.025 180.790 181.345 180.850 ;
        RECT 181.960 180.805 182.250 180.850 ;
        RECT 182.405 180.790 182.725 181.050 ;
        RECT 186.545 180.990 186.865 181.050 ;
        RECT 187.020 180.990 187.310 181.035 ;
        RECT 192.080 180.990 192.370 181.035 ;
        RECT 192.525 180.990 192.845 181.050 ;
        RECT 182.955 180.850 184.475 180.990 ;
        RECT 166.765 180.650 167.085 180.710 ;
        RECT 175.505 180.650 175.825 180.710 ;
        RECT 166.765 180.510 175.825 180.650 ;
        RECT 166.765 180.450 167.085 180.510 ;
        RECT 175.505 180.450 175.825 180.510 ;
        RECT 177.805 180.450 178.125 180.710 ;
        RECT 179.645 180.650 179.965 180.710 ;
        RECT 182.955 180.650 183.095 180.850 ;
        RECT 179.645 180.510 183.095 180.650 ;
        RECT 179.645 180.450 179.965 180.510 ;
        RECT 183.785 180.450 184.105 180.710 ;
        RECT 184.335 180.650 184.475 180.850 ;
        RECT 186.545 180.850 192.845 180.990 ;
        RECT 186.545 180.790 186.865 180.850 ;
        RECT 187.020 180.805 187.310 180.850 ;
        RECT 192.080 180.805 192.370 180.850 ;
        RECT 192.525 180.790 192.845 180.850 ;
        RECT 195.375 180.650 195.515 181.145 ;
        RECT 198.505 181.130 198.825 181.190 ;
        RECT 199.440 181.145 199.730 181.190 ;
        RECT 199.900 181.145 200.190 181.375 ;
        RECT 201.280 181.145 201.570 181.375 ;
        RECT 202.185 181.330 202.505 181.390 ;
        RECT 202.660 181.330 202.950 181.375 ;
        RECT 202.185 181.190 202.950 181.330 ;
        RECT 196.680 180.805 196.970 181.035 ;
        RECT 199.975 180.990 200.115 181.145 ;
        RECT 202.185 181.130 202.505 181.190 ;
        RECT 202.660 181.145 202.950 181.190 ;
        RECT 204.025 181.130 204.345 181.390 ;
        RECT 206.345 181.330 206.635 181.375 ;
        RECT 208.185 181.330 208.475 181.375 ;
        RECT 206.345 181.190 208.475 181.330 ;
        RECT 206.345 181.145 206.635 181.190 ;
        RECT 208.185 181.145 208.475 181.190 ;
        RECT 208.625 181.130 208.945 181.390 ;
        RECT 209.330 181.330 209.620 181.375 ;
        RECT 209.300 181.310 209.620 181.330 ;
        RECT 209.085 181.145 209.620 181.310 ;
        RECT 209.085 181.110 209.440 181.145 ;
        RECT 210.005 181.130 210.325 181.390 ;
        RECT 210.530 181.330 210.820 181.375 ;
        RECT 212.370 181.330 212.660 181.375 ;
        RECT 210.530 181.190 212.660 181.330 ;
        RECT 210.530 181.145 210.820 181.190 ;
        RECT 212.370 181.145 212.660 181.190 ;
        RECT 214.145 181.130 214.465 181.390 ;
        RECT 216.465 181.330 216.755 181.375 ;
        RECT 218.305 181.330 218.595 181.375 ;
        RECT 216.465 181.190 218.595 181.330 ;
        RECT 216.465 181.145 216.755 181.190 ;
        RECT 218.305 181.145 218.595 181.190 ;
        RECT 220.650 181.330 220.940 181.375 ;
        RECT 222.490 181.330 222.780 181.375 ;
        RECT 220.650 181.190 222.780 181.330 ;
        RECT 220.650 181.145 220.940 181.190 ;
        RECT 222.490 181.145 222.780 181.190 ;
        RECT 223.345 181.330 223.665 181.390 ;
        RECT 223.820 181.330 224.110 181.375 ;
        RECT 226.125 181.330 226.415 181.375 ;
        RECT 227.965 181.330 228.255 181.375 ;
        RECT 228.510 181.330 228.800 181.375 ;
        RECT 223.345 181.190 224.110 181.330 ;
        RECT 223.345 181.130 223.665 181.190 ;
        RECT 223.820 181.145 224.110 181.190 ;
        RECT 224.355 181.190 225.415 181.330 ;
        RECT 209.085 181.050 209.405 181.110 ;
        RECT 224.355 181.050 224.495 181.190 ;
        RECT 201.725 180.990 202.045 181.050 ;
        RECT 204.960 180.990 205.250 181.035 ;
        RECT 199.975 180.850 201.495 180.990 ;
        RECT 184.335 180.510 195.515 180.650 ;
        RECT 164.465 180.310 164.785 180.370 ;
        RECT 167.685 180.310 168.005 180.370 ;
        RECT 164.465 180.170 168.005 180.310 ;
        RECT 164.465 180.110 164.785 180.170 ;
        RECT 167.685 180.110 168.005 180.170 ;
        RECT 169.065 180.310 169.385 180.370 ;
        RECT 179.185 180.310 179.505 180.370 ;
        RECT 169.065 180.170 179.505 180.310 ;
        RECT 169.065 180.110 169.385 180.170 ;
        RECT 179.185 180.110 179.505 180.170 ;
        RECT 181.945 180.310 182.265 180.370 ;
        RECT 186.085 180.310 186.405 180.370 ;
        RECT 181.945 180.170 186.405 180.310 ;
        RECT 196.755 180.310 196.895 180.805 ;
        RECT 200.805 180.450 201.125 180.710 ;
        RECT 201.355 180.650 201.495 180.850 ;
        RECT 201.725 180.850 205.250 180.990 ;
        RECT 201.725 180.790 202.045 180.850 ;
        RECT 204.960 180.805 205.250 180.850 ;
        RECT 213.685 180.990 214.005 181.050 ;
        RECT 215.080 180.990 215.370 181.035 ;
        RECT 213.685 180.850 215.370 180.990 ;
        RECT 213.685 180.790 214.005 180.850 ;
        RECT 215.080 180.805 215.370 180.850 ;
        RECT 217.380 180.805 217.670 181.035 ;
        RECT 204.025 180.650 204.345 180.710 ;
        RECT 201.355 180.510 204.345 180.650 ;
        RECT 204.025 180.450 204.345 180.510 ;
        RECT 206.325 180.650 206.645 180.710 ;
        RECT 207.260 180.650 207.550 180.695 ;
        RECT 206.325 180.510 207.550 180.650 ;
        RECT 206.325 180.450 206.645 180.510 ;
        RECT 206.875 180.310 207.015 180.510 ;
        RECT 207.260 180.465 207.550 180.510 ;
        RECT 208.220 180.650 208.510 180.695 ;
        RECT 211.450 180.650 211.740 180.695 ;
        RECT 217.455 180.650 217.595 180.805 ;
        RECT 218.745 180.790 219.065 181.050 ;
        RECT 219.665 181.035 219.985 181.050 ;
        RECT 219.450 180.805 219.985 181.035 ;
        RECT 220.140 180.990 220.430 181.035 ;
        RECT 221.045 180.990 221.365 181.050 ;
        RECT 224.265 180.990 224.585 181.050 ;
        RECT 220.140 180.850 224.585 180.990 ;
        RECT 220.140 180.805 220.430 180.850 ;
        RECT 219.665 180.790 219.985 180.805 ;
        RECT 221.045 180.790 221.365 180.850 ;
        RECT 224.265 180.790 224.585 180.850 ;
        RECT 224.725 180.790 225.045 181.050 ;
        RECT 225.275 180.990 225.415 181.190 ;
        RECT 226.125 181.190 228.255 181.330 ;
        RECT 228.495 181.310 228.800 181.330 ;
        RECT 226.125 181.145 226.415 181.190 ;
        RECT 227.965 181.145 228.255 181.190 ;
        RECT 228.405 181.145 228.800 181.310 ;
        RECT 230.310 181.330 230.600 181.375 ;
        RECT 232.150 181.330 232.440 181.375 ;
        RECT 230.310 181.190 232.440 181.330 ;
        RECT 230.310 181.145 230.600 181.190 ;
        RECT 232.150 181.145 232.440 181.190 ;
        RECT 228.405 181.050 228.725 181.145 ;
        RECT 234.385 181.130 234.705 181.390 ;
        RECT 229.325 181.035 229.645 181.050 ;
        RECT 225.275 180.850 227.715 180.990 ;
        RECT 218.340 180.650 218.630 180.695 ;
        RECT 221.570 180.650 221.860 180.695 ;
        RECT 227.040 180.650 227.330 180.695 ;
        RECT 208.220 180.510 211.740 180.650 ;
        RECT 208.220 180.465 208.510 180.510 ;
        RECT 211.450 180.465 211.740 180.510 ;
        RECT 214.695 180.510 218.055 180.650 ;
        RECT 210.005 180.310 210.325 180.370 ;
        RECT 214.695 180.310 214.835 180.510 ;
        RECT 196.755 180.170 214.835 180.310 ;
        RECT 215.525 180.310 215.845 180.370 ;
        RECT 217.365 180.310 217.685 180.370 ;
        RECT 215.525 180.170 217.685 180.310 ;
        RECT 217.915 180.310 218.055 180.510 ;
        RECT 218.340 180.510 221.860 180.650 ;
        RECT 218.340 180.465 218.630 180.510 ;
        RECT 221.570 180.465 221.860 180.510 ;
        RECT 222.975 180.510 227.330 180.650 ;
        RECT 222.975 180.310 223.115 180.510 ;
        RECT 227.040 180.465 227.330 180.510 ;
        RECT 217.915 180.170 223.115 180.310 ;
        RECT 181.945 180.110 182.265 180.170 ;
        RECT 186.085 180.110 186.405 180.170 ;
        RECT 210.005 180.110 210.325 180.170 ;
        RECT 215.525 180.110 215.845 180.170 ;
        RECT 217.365 180.110 217.685 180.170 ;
        RECT 223.345 180.110 223.665 180.370 ;
        RECT 223.805 180.310 224.125 180.370 ;
        RECT 225.645 180.310 225.965 180.370 ;
        RECT 223.805 180.170 225.965 180.310 ;
        RECT 227.575 180.310 227.715 180.850 ;
        RECT 229.110 180.805 229.645 181.035 ;
        RECT 229.800 180.990 230.090 181.035 ;
        RECT 229.800 180.850 231.855 180.990 ;
        RECT 229.800 180.805 230.090 180.850 ;
        RECT 229.325 180.790 229.645 180.805 ;
        RECT 228.000 180.650 228.290 180.695 ;
        RECT 231.230 180.650 231.520 180.695 ;
        RECT 228.000 180.510 231.520 180.650 ;
        RECT 228.000 180.465 228.290 180.510 ;
        RECT 231.230 180.465 231.520 180.510 ;
        RECT 231.715 180.310 231.855 180.850 ;
        RECT 227.575 180.170 231.855 180.310 ;
        RECT 223.805 180.110 224.125 180.170 ;
        RECT 225.645 180.110 225.965 180.170 ;
        RECT 233.005 180.110 233.325 180.370 ;
        RECT 77.595 179.815 78.595 180.050 ;
        RECT 83.345 179.815 84.345 180.050 ;
        RECT 64.175 179.585 80.135 179.815 ;
        RECT 81.805 179.585 97.765 179.815 ;
        RECT 63.895 178.380 64.595 179.380 ;
        RECT 77.595 179.350 78.595 179.585 ;
        RECT 77.595 178.175 78.595 178.410 ;
        RECT 80.185 178.380 81.755 179.380 ;
        RECT 83.345 179.350 84.345 179.585 ;
        RECT 83.345 178.175 84.345 178.410 ;
        RECT 97.345 178.380 98.045 179.380 ;
        RECT 64.175 177.945 80.135 178.175 ;
        RECT 81.805 177.945 97.765 178.175 ;
        RECT 77.595 177.710 78.595 177.945 ;
        RECT 83.345 177.710 84.345 177.945 ;
        RECT 77.595 176.795 78.595 177.030 ;
        RECT 83.345 176.795 84.345 177.030 ;
        RECT 64.175 176.565 80.135 176.795 ;
        RECT 81.805 176.565 97.765 176.795 ;
        RECT 63.895 175.360 64.595 176.360 ;
        RECT 77.595 176.330 78.595 176.565 ;
        RECT 77.595 175.155 78.595 175.390 ;
        RECT 80.185 175.360 81.755 176.360 ;
        RECT 83.345 176.330 84.345 176.565 ;
        RECT 83.345 175.155 84.345 175.390 ;
        RECT 97.345 175.360 98.045 176.360 ;
        RECT 64.175 174.925 80.135 175.155 ;
        RECT 81.805 174.925 97.765 175.155 ;
        RECT 77.595 174.690 78.595 174.925 ;
        RECT 83.345 174.690 84.345 174.925 ;
        RECT 64.175 173.545 80.135 173.775 ;
        RECT 81.805 173.545 97.765 173.775 ;
        RECT 63.895 172.340 64.125 173.340 ;
        RECT 80.185 172.340 81.755 173.340 ;
        RECT 97.815 172.340 98.045 173.340 ;
        RECT 64.175 171.905 80.135 172.135 ;
        RECT 81.805 171.905 97.765 172.135 ;
        RECT 98.485 171.445 100.480 180.110 ;
        RECT 62.865 160.555 100.480 171.445 ;
        RECT 5.910 143.155 58.705 143.745 ;
        RECT 5.910 140.725 23.785 143.155 ;
        RECT 24.505 143.045 25.505 143.155 ;
        RECT 24.255 142.435 57.645 142.665 ;
        RECT 24.255 141.275 24.485 142.435 ;
        RECT 28.015 141.965 29.015 142.435 ;
        RECT 32.545 141.275 32.775 142.435 ;
        RECT 36.305 141.965 37.305 142.435 ;
        RECT 40.835 141.275 41.065 142.435 ;
        RECT 44.595 141.965 45.595 142.435 ;
        RECT 49.125 141.275 49.355 142.435 ;
        RECT 52.885 141.965 53.885 142.435 ;
        RECT 57.415 141.275 57.645 142.435 ;
        RECT 24.535 140.885 32.495 141.115 ;
        RECT 32.825 140.885 40.785 141.115 ;
        RECT 41.115 140.885 49.075 141.115 ;
        RECT 49.405 140.885 57.365 141.115 ;
        RECT 5.910 139.725 24.955 140.725 ;
        RECT 32.545 139.725 32.775 140.725 ;
        RECT 40.835 139.725 41.065 140.725 ;
        RECT 49.125 139.725 49.355 140.725 ;
        RECT 56.545 139.725 57.645 140.725 ;
        RECT 5.910 139.175 23.785 139.725 ;
        RECT 24.535 139.335 32.495 139.565 ;
        RECT 32.825 139.335 40.785 139.565 ;
        RECT 41.115 139.335 49.075 139.565 ;
        RECT 49.405 139.335 57.365 139.565 ;
        RECT 5.910 138.175 24.955 139.175 ;
        RECT 32.545 138.175 32.775 139.175 ;
        RECT 40.835 138.175 41.065 139.175 ;
        RECT 49.125 138.175 49.355 139.175 ;
        RECT 53.035 138.175 57.645 139.175 ;
        RECT 5.910 137.925 23.785 138.175 ;
        RECT 5.910 137.075 9.990 137.925 ;
        RECT 11.145 137.465 11.845 137.535 ;
        RECT 14.080 137.465 14.780 137.535 ;
        RECT 15.370 137.465 16.070 137.535 ;
        RECT 18.305 137.465 19.005 137.535 ;
        RECT 11.015 137.235 11.975 137.465 ;
        RECT 13.950 137.235 14.910 137.465 ;
        RECT 15.240 137.235 16.200 137.465 ;
        RECT 18.175 137.235 19.135 137.465 ;
        RECT 5.910 136.075 10.965 137.075 ;
        RECT 12.025 136.925 12.255 137.075 ;
        RECT 11.990 136.225 12.290 136.925 ;
        RECT 12.025 136.075 12.255 136.225 ;
        RECT 5.910 135.225 9.990 136.075 ;
        RECT 13.670 135.825 13.900 137.075 ;
        RECT 14.960 136.925 15.190 137.075 ;
        RECT 16.250 136.925 16.480 137.075 ;
        RECT 14.925 136.225 15.225 136.925 ;
        RECT 16.215 136.225 16.515 136.925 ;
        RECT 14.960 136.075 15.190 136.225 ;
        RECT 16.250 136.075 16.480 136.225 ;
        RECT 13.435 135.525 14.135 135.825 ;
        RECT 17.895 135.225 18.125 137.075 ;
        RECT 19.185 136.775 19.415 137.075 ;
        RECT 19.150 136.075 19.450 136.775 ;
        RECT 20.160 135.745 23.785 137.925 ;
        RECT 24.535 137.785 32.495 138.015 ;
        RECT 32.825 137.785 40.785 138.015 ;
        RECT 41.115 137.785 49.075 138.015 ;
        RECT 49.405 137.785 57.365 138.015 ;
        RECT 24.255 136.465 24.485 137.625 ;
        RECT 28.015 136.465 29.015 136.935 ;
        RECT 32.545 136.465 32.775 137.625 ;
        RECT 36.305 136.465 37.305 136.935 ;
        RECT 40.835 136.465 41.065 137.625 ;
        RECT 44.595 136.465 45.595 136.935 ;
        RECT 49.125 136.465 49.355 137.625 ;
        RECT 52.885 136.465 53.885 136.935 ;
        RECT 57.415 136.465 57.645 137.625 ;
        RECT 24.255 136.235 57.645 136.465 ;
        RECT 24.505 135.745 25.505 135.855 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 20.160 135.225 58.705 135.745 ;
        RECT 5.910 132.225 58.705 135.225 ;
        RECT 62.865 139.455 69.970 160.555 ;
        RECT 71.220 157.040 89.820 159.315 ;
        RECT 71.220 142.990 73.495 157.040 ;
        RECT 76.385 157.030 77.215 157.040 ;
        RECT 80.105 157.030 80.935 157.040 ;
        RECT 83.825 157.030 84.655 157.040 ;
        RECT 74.940 154.420 86.100 155.595 ;
        RECT 74.940 153.050 76.115 154.420 ;
        RECT 76.385 153.310 77.215 154.140 ;
        RECT 77.485 153.050 79.835 154.420 ;
        RECT 80.105 153.310 80.935 154.140 ;
        RECT 81.205 153.050 83.555 154.420 ;
        RECT 83.825 153.310 84.655 154.140 ;
        RECT 84.925 153.050 86.100 154.420 ;
        RECT 74.940 150.700 86.100 153.050 ;
        RECT 74.940 149.330 76.115 150.700 ;
        RECT 76.385 149.590 77.215 150.420 ;
        RECT 77.485 149.330 79.835 150.700 ;
        RECT 80.105 149.590 80.935 150.420 ;
        RECT 81.205 149.330 83.555 150.700 ;
        RECT 83.825 149.590 84.655 150.420 ;
        RECT 84.925 149.330 86.100 150.700 ;
        RECT 74.940 146.980 86.100 149.330 ;
        RECT 74.940 145.610 76.115 146.980 ;
        RECT 76.385 145.870 77.215 146.700 ;
        RECT 77.485 145.610 79.835 146.980 ;
        RECT 80.105 145.870 80.935 146.700 ;
        RECT 81.205 145.610 83.555 146.980 ;
        RECT 83.825 145.870 84.655 146.700 ;
        RECT 84.925 145.610 86.100 146.980 ;
        RECT 74.940 144.435 86.100 145.610 ;
        RECT 87.545 142.990 89.820 157.040 ;
        RECT 71.220 140.715 89.820 142.990 ;
        RECT 91.070 139.455 100.480 160.555 ;
        RECT 101.935 176.325 152.755 178.210 ;
        RECT 101.935 174.870 114.420 176.325 ;
        RECT 115.200 175.635 118.030 176.165 ;
        RECT 119.820 175.635 122.650 176.165 ;
        RECT 124.440 175.635 127.270 176.165 ;
        RECT 129.060 175.635 131.890 176.165 ;
        RECT 133.680 175.635 136.510 176.165 ;
        RECT 138.300 175.635 141.130 176.165 ;
        RECT 142.920 175.635 145.750 176.165 ;
        RECT 147.540 175.635 150.370 176.165 ;
        RECT 114.920 174.870 115.150 175.475 ;
        RECT 101.935 172.215 115.185 174.870 ;
        RECT 101.935 162.685 103.025 172.215 ;
        RECT 103.715 171.610 104.675 171.840 ;
        RECT 105.005 171.610 105.965 171.840 ;
        RECT 103.435 170.840 103.665 171.450 ;
        RECT 103.400 168.540 103.700 170.840 ;
        RECT 103.435 163.450 103.665 168.540 ;
        RECT 104.725 167.140 104.955 171.450 ;
        RECT 106.015 170.840 106.245 171.450 ;
        RECT 105.980 168.540 106.280 170.840 ;
        RECT 104.690 164.840 104.990 167.140 ;
        RECT 104.725 163.450 104.955 164.840 ;
        RECT 106.015 163.450 106.245 168.540 ;
        RECT 103.715 163.060 104.675 163.290 ;
        RECT 105.005 163.060 105.965 163.290 ;
        RECT 103.715 162.990 104.415 163.060 ;
        RECT 105.265 162.990 105.965 163.060 ;
        RECT 106.655 162.685 107.055 172.215 ;
        RECT 110.685 172.070 115.185 172.215 ;
        RECT 107.745 171.610 108.705 171.840 ;
        RECT 109.035 171.610 109.995 171.840 ;
        RECT 107.465 170.840 107.695 171.450 ;
        RECT 107.430 168.540 107.730 170.840 ;
        RECT 107.465 163.450 107.695 168.540 ;
        RECT 108.755 167.140 108.985 171.450 ;
        RECT 110.045 170.840 110.275 171.450 ;
        RECT 110.010 168.540 110.310 170.840 ;
        RECT 108.720 164.840 109.020 167.140 ;
        RECT 108.755 163.450 108.985 164.840 ;
        RECT 110.045 163.450 110.275 168.540 ;
        RECT 110.685 166.625 114.420 172.070 ;
        RECT 114.920 167.475 115.150 172.070 ;
        RECT 115.710 170.895 115.940 175.475 ;
        RECT 116.500 174.870 116.730 175.475 ;
        RECT 116.465 172.070 116.765 174.870 ;
        RECT 115.675 168.095 115.975 170.895 ;
        RECT 115.710 167.475 115.940 168.095 ;
        RECT 116.500 167.475 116.730 172.070 ;
        RECT 117.290 170.895 117.520 175.475 ;
        RECT 118.080 174.870 118.310 175.475 ;
        RECT 119.540 174.870 119.770 175.475 ;
        RECT 118.045 172.070 118.345 174.870 ;
        RECT 119.505 172.070 119.805 174.870 ;
        RECT 117.255 168.095 117.555 170.895 ;
        RECT 117.290 167.475 117.520 168.095 ;
        RECT 118.080 167.475 118.310 172.070 ;
        RECT 119.540 167.475 119.770 172.070 ;
        RECT 120.330 170.895 120.560 175.475 ;
        RECT 121.120 174.870 121.350 175.475 ;
        RECT 121.085 172.070 121.385 174.870 ;
        RECT 120.295 168.095 120.595 170.895 ;
        RECT 120.330 167.475 120.560 168.095 ;
        RECT 121.120 167.475 121.350 172.070 ;
        RECT 121.910 170.895 122.140 175.475 ;
        RECT 122.700 174.870 122.930 175.475 ;
        RECT 124.160 174.870 124.390 175.475 ;
        RECT 122.665 172.070 122.965 174.870 ;
        RECT 124.125 172.070 124.425 174.870 ;
        RECT 121.875 168.095 122.175 170.895 ;
        RECT 121.910 167.475 122.140 168.095 ;
        RECT 122.700 167.475 122.930 172.070 ;
        RECT 124.160 167.475 124.390 172.070 ;
        RECT 124.950 170.895 125.180 175.475 ;
        RECT 125.740 174.870 125.970 175.475 ;
        RECT 125.705 172.070 126.005 174.870 ;
        RECT 124.915 168.095 125.215 170.895 ;
        RECT 124.950 167.475 125.180 168.095 ;
        RECT 125.740 167.475 125.970 172.070 ;
        RECT 126.530 170.895 126.760 175.475 ;
        RECT 127.320 174.870 127.550 175.475 ;
        RECT 128.780 174.870 129.010 175.475 ;
        RECT 127.285 172.070 127.585 174.870 ;
        RECT 128.745 172.070 129.045 174.870 ;
        RECT 126.495 168.095 126.795 170.895 ;
        RECT 126.530 167.475 126.760 168.095 ;
        RECT 127.320 167.475 127.550 172.070 ;
        RECT 128.780 167.475 129.010 172.070 ;
        RECT 129.570 170.895 129.800 175.475 ;
        RECT 130.360 174.870 130.590 175.475 ;
        RECT 130.325 172.070 130.625 174.870 ;
        RECT 129.535 168.095 129.835 170.895 ;
        RECT 129.570 167.475 129.800 168.095 ;
        RECT 130.360 167.475 130.590 172.070 ;
        RECT 131.150 170.895 131.380 175.475 ;
        RECT 131.940 174.870 132.170 175.475 ;
        RECT 133.400 174.870 133.630 175.475 ;
        RECT 131.905 172.070 132.205 174.870 ;
        RECT 133.365 172.070 133.665 174.870 ;
        RECT 131.115 168.095 131.415 170.895 ;
        RECT 131.150 167.475 131.380 168.095 ;
        RECT 131.940 167.475 132.170 172.070 ;
        RECT 133.400 167.475 133.630 172.070 ;
        RECT 134.190 170.895 134.420 175.475 ;
        RECT 134.980 174.870 135.210 175.475 ;
        RECT 134.945 172.070 135.245 174.870 ;
        RECT 134.155 168.095 134.455 170.895 ;
        RECT 134.190 167.475 134.420 168.095 ;
        RECT 134.980 167.475 135.210 172.070 ;
        RECT 135.770 170.895 136.000 175.475 ;
        RECT 136.560 174.870 136.790 175.475 ;
        RECT 138.020 174.870 138.250 175.475 ;
        RECT 136.525 172.070 136.825 174.870 ;
        RECT 137.985 172.070 138.285 174.870 ;
        RECT 135.735 168.095 136.035 170.895 ;
        RECT 135.770 167.475 136.000 168.095 ;
        RECT 136.560 167.475 136.790 172.070 ;
        RECT 138.020 167.475 138.250 172.070 ;
        RECT 138.810 170.895 139.040 175.475 ;
        RECT 139.600 174.870 139.830 175.475 ;
        RECT 139.565 172.070 139.865 174.870 ;
        RECT 138.775 168.095 139.075 170.895 ;
        RECT 138.810 167.475 139.040 168.095 ;
        RECT 139.600 167.475 139.830 172.070 ;
        RECT 140.390 170.895 140.620 175.475 ;
        RECT 141.180 174.870 141.410 175.475 ;
        RECT 142.640 174.870 142.870 175.475 ;
        RECT 141.145 172.070 141.445 174.870 ;
        RECT 142.605 172.070 142.905 174.870 ;
        RECT 140.355 168.095 140.655 170.895 ;
        RECT 140.390 167.475 140.620 168.095 ;
        RECT 141.180 167.475 141.410 172.070 ;
        RECT 142.640 167.475 142.870 172.070 ;
        RECT 143.430 170.895 143.660 175.475 ;
        RECT 144.220 174.870 144.450 175.475 ;
        RECT 144.185 172.070 144.485 174.870 ;
        RECT 143.395 168.095 143.695 170.895 ;
        RECT 143.430 167.475 143.660 168.095 ;
        RECT 144.220 167.475 144.450 172.070 ;
        RECT 145.010 170.895 145.240 175.475 ;
        RECT 145.800 174.870 146.030 175.475 ;
        RECT 147.260 174.870 147.490 175.475 ;
        RECT 145.765 172.070 146.065 174.870 ;
        RECT 147.225 172.070 147.525 174.870 ;
        RECT 144.975 168.095 145.275 170.895 ;
        RECT 145.010 167.475 145.240 168.095 ;
        RECT 145.800 167.475 146.030 172.070 ;
        RECT 147.260 167.475 147.490 172.070 ;
        RECT 148.050 170.895 148.280 175.475 ;
        RECT 148.840 174.870 149.070 175.475 ;
        RECT 148.805 172.070 149.105 174.870 ;
        RECT 148.015 168.095 148.315 170.895 ;
        RECT 148.050 167.475 148.280 168.095 ;
        RECT 148.840 167.475 149.070 172.070 ;
        RECT 149.630 170.895 149.860 175.475 ;
        RECT 150.420 174.870 150.650 175.475 ;
        RECT 150.385 172.070 150.685 174.870 ;
        RECT 149.595 168.095 149.895 170.895 ;
        RECT 149.630 167.475 149.860 168.095 ;
        RECT 150.420 167.475 150.650 172.070 ;
        RECT 115.200 167.085 115.660 167.315 ;
        RECT 115.990 167.085 116.450 167.315 ;
        RECT 116.780 167.085 117.240 167.315 ;
        RECT 117.570 167.085 118.030 167.315 ;
        RECT 119.820 167.085 120.280 167.315 ;
        RECT 120.610 167.085 121.070 167.315 ;
        RECT 121.400 167.085 121.860 167.315 ;
        RECT 122.190 167.085 122.650 167.315 ;
        RECT 124.440 167.085 124.900 167.315 ;
        RECT 125.230 167.085 125.690 167.315 ;
        RECT 126.020 167.085 126.480 167.315 ;
        RECT 126.810 167.085 127.270 167.315 ;
        RECT 129.060 167.085 129.520 167.315 ;
        RECT 129.850 167.085 130.310 167.315 ;
        RECT 130.640 167.085 131.100 167.315 ;
        RECT 131.430 167.085 131.890 167.315 ;
        RECT 133.680 167.085 134.140 167.315 ;
        RECT 134.470 167.085 134.930 167.315 ;
        RECT 135.260 167.085 135.720 167.315 ;
        RECT 136.050 167.085 136.510 167.315 ;
        RECT 138.300 167.085 138.760 167.315 ;
        RECT 139.090 167.085 139.550 167.315 ;
        RECT 139.880 167.085 140.340 167.315 ;
        RECT 140.670 167.085 141.130 167.315 ;
        RECT 142.920 167.085 143.380 167.315 ;
        RECT 143.710 167.085 144.170 167.315 ;
        RECT 144.500 167.085 144.960 167.315 ;
        RECT 145.290 167.085 145.750 167.315 ;
        RECT 147.540 167.085 148.000 167.315 ;
        RECT 148.330 167.085 148.790 167.315 ;
        RECT 149.120 167.085 149.580 167.315 ;
        RECT 149.910 167.085 150.370 167.315 ;
        RECT 151.150 166.625 152.755 176.325 ;
        RECT 110.685 166.035 152.755 166.625 ;
        RECT 107.745 163.060 108.705 163.290 ;
        RECT 109.035 163.060 109.995 163.290 ;
        RECT 107.745 162.990 108.445 163.060 ;
        RECT 109.295 162.990 109.995 163.060 ;
        RECT 110.685 162.685 114.420 166.035 ;
        RECT 134.745 165.030 135.445 165.080 ;
        RECT 146.905 165.030 147.605 165.080 ;
        RECT 134.745 164.430 147.605 165.030 ;
        RECT 134.745 164.380 135.445 164.430 ;
        RECT 146.905 164.380 147.605 164.430 ;
        RECT 133.735 163.740 134.435 163.790 ;
        RECT 143.985 163.740 144.685 163.790 ;
        RECT 133.735 163.140 144.685 163.740 ;
        RECT 133.735 163.090 134.435 163.140 ;
        RECT 143.985 163.090 144.685 163.140 ;
        RECT 101.935 162.285 114.420 162.685 ;
        RECT 101.935 158.755 103.025 162.285 ;
        RECT 103.435 160.445 103.665 161.520 ;
        RECT 103.400 159.745 103.700 160.445 ;
        RECT 103.435 159.520 103.665 159.745 ;
        RECT 104.725 159.520 104.955 162.285 ;
        RECT 106.015 160.445 106.245 161.520 ;
        RECT 105.980 159.745 106.280 160.445 ;
        RECT 106.015 159.520 106.245 159.745 ;
        RECT 103.715 159.130 104.675 159.360 ;
        RECT 105.005 159.130 105.965 159.360 ;
        RECT 103.845 159.060 104.545 159.130 ;
        RECT 105.135 159.060 105.835 159.130 ;
        RECT 106.655 158.755 107.055 162.285 ;
        RECT 107.465 160.445 107.695 161.520 ;
        RECT 107.430 159.745 107.730 160.445 ;
        RECT 107.465 159.520 107.695 159.745 ;
        RECT 108.755 159.520 108.985 162.285 ;
        RECT 110.045 160.445 110.275 161.520 ;
        RECT 110.010 159.745 110.310 160.445 ;
        RECT 110.045 159.520 110.275 159.745 ;
        RECT 107.745 159.130 108.705 159.360 ;
        RECT 109.035 159.130 109.995 159.360 ;
        RECT 107.875 159.060 108.575 159.130 ;
        RECT 109.165 159.060 109.865 159.130 ;
        RECT 110.685 158.755 114.420 162.285 ;
        RECT 136.825 162.330 137.525 162.400 ;
        RECT 143.985 162.330 144.685 162.400 ;
        RECT 136.825 161.730 144.685 162.330 ;
        RECT 136.825 161.700 137.525 161.730 ;
        RECT 143.985 161.700 144.685 161.730 ;
        RECT 134.745 160.160 135.445 160.210 ;
        RECT 145.575 160.160 146.275 160.210 ;
        RECT 134.745 159.560 146.275 160.160 ;
        RECT 134.745 159.510 135.445 159.560 ;
        RECT 145.575 159.510 146.275 159.560 ;
        RECT 101.935 157.850 114.420 158.755 ;
        RECT 141.665 159.150 142.365 159.200 ;
        RECT 148.605 159.150 149.305 159.200 ;
        RECT 141.665 158.550 149.305 159.150 ;
        RECT 141.665 158.500 142.365 158.550 ;
        RECT 148.605 158.500 149.305 158.550 ;
        RECT 153.960 158.060 155.900 180.110 ;
        RECT 162.095 179.490 236.155 179.970 ;
        RECT 164.480 179.290 164.770 179.335 ;
        RECT 167.225 179.290 167.545 179.350 ;
        RECT 164.480 179.150 167.545 179.290 ;
        RECT 164.480 179.105 164.770 179.150 ;
        RECT 167.225 179.090 167.545 179.150 ;
        RECT 168.145 179.090 168.465 179.350 ;
        RECT 173.665 179.290 173.985 179.350 ;
        RECT 176.440 179.290 176.730 179.335 ;
        RECT 173.665 179.150 176.730 179.290 ;
        RECT 173.665 179.090 173.985 179.150 ;
        RECT 176.440 179.105 176.730 179.150 ;
        RECT 179.200 179.290 179.490 179.335 ;
        RECT 179.645 179.290 179.965 179.350 ;
        RECT 179.200 179.150 179.965 179.290 ;
        RECT 179.200 179.105 179.490 179.150 ;
        RECT 179.645 179.090 179.965 179.150 ;
        RECT 180.580 179.290 180.870 179.335 ;
        RECT 181.025 179.290 181.345 179.350 ;
        RECT 180.580 179.150 181.345 179.290 ;
        RECT 180.580 179.105 180.870 179.150 ;
        RECT 181.025 179.090 181.345 179.150 ;
        RECT 181.945 179.090 182.265 179.350 ;
        RECT 185.165 179.290 185.485 179.350 ;
        RECT 191.620 179.290 191.910 179.335 ;
        RECT 192.065 179.290 192.385 179.350 ;
        RECT 185.165 179.150 190.915 179.290 ;
        RECT 185.165 179.090 185.485 179.150 ;
        RECT 166.780 178.765 167.070 178.995 ;
        RECT 170.460 178.950 170.750 178.995 ;
        RECT 172.745 178.950 173.065 179.010 ;
        RECT 170.460 178.810 173.065 178.950 ;
        RECT 170.460 178.765 170.750 178.810 ;
        RECT 166.855 178.610 166.995 178.765 ;
        RECT 172.745 178.750 173.065 178.810 ;
        RECT 173.220 178.950 173.510 178.995 ;
        RECT 186.545 178.950 186.865 179.010 ;
        RECT 187.480 178.950 187.770 178.995 ;
        RECT 173.220 178.810 186.865 178.950 ;
        RECT 173.220 178.765 173.510 178.810 ;
        RECT 186.545 178.750 186.865 178.810 ;
        RECT 187.095 178.810 187.770 178.950 ;
        RECT 182.405 178.610 182.725 178.670 ;
        RECT 185.640 178.610 185.930 178.655 ;
        RECT 186.085 178.610 186.405 178.670 ;
        RECT 166.855 178.470 174.815 178.610 ;
        RECT 163.545 178.070 163.865 178.330 ;
        RECT 165.845 178.070 166.165 178.330 ;
        RECT 168.605 178.270 168.925 178.330 ;
        RECT 168.410 178.130 168.925 178.270 ;
        RECT 168.605 178.070 168.925 178.130 ;
        RECT 169.065 178.070 169.385 178.330 ;
        RECT 169.525 178.070 169.845 178.330 ;
        RECT 170.920 178.270 171.210 178.315 ;
        RECT 171.365 178.270 171.685 178.330 ;
        RECT 170.920 178.130 171.685 178.270 ;
        RECT 170.920 178.085 171.210 178.130 ;
        RECT 171.365 178.070 171.685 178.130 ;
        RECT 172.300 178.085 172.590 178.315 ;
        RECT 173.205 178.270 173.525 178.330 ;
        RECT 173.680 178.270 173.970 178.315 ;
        RECT 173.205 178.130 173.970 178.270 ;
        RECT 174.675 178.270 174.815 178.470 ;
        RECT 182.405 178.470 186.405 178.610 ;
        RECT 182.405 178.410 182.725 178.470 ;
        RECT 185.640 178.425 185.930 178.470 ;
        RECT 186.085 178.410 186.405 178.470 ;
        RECT 187.095 178.330 187.235 178.810 ;
        RECT 187.480 178.765 187.770 178.810 ;
        RECT 189.765 178.950 190.085 179.010 ;
        RECT 190.240 178.950 190.530 178.995 ;
        RECT 189.765 178.810 190.530 178.950 ;
        RECT 190.775 178.950 190.915 179.150 ;
        RECT 191.620 179.150 192.385 179.290 ;
        RECT 191.620 179.105 191.910 179.150 ;
        RECT 192.065 179.090 192.385 179.150 ;
        RECT 193.000 179.290 193.290 179.335 ;
        RECT 193.445 179.290 193.765 179.350 ;
        RECT 193.000 179.150 193.765 179.290 ;
        RECT 193.000 179.105 193.290 179.150 ;
        RECT 193.445 179.090 193.765 179.150 ;
        RECT 195.745 179.090 196.065 179.350 ;
        RECT 200.805 179.290 201.125 179.350 ;
        RECT 200.805 179.150 214.375 179.290 ;
        RECT 200.805 179.090 201.125 179.150 ;
        RECT 194.365 178.950 194.685 179.010 ;
        RECT 190.775 178.810 194.685 178.950 ;
        RECT 195.835 178.950 195.975 179.090 ;
        RECT 200.360 178.950 200.650 178.995 ;
        RECT 204.485 178.950 204.805 179.010 ;
        RECT 195.835 178.810 200.115 178.950 ;
        RECT 189.765 178.750 190.085 178.810 ;
        RECT 190.240 178.765 190.530 178.810 ;
        RECT 194.365 178.750 194.685 178.810 ;
        RECT 192.525 178.610 192.845 178.670 ;
        RECT 195.760 178.610 196.050 178.655 ;
        RECT 189.395 178.470 196.050 178.610 ;
        RECT 199.975 178.610 200.115 178.810 ;
        RECT 200.360 178.810 204.805 178.950 ;
        RECT 200.360 178.765 200.650 178.810 ;
        RECT 204.485 178.750 204.805 178.810 ;
        RECT 205.830 178.950 206.120 178.995 ;
        RECT 209.060 178.950 209.350 178.995 ;
        RECT 205.830 178.810 209.350 178.950 ;
        RECT 205.830 178.765 206.120 178.810 ;
        RECT 209.060 178.765 209.350 178.810 ;
        RECT 210.005 178.750 210.325 179.010 ;
        RECT 214.235 178.950 214.375 179.150 ;
        RECT 216.445 179.090 216.765 179.350 ;
        RECT 219.665 179.290 219.985 179.350 ;
        RECT 226.120 179.290 226.410 179.335 ;
        RECT 226.565 179.290 226.885 179.350 ;
        RECT 219.665 179.150 225.875 179.290 ;
        RECT 219.665 179.090 219.985 179.150 ;
        RECT 220.140 178.950 220.430 178.995 ;
        RECT 220.585 178.950 220.905 179.010 ;
        RECT 214.235 178.810 218.055 178.950 ;
        RECT 204.040 178.610 204.330 178.655 ;
        RECT 199.975 178.470 204.330 178.610 ;
        RECT 174.675 178.250 175.275 178.270 ;
        RECT 175.520 178.250 175.810 178.315 ;
        RECT 174.675 178.130 175.810 178.250 ;
        RECT 172.375 177.930 172.515 178.085 ;
        RECT 173.205 178.070 173.525 178.130 ;
        RECT 173.680 178.085 173.970 178.130 ;
        RECT 175.135 178.110 175.810 178.130 ;
        RECT 175.520 178.085 175.810 178.110 ;
        RECT 175.965 178.270 176.285 178.330 ;
        RECT 178.280 178.270 178.570 178.315 ;
        RECT 178.725 178.270 179.045 178.330 ;
        RECT 175.965 178.130 176.480 178.270 ;
        RECT 178.280 178.130 179.045 178.270 ;
        RECT 175.965 178.070 176.285 178.130 ;
        RECT 178.280 178.085 178.570 178.130 ;
        RECT 178.725 178.070 179.045 178.130 ;
        RECT 179.645 178.070 179.965 178.330 ;
        RECT 181.040 178.270 181.330 178.315 ;
        RECT 184.720 178.270 185.010 178.315 ;
        RECT 185.165 178.270 185.485 178.330 ;
        RECT 181.040 178.130 184.475 178.270 ;
        RECT 181.040 178.085 181.330 178.130 ;
        RECT 174.125 177.930 174.445 177.990 ;
        RECT 184.335 177.930 184.475 178.130 ;
        RECT 184.720 178.130 185.485 178.270 ;
        RECT 184.720 178.085 185.010 178.130 ;
        RECT 185.165 178.070 185.485 178.130 ;
        RECT 186.560 178.085 186.850 178.315 ;
        RECT 186.635 177.930 186.775 178.085 ;
        RECT 187.005 178.070 187.325 178.330 ;
        RECT 187.925 178.270 188.245 178.330 ;
        RECT 189.395 178.315 189.535 178.470 ;
        RECT 188.400 178.270 188.690 178.315 ;
        RECT 187.925 178.130 188.690 178.270 ;
        RECT 187.925 178.070 188.245 178.130 ;
        RECT 188.400 178.085 188.690 178.130 ;
        RECT 189.170 178.130 189.535 178.315 ;
        RECT 189.170 178.085 189.460 178.130 ;
        RECT 190.685 178.070 191.005 178.330 ;
        RECT 191.695 178.315 191.835 178.470 ;
        RECT 192.525 178.410 192.845 178.470 ;
        RECT 195.760 178.425 196.050 178.470 ;
        RECT 204.040 178.425 204.330 178.470 ;
        RECT 205.405 178.610 205.725 178.670 ;
        RECT 207.245 178.610 207.565 178.670 ;
        RECT 208.165 178.655 208.485 178.670 ;
        RECT 205.405 178.470 207.565 178.610 ;
        RECT 205.405 178.410 205.725 178.470 ;
        RECT 207.245 178.410 207.565 178.470 ;
        RECT 208.055 178.425 208.485 178.655 ;
        RECT 211.845 178.610 212.165 178.670 ;
        RECT 208.165 178.410 208.485 178.425 ;
        RECT 208.715 178.470 212.165 178.610 ;
        RECT 191.470 178.130 191.835 178.315 ;
        RECT 191.470 178.085 191.760 178.130 ;
        RECT 194.825 178.070 195.145 178.330 ;
        RECT 195.300 178.270 195.590 178.315 ;
        RECT 196.205 178.270 196.525 178.330 ;
        RECT 195.300 178.130 196.525 178.270 ;
        RECT 195.300 178.085 195.590 178.130 ;
        RECT 196.205 178.070 196.525 178.130 ;
        RECT 198.060 178.270 198.350 178.315 ;
        RECT 198.965 178.270 199.285 178.330 ;
        RECT 198.060 178.130 199.285 178.270 ;
        RECT 198.060 178.085 198.350 178.130 ;
        RECT 198.965 178.070 199.285 178.130 ;
        RECT 199.440 178.270 199.730 178.315 ;
        RECT 200.345 178.270 200.665 178.330 ;
        RECT 199.440 178.130 200.665 178.270 ;
        RECT 199.440 178.085 199.730 178.130 ;
        RECT 200.345 178.070 200.665 178.130 ;
        RECT 201.265 178.270 201.585 178.330 ;
        RECT 208.715 178.315 208.855 178.470 ;
        RECT 211.845 178.410 212.165 178.470 ;
        RECT 212.305 178.410 212.625 178.670 ;
        RECT 213.225 178.410 213.545 178.670 ;
        RECT 215.065 178.610 215.385 178.670 ;
        RECT 217.915 178.655 218.055 178.810 ;
        RECT 220.140 178.810 220.905 178.950 ;
        RECT 220.140 178.765 220.430 178.810 ;
        RECT 220.585 178.750 220.905 178.810 ;
        RECT 221.100 178.950 221.390 178.995 ;
        RECT 224.330 178.950 224.620 178.995 ;
        RECT 221.100 178.810 224.620 178.950 ;
        RECT 225.735 178.950 225.875 179.150 ;
        RECT 226.120 179.150 226.885 179.290 ;
        RECT 226.120 179.105 226.410 179.150 ;
        RECT 226.565 179.090 226.885 179.150 ;
        RECT 228.420 179.290 228.710 179.335 ;
        RECT 228.865 179.290 229.185 179.350 ;
        RECT 228.420 179.150 229.185 179.290 ;
        RECT 228.420 179.105 228.710 179.150 ;
        RECT 228.865 179.090 229.185 179.150 ;
        RECT 229.325 179.290 229.645 179.350 ;
        RECT 231.180 179.290 231.470 179.335 ;
        RECT 229.325 179.150 231.470 179.290 ;
        RECT 229.325 179.090 229.645 179.150 ;
        RECT 231.180 179.105 231.470 179.150 ;
        RECT 229.800 178.950 230.090 178.995 ;
        RECT 225.735 178.810 230.090 178.950 ;
        RECT 221.100 178.765 221.390 178.810 ;
        RECT 224.330 178.765 224.620 178.810 ;
        RECT 229.800 178.765 230.090 178.810 ;
        RECT 232.560 178.765 232.850 178.995 ;
        RECT 216.920 178.610 217.210 178.655 ;
        RECT 215.065 178.470 217.210 178.610 ;
        RECT 215.065 178.410 215.385 178.470 ;
        RECT 216.920 178.425 217.210 178.470 ;
        RECT 217.840 178.425 218.130 178.655 ;
        RECT 221.505 178.410 221.825 178.670 ;
        RECT 222.210 178.610 222.500 178.655 ;
        RECT 232.635 178.610 232.775 178.765 ;
        RECT 222.210 178.470 232.775 178.610 ;
        RECT 222.210 178.425 222.500 178.470 ;
        RECT 201.740 178.270 202.030 178.315 ;
        RECT 201.265 178.130 202.030 178.270 ;
        RECT 201.265 178.070 201.585 178.130 ;
        RECT 201.740 178.085 202.030 178.130 ;
        RECT 204.910 178.270 205.200 178.315 ;
        RECT 206.750 178.270 207.040 178.315 ;
        RECT 204.910 178.130 207.040 178.270 ;
        RECT 204.910 178.085 205.200 178.130 ;
        RECT 206.750 178.085 207.040 178.130 ;
        RECT 208.640 178.085 208.930 178.315 ;
        RECT 209.095 178.270 209.385 178.315 ;
        RECT 210.935 178.270 211.225 178.315 ;
        RECT 209.095 178.130 211.225 178.270 ;
        RECT 209.095 178.085 209.385 178.130 ;
        RECT 210.935 178.085 211.225 178.130 ;
        RECT 214.160 178.085 214.450 178.315 ;
        RECT 214.605 178.270 214.925 178.330 ;
        RECT 215.540 178.270 215.830 178.315 ;
        RECT 214.605 178.130 215.830 178.270 ;
        RECT 195.745 177.930 196.065 177.990 ;
        RECT 172.375 177.790 174.445 177.930 ;
        RECT 174.125 177.730 174.445 177.790 ;
        RECT 174.675 177.790 183.095 177.930 ;
        RECT 184.335 177.790 186.315 177.930 ;
        RECT 186.635 177.790 196.065 177.930 ;
        RECT 171.840 177.590 172.130 177.635 ;
        RECT 172.285 177.590 172.605 177.650 ;
        RECT 174.675 177.635 174.815 177.790 ;
        RECT 171.840 177.450 172.605 177.590 ;
        RECT 171.840 177.405 172.130 177.450 ;
        RECT 172.285 177.390 172.605 177.450 ;
        RECT 174.600 177.405 174.890 177.635 ;
        RECT 177.805 177.590 178.125 177.650 ;
        RECT 182.420 177.590 182.710 177.635 ;
        RECT 177.805 177.450 182.710 177.590 ;
        RECT 182.955 177.590 183.095 177.790 ;
        RECT 184.260 177.590 184.550 177.635 ;
        RECT 182.955 177.450 184.550 177.590 ;
        RECT 186.175 177.590 186.315 177.790 ;
        RECT 195.745 177.730 196.065 177.790 ;
        RECT 205.415 177.930 205.705 177.975 ;
        RECT 206.335 177.930 206.625 177.975 ;
        RECT 211.855 177.930 212.145 177.975 ;
        RECT 205.415 177.790 212.145 177.930 ;
        RECT 205.415 177.745 205.705 177.790 ;
        RECT 206.335 177.745 206.625 177.790 ;
        RECT 211.855 177.745 212.145 177.790 ;
        RECT 193.905 177.590 194.225 177.650 ;
        RECT 186.175 177.450 194.225 177.590 ;
        RECT 177.805 177.390 178.125 177.450 ;
        RECT 182.420 177.405 182.710 177.450 ;
        RECT 184.260 177.405 184.550 177.450 ;
        RECT 193.905 177.390 194.225 177.450 ;
        RECT 198.980 177.590 199.270 177.635 ;
        RECT 201.725 177.590 202.045 177.650 ;
        RECT 198.980 177.450 202.045 177.590 ;
        RECT 198.980 177.405 199.270 177.450 ;
        RECT 201.725 177.390 202.045 177.450 ;
        RECT 202.645 177.390 202.965 177.650 ;
        RECT 204.945 177.590 205.265 177.650 ;
        RECT 214.235 177.590 214.375 178.085 ;
        RECT 214.605 178.070 214.925 178.130 ;
        RECT 215.540 178.085 215.830 178.130 ;
        RECT 219.225 178.270 219.515 178.315 ;
        RECT 221.065 178.270 221.355 178.315 ;
        RECT 219.225 178.130 221.355 178.270 ;
        RECT 219.225 178.085 219.515 178.130 ;
        RECT 221.065 178.085 221.355 178.130 ;
        RECT 222.885 178.070 223.205 178.330 ;
        RECT 223.410 178.270 223.700 178.315 ;
        RECT 225.250 178.270 225.540 178.315 ;
        RECT 223.410 178.130 225.540 178.270 ;
        RECT 223.410 178.085 223.700 178.130 ;
        RECT 225.250 178.085 225.540 178.130 ;
        RECT 226.565 178.270 226.885 178.330 ;
        RECT 227.960 178.270 228.250 178.315 ;
        RECT 226.565 178.130 228.250 178.270 ;
        RECT 226.565 178.070 226.885 178.130 ;
        RECT 227.960 178.085 228.250 178.130 ;
        RECT 229.325 178.070 229.645 178.330 ;
        RECT 230.705 178.070 231.025 178.330 ;
        RECT 232.085 178.070 232.405 178.330 ;
        RECT 233.465 178.070 233.785 178.330 ;
        RECT 218.305 177.930 218.595 177.975 ;
        RECT 223.825 177.930 224.115 177.975 ;
        RECT 224.745 177.930 225.035 177.975 ;
        RECT 218.305 177.790 225.035 177.930 ;
        RECT 218.305 177.745 218.595 177.790 ;
        RECT 223.825 177.745 224.115 177.790 ;
        RECT 224.745 177.745 225.035 177.790 ;
        RECT 204.945 177.450 214.375 177.590 ;
        RECT 215.080 177.590 215.370 177.635 ;
        RECT 215.525 177.590 215.845 177.650 ;
        RECT 215.080 177.450 215.845 177.590 ;
        RECT 204.945 177.390 205.265 177.450 ;
        RECT 215.080 177.405 215.370 177.450 ;
        RECT 215.525 177.390 215.845 177.450 ;
        RECT 223.345 177.590 223.665 177.650 ;
        RECT 227.040 177.590 227.330 177.635 ;
        RECT 223.345 177.450 227.330 177.590 ;
        RECT 223.345 177.390 223.665 177.450 ;
        RECT 227.040 177.405 227.330 177.450 ;
        RECT 162.095 176.770 236.155 177.250 ;
        RECT 163.085 176.570 163.405 176.630 ;
        RECT 172.285 176.570 172.605 176.630 ;
        RECT 163.085 176.430 172.605 176.570 ;
        RECT 163.085 176.370 163.405 176.430 ;
        RECT 172.285 176.370 172.605 176.430 ;
        RECT 180.565 176.370 180.885 176.630 ;
        RECT 187.005 176.570 187.325 176.630 ;
        RECT 198.045 176.570 198.365 176.630 ;
        RECT 187.005 176.430 198.365 176.570 ;
        RECT 187.005 176.370 187.325 176.430 ;
        RECT 198.045 176.370 198.365 176.430 ;
        RECT 202.645 176.570 202.965 176.630 ;
        RECT 212.765 176.570 213.085 176.630 ;
        RECT 202.645 176.430 213.085 176.570 ;
        RECT 202.645 176.370 202.965 176.430 ;
        RECT 212.765 176.370 213.085 176.430 ;
        RECT 219.205 176.570 219.525 176.630 ;
        RECT 232.085 176.570 232.405 176.630 ;
        RECT 219.205 176.430 232.405 176.570 ;
        RECT 219.205 176.370 219.525 176.430 ;
        RECT 232.085 176.370 232.405 176.430 ;
        RECT 171.365 176.230 171.685 176.290 ;
        RECT 180.655 176.230 180.795 176.370 ;
        RECT 171.365 176.090 180.795 176.230 ;
        RECT 206.325 176.230 206.645 176.290 ;
        RECT 214.605 176.230 214.925 176.290 ;
        RECT 206.325 176.090 214.925 176.230 ;
        RECT 171.365 176.030 171.685 176.090 ;
        RECT 206.325 176.030 206.645 176.090 ;
        RECT 214.605 176.030 214.925 176.090 ;
        RECT 218.285 176.230 218.605 176.290 ;
        RECT 233.465 176.230 233.785 176.290 ;
        RECT 218.285 176.090 233.785 176.230 ;
        RECT 218.285 176.030 218.605 176.090 ;
        RECT 233.465 176.030 233.785 176.090 ;
        RECT 174.125 175.890 174.445 175.950 ;
        RECT 184.245 175.890 184.565 175.950 ;
        RECT 174.125 175.750 184.565 175.890 ;
        RECT 174.125 175.690 174.445 175.750 ;
        RECT 184.245 175.690 184.565 175.750 ;
        RECT 216.445 175.890 216.765 175.950 ;
        RECT 230.705 175.890 231.025 175.950 ;
        RECT 216.445 175.750 231.025 175.890 ;
        RECT 216.445 175.690 216.765 175.750 ;
        RECT 230.705 175.690 231.025 175.750 ;
        RECT 165.845 175.550 166.165 175.610 ;
        RECT 177.805 175.550 178.125 175.610 ;
        RECT 165.845 175.410 178.125 175.550 ;
        RECT 165.845 175.350 166.165 175.410 ;
        RECT 177.805 175.350 178.125 175.410 ;
        RECT 179.645 175.550 179.965 175.610 ;
        RECT 191.605 175.550 191.925 175.610 ;
        RECT 179.645 175.410 191.925 175.550 ;
        RECT 179.645 175.350 179.965 175.410 ;
        RECT 191.605 175.350 191.925 175.410 ;
        RECT 215.525 175.550 215.845 175.610 ;
        RECT 229.325 175.550 229.645 175.610 ;
        RECT 215.525 175.410 229.645 175.550 ;
        RECT 215.525 175.350 215.845 175.410 ;
        RECT 229.325 175.350 229.645 175.410 ;
        RECT 167.685 175.210 168.005 175.270 ;
        RECT 175.045 175.210 175.365 175.270 ;
        RECT 167.685 175.070 175.365 175.210 ;
        RECT 167.685 175.010 168.005 175.070 ;
        RECT 175.045 175.010 175.365 175.070 ;
        RECT 178.725 175.210 179.045 175.270 ;
        RECT 190.685 175.210 191.005 175.270 ;
        RECT 178.725 175.070 191.005 175.210 ;
        RECT 178.725 175.010 179.045 175.070 ;
        RECT 190.685 175.010 191.005 175.070 ;
        RECT 213.685 175.210 214.005 175.270 ;
        RECT 226.565 175.210 226.885 175.270 ;
        RECT 213.685 175.070 226.885 175.210 ;
        RECT 213.685 175.010 214.005 175.070 ;
        RECT 226.565 175.010 226.885 175.070 ;
        RECT 221.045 174.870 221.365 174.930 ;
        RECT 231.625 174.870 231.945 174.930 ;
        RECT 221.045 174.730 231.945 174.870 ;
        RECT 221.045 174.670 221.365 174.730 ;
        RECT 231.625 174.670 231.945 174.730 ;
        RECT 173.205 174.530 173.525 174.590 ;
        RECT 185.165 174.530 185.485 174.590 ;
        RECT 173.205 174.390 185.485 174.530 ;
        RECT 173.205 174.330 173.525 174.390 ;
        RECT 185.165 174.330 185.485 174.390 ;
        RECT 207.245 174.530 207.565 174.590 ;
        RECT 210.925 174.530 211.245 174.590 ;
        RECT 207.245 174.390 211.245 174.530 ;
        RECT 207.245 174.330 207.565 174.390 ;
        RECT 210.925 174.330 211.245 174.390 ;
        RECT 115.985 156.185 155.900 158.060 ;
        RECT 115.985 156.060 116.575 156.185 ;
        RECT 102.625 155.660 116.575 156.060 ;
        RECT 102.625 152.040 103.025 155.660 ;
        RECT 103.715 155.055 104.675 155.385 ;
        RECT 105.005 155.055 105.965 155.385 ;
        RECT 103.435 153.515 103.665 154.850 ;
        RECT 103.400 152.815 103.700 153.515 ;
        RECT 104.725 152.040 104.955 154.850 ;
        RECT 106.015 154.585 106.245 154.850 ;
        RECT 105.980 153.885 106.280 154.585 ;
        RECT 106.015 152.850 106.245 153.885 ;
        RECT 106.655 152.040 107.055 155.660 ;
        RECT 107.745 155.055 108.705 155.385 ;
        RECT 109.035 155.055 109.995 155.385 ;
        RECT 107.465 153.515 107.695 154.850 ;
        RECT 107.430 152.815 107.730 153.515 ;
        RECT 108.755 152.040 108.985 154.850 ;
        RECT 110.045 154.585 110.275 154.850 ;
        RECT 110.010 153.885 110.310 154.585 ;
        RECT 110.045 152.850 110.275 153.885 ;
        RECT 110.685 152.040 116.575 155.660 ;
        RECT 102.625 151.550 116.575 152.040 ;
        RECT 102.625 142.020 103.025 151.550 ;
        RECT 103.715 151.035 104.675 151.365 ;
        RECT 105.005 151.035 105.965 151.365 ;
        RECT 103.435 145.785 103.665 150.830 ;
        RECT 104.725 149.485 104.955 150.830 ;
        RECT 104.690 147.185 104.990 149.485 ;
        RECT 103.400 143.485 103.700 145.785 ;
        RECT 103.435 142.830 103.665 143.485 ;
        RECT 104.725 142.830 104.955 147.185 ;
        RECT 106.015 145.785 106.245 150.830 ;
        RECT 105.980 143.485 106.280 145.785 ;
        RECT 106.015 142.830 106.245 143.485 ;
        RECT 103.715 142.395 104.675 142.625 ;
        RECT 105.005 142.395 105.965 142.625 ;
        RECT 106.655 142.020 107.055 151.550 ;
        RECT 107.745 151.035 108.705 151.365 ;
        RECT 109.035 151.035 109.995 151.365 ;
        RECT 107.465 145.785 107.695 150.830 ;
        RECT 108.755 149.485 108.985 150.830 ;
        RECT 108.720 147.185 109.020 149.485 ;
        RECT 107.430 143.485 107.730 145.785 ;
        RECT 107.465 142.830 107.695 143.485 ;
        RECT 108.755 142.830 108.985 147.185 ;
        RECT 110.045 145.785 110.275 150.830 ;
        RECT 110.010 143.485 110.310 145.785 ;
        RECT 110.045 142.830 110.275 143.485 ;
        RECT 107.745 142.395 108.705 142.625 ;
        RECT 109.035 142.395 109.995 142.625 ;
        RECT 110.685 142.020 116.575 151.550 ;
        RECT 117.160 142.145 119.265 155.605 ;
        RECT 122.405 146.245 124.510 155.605 ;
        RECT 125.090 146.825 127.195 155.605 ;
        RECT 130.335 146.825 132.440 155.605 ;
        RECT 133.020 154.960 135.125 155.660 ;
        RECT 133.020 152.675 135.125 154.435 ;
        RECT 138.265 153.845 140.370 155.605 ;
        RECT 133.020 151.450 135.125 152.150 ;
        RECT 138.265 151.505 140.370 153.265 ;
        RECT 140.950 152.675 143.055 156.185 ;
        RECT 146.195 152.675 148.300 156.185 ;
        RECT 140.950 151.460 143.055 152.160 ;
        RECT 133.020 150.280 135.125 150.980 ;
        RECT 133.020 149.110 135.125 149.810 ;
        RECT 138.265 149.165 140.370 150.925 ;
        RECT 140.950 149.165 143.055 150.925 ;
        RECT 146.195 150.335 148.300 152.095 ;
        RECT 133.020 146.825 135.125 148.585 ;
        RECT 138.265 146.825 140.370 148.585 ;
        RECT 140.950 146.825 143.055 148.585 ;
        RECT 146.195 147.995 148.300 149.755 ;
        RECT 122.405 142.145 127.195 146.245 ;
        RECT 130.335 142.145 132.440 146.245 ;
        RECT 133.020 142.145 135.125 146.245 ;
        RECT 138.265 142.145 140.370 146.245 ;
        RECT 140.950 144.485 143.055 146.245 ;
        RECT 146.195 145.655 148.300 147.415 ;
        RECT 140.950 143.290 143.055 143.990 ;
        RECT 146.195 143.315 148.300 145.075 ;
        RECT 140.950 142.040 143.055 142.740 ;
        RECT 146.195 142.080 148.300 142.780 ;
        RECT 102.625 141.620 116.575 142.020 ;
        RECT 62.865 130.990 100.480 139.455 ;
        RECT 111.085 141.565 116.575 141.620 ;
        RECT 148.885 141.565 155.900 156.185 ;
        RECT 111.085 137.690 155.900 141.565 ;
        RECT 111.085 130.990 135.120 137.690 ;
        RECT 62.865 127.485 135.120 130.990 ;
        RECT 138.080 134.100 145.960 137.690 ;
        RECT 138.080 130.310 138.670 134.100 ;
        RECT 139.615 133.640 140.315 133.760 ;
        RECT 140.905 133.640 141.605 133.760 ;
        RECT 139.485 133.410 140.445 133.640 ;
        RECT 140.775 133.410 141.735 133.640 ;
        RECT 139.205 132.990 139.435 133.205 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 139.205 131.205 139.435 131.390 ;
        RECT 140.495 130.310 140.725 133.205 ;
        RECT 141.785 132.990 142.015 133.205 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 143.315 132.640 143.545 133.205 ;
        RECT 143.280 131.940 143.580 132.640 ;
        RECT 141.785 131.205 142.015 131.390 ;
        RECT 143.315 131.205 143.545 131.940 ;
        RECT 144.605 131.205 144.835 134.100 ;
        RECT 143.595 130.770 144.555 131.000 ;
        RECT 143.725 130.700 144.425 130.770 ;
        RECT 145.370 130.310 145.960 134.100 ;
        RECT 138.080 129.720 145.960 130.310 ;
        RECT 4.100 124.285 135.120 127.485 ;
        RECT 4.100 44.835 4.900 124.285 ;
        RECT 8.665 123.695 70.175 124.285 ;
        RECT 8.665 122.800 10.615 123.695 ;
        RECT 11.335 123.005 13.295 123.235 ;
        RECT 13.625 123.005 15.585 123.235 ;
        RECT 17.255 123.005 19.215 123.305 ;
        RECT 19.545 123.005 21.505 123.305 ;
        RECT 23.175 123.005 25.135 123.305 ;
        RECT 25.465 123.005 27.425 123.305 ;
        RECT 29.095 123.005 31.055 123.305 ;
        RECT 31.385 123.005 33.345 123.305 ;
        RECT 35.015 123.005 36.975 123.305 ;
        RECT 37.305 123.005 39.265 123.305 ;
        RECT 40.935 123.005 42.895 123.305 ;
        RECT 43.225 123.005 45.185 123.305 ;
        RECT 46.855 123.005 48.815 123.305 ;
        RECT 49.145 123.005 51.105 123.305 ;
        RECT 52.775 123.005 54.735 123.305 ;
        RECT 55.065 123.005 57.025 123.305 ;
        RECT 58.695 123.005 60.655 123.305 ;
        RECT 60.985 123.005 62.945 123.305 ;
        RECT 64.615 123.005 66.575 123.235 ;
        RECT 66.905 123.005 68.865 123.235 ;
        RECT 69.585 122.800 70.175 123.695 ;
        RECT 8.665 117.050 11.285 122.800 ;
        RECT 13.345 117.050 13.575 122.800 ;
        RECT 15.635 117.050 15.865 122.800 ;
        RECT 16.975 117.050 17.205 122.800 ;
        RECT 19.265 122.050 19.495 122.800 ;
        RECT 19.030 120.550 19.730 122.050 ;
        RECT 8.665 115.550 11.520 117.050 ;
        RECT 13.110 115.550 13.810 117.050 ;
        RECT 15.400 115.550 16.100 117.050 ;
        RECT 16.740 115.550 17.440 117.050 ;
        RECT 8.665 114.595 11.285 115.550 ;
        RECT 13.345 114.595 13.575 115.550 ;
        RECT 15.635 114.595 15.865 115.550 ;
        RECT 16.975 114.800 17.205 115.550 ;
        RECT 19.265 114.800 19.495 120.550 ;
        RECT 21.555 117.050 21.785 122.800 ;
        RECT 22.895 117.050 23.125 122.800 ;
        RECT 25.185 119.550 25.415 122.800 ;
        RECT 24.950 118.050 25.650 119.550 ;
        RECT 21.320 115.550 22.020 117.050 ;
        RECT 22.660 115.550 23.360 117.050 ;
        RECT 21.555 114.800 21.785 115.550 ;
        RECT 22.895 114.800 23.125 115.550 ;
        RECT 25.185 114.800 25.415 118.050 ;
        RECT 27.475 117.050 27.705 122.800 ;
        RECT 28.815 117.050 29.045 122.800 ;
        RECT 27.240 115.550 27.940 117.050 ;
        RECT 28.580 115.550 29.280 117.050 ;
        RECT 27.475 114.800 27.705 115.550 ;
        RECT 28.815 114.800 29.045 115.550 ;
        RECT 31.105 114.595 31.335 122.800 ;
        RECT 33.395 117.050 33.625 122.800 ;
        RECT 34.735 117.050 34.965 122.800 ;
        RECT 37.025 122.050 37.255 122.800 ;
        RECT 36.790 120.550 37.490 122.050 ;
        RECT 33.160 115.550 33.860 117.050 ;
        RECT 34.500 115.550 35.200 117.050 ;
        RECT 33.395 114.800 33.625 115.550 ;
        RECT 34.735 114.800 34.965 115.550 ;
        RECT 37.025 114.800 37.255 120.550 ;
        RECT 39.315 117.050 39.545 122.800 ;
        RECT 40.655 117.050 40.885 122.800 ;
        RECT 42.945 122.050 43.175 122.800 ;
        RECT 42.710 120.550 43.410 122.050 ;
        RECT 39.080 115.550 39.780 117.050 ;
        RECT 40.420 115.550 41.120 117.050 ;
        RECT 39.315 114.800 39.545 115.550 ;
        RECT 40.655 114.800 40.885 115.550 ;
        RECT 42.945 114.800 43.175 120.550 ;
        RECT 45.235 117.050 45.465 122.800 ;
        RECT 46.575 117.050 46.805 122.800 ;
        RECT 45.000 115.550 45.700 117.050 ;
        RECT 46.340 115.550 47.040 117.050 ;
        RECT 45.235 114.800 45.465 115.550 ;
        RECT 46.575 114.800 46.805 115.550 ;
        RECT 48.865 114.595 49.095 122.800 ;
        RECT 51.155 117.050 51.385 122.800 ;
        RECT 52.495 117.050 52.725 122.800 ;
        RECT 54.785 119.550 55.015 122.800 ;
        RECT 54.550 118.050 55.250 119.550 ;
        RECT 50.920 115.550 51.620 117.050 ;
        RECT 52.260 115.550 52.960 117.050 ;
        RECT 51.155 114.800 51.385 115.550 ;
        RECT 52.495 114.800 52.725 115.550 ;
        RECT 54.785 114.800 55.015 118.050 ;
        RECT 57.075 117.050 57.305 122.800 ;
        RECT 58.415 117.050 58.645 122.800 ;
        RECT 60.705 122.050 60.935 122.800 ;
        RECT 60.470 120.550 61.170 122.050 ;
        RECT 56.840 115.550 57.540 117.050 ;
        RECT 58.180 115.550 58.880 117.050 ;
        RECT 57.075 114.800 57.305 115.550 ;
        RECT 58.415 114.800 58.645 115.550 ;
        RECT 60.705 114.800 60.935 120.550 ;
        RECT 62.995 117.050 63.225 122.800 ;
        RECT 64.335 117.050 64.565 122.800 ;
        RECT 66.625 117.050 66.855 122.800 ;
        RECT 68.915 117.050 70.175 122.800 ;
        RECT 62.760 115.550 63.460 117.050 ;
        RECT 64.100 115.550 64.800 117.050 ;
        RECT 66.390 115.550 67.090 117.050 ;
        RECT 68.680 115.550 70.175 117.050 ;
        RECT 62.995 114.800 63.225 115.550 ;
        RECT 64.335 114.595 64.565 115.550 ;
        RECT 66.625 114.595 66.855 115.550 ;
        RECT 68.915 114.595 70.175 115.550 ;
        RECT 8.665 114.365 15.865 114.595 ;
        RECT 8.665 113.215 10.615 114.365 ;
        RECT 17.255 114.295 19.215 114.595 ;
        RECT 19.545 114.295 21.505 114.595 ;
        RECT 23.175 114.295 25.135 114.595 ;
        RECT 25.465 114.295 27.425 114.595 ;
        RECT 29.095 114.365 33.345 114.595 ;
        RECT 29.095 114.295 31.055 114.365 ;
        RECT 31.385 114.295 33.345 114.365 ;
        RECT 35.015 114.295 36.975 114.595 ;
        RECT 37.305 114.295 39.265 114.595 ;
        RECT 40.935 114.295 42.895 114.595 ;
        RECT 43.225 114.295 45.185 114.595 ;
        RECT 46.855 114.365 51.105 114.595 ;
        RECT 46.855 114.295 48.815 114.365 ;
        RECT 49.145 114.295 51.105 114.365 ;
        RECT 52.775 114.295 54.735 114.595 ;
        RECT 55.065 114.295 57.025 114.595 ;
        RECT 58.695 114.295 60.655 114.595 ;
        RECT 60.985 114.295 62.945 114.595 ;
        RECT 64.335 114.365 70.175 114.595 ;
        RECT 8.665 112.985 15.865 113.215 ;
        RECT 17.255 112.985 19.215 113.285 ;
        RECT 19.545 112.985 21.505 113.285 ;
        RECT 23.175 112.985 25.135 113.285 ;
        RECT 25.465 112.985 27.425 113.285 ;
        RECT 29.095 113.215 31.055 113.285 ;
        RECT 31.385 113.215 33.345 113.285 ;
        RECT 29.095 112.985 33.345 113.215 ;
        RECT 35.015 112.985 36.975 113.285 ;
        RECT 37.305 112.985 39.265 113.285 ;
        RECT 40.935 112.985 42.895 113.285 ;
        RECT 43.225 112.985 45.185 113.285 ;
        RECT 46.855 113.215 48.815 113.285 ;
        RECT 49.145 113.215 51.105 113.285 ;
        RECT 46.855 112.985 51.105 113.215 ;
        RECT 52.775 112.985 54.735 113.285 ;
        RECT 55.065 112.985 57.025 113.285 ;
        RECT 58.695 112.985 60.655 113.285 ;
        RECT 60.985 112.985 62.945 113.285 ;
        RECT 69.585 113.215 70.175 114.365 ;
        RECT 64.335 112.985 70.175 113.215 ;
        RECT 8.665 112.030 11.285 112.985 ;
        RECT 13.345 112.030 13.575 112.985 ;
        RECT 15.635 112.030 15.865 112.985 ;
        RECT 16.975 112.030 17.205 112.780 ;
        RECT 8.665 110.530 11.520 112.030 ;
        RECT 13.110 110.530 13.810 112.030 ;
        RECT 15.400 110.530 16.100 112.030 ;
        RECT 16.740 110.530 17.440 112.030 ;
        RECT 8.665 104.780 11.285 110.530 ;
        RECT 13.345 104.780 13.575 110.530 ;
        RECT 15.635 104.780 15.865 110.530 ;
        RECT 16.975 104.780 17.205 110.530 ;
        RECT 19.265 107.030 19.495 112.780 ;
        RECT 21.555 112.030 21.785 112.780 ;
        RECT 22.895 112.030 23.125 112.780 ;
        RECT 21.320 110.530 22.020 112.030 ;
        RECT 22.660 110.530 23.360 112.030 ;
        RECT 19.030 105.530 19.730 107.030 ;
        RECT 19.265 104.780 19.495 105.530 ;
        RECT 21.555 104.780 21.785 110.530 ;
        RECT 22.895 104.780 23.125 110.530 ;
        RECT 25.185 109.530 25.415 112.780 ;
        RECT 27.475 112.030 27.705 112.780 ;
        RECT 28.815 112.030 29.045 112.780 ;
        RECT 27.240 110.530 27.940 112.030 ;
        RECT 28.580 110.530 29.280 112.030 ;
        RECT 24.950 108.030 25.650 109.530 ;
        RECT 25.185 104.780 25.415 108.030 ;
        RECT 27.475 104.780 27.705 110.530 ;
        RECT 28.815 104.780 29.045 110.530 ;
        RECT 31.105 104.780 31.335 112.985 ;
        RECT 33.395 112.030 33.625 112.780 ;
        RECT 34.735 112.030 34.965 112.780 ;
        RECT 33.160 110.530 33.860 112.030 ;
        RECT 34.500 110.530 35.200 112.030 ;
        RECT 33.395 104.780 33.625 110.530 ;
        RECT 34.735 104.780 34.965 110.530 ;
        RECT 37.025 107.030 37.255 112.780 ;
        RECT 39.315 112.030 39.545 112.780 ;
        RECT 40.655 112.030 40.885 112.780 ;
        RECT 39.080 110.530 39.780 112.030 ;
        RECT 40.420 110.530 41.120 112.030 ;
        RECT 36.790 105.530 37.490 107.030 ;
        RECT 37.025 104.780 37.255 105.530 ;
        RECT 39.315 104.780 39.545 110.530 ;
        RECT 40.655 104.780 40.885 110.530 ;
        RECT 42.945 107.030 43.175 112.780 ;
        RECT 45.235 112.030 45.465 112.780 ;
        RECT 46.575 112.030 46.805 112.780 ;
        RECT 45.000 110.530 45.700 112.030 ;
        RECT 46.340 110.530 47.040 112.030 ;
        RECT 42.710 105.530 43.410 107.030 ;
        RECT 42.945 104.780 43.175 105.530 ;
        RECT 45.235 104.780 45.465 110.530 ;
        RECT 46.575 104.780 46.805 110.530 ;
        RECT 48.865 104.780 49.095 112.985 ;
        RECT 51.155 112.030 51.385 112.780 ;
        RECT 52.495 112.030 52.725 112.780 ;
        RECT 50.920 110.530 51.620 112.030 ;
        RECT 52.260 110.530 52.960 112.030 ;
        RECT 51.155 104.780 51.385 110.530 ;
        RECT 52.495 104.780 52.725 110.530 ;
        RECT 54.785 109.530 55.015 112.780 ;
        RECT 57.075 112.030 57.305 112.780 ;
        RECT 58.415 112.030 58.645 112.780 ;
        RECT 56.840 110.530 57.540 112.030 ;
        RECT 58.180 110.530 58.880 112.030 ;
        RECT 54.550 108.030 55.250 109.530 ;
        RECT 54.785 104.780 55.015 108.030 ;
        RECT 57.075 104.780 57.305 110.530 ;
        RECT 58.415 104.780 58.645 110.530 ;
        RECT 60.705 107.030 60.935 112.780 ;
        RECT 62.995 112.030 63.225 112.780 ;
        RECT 64.335 112.030 64.565 112.985 ;
        RECT 66.625 112.030 66.855 112.985 ;
        RECT 68.915 112.030 70.175 112.985 ;
        RECT 62.760 110.530 63.460 112.030 ;
        RECT 64.100 110.530 64.800 112.030 ;
        RECT 66.390 110.530 67.090 112.030 ;
        RECT 68.680 110.530 70.175 112.030 ;
        RECT 60.470 105.530 61.170 107.030 ;
        RECT 60.705 104.780 60.935 105.530 ;
        RECT 62.995 104.780 63.225 110.530 ;
        RECT 64.335 104.780 64.565 110.530 ;
        RECT 66.625 104.780 66.855 110.530 ;
        RECT 68.915 104.780 70.175 110.530 ;
        RECT 8.665 103.885 10.615 104.780 ;
        RECT 11.335 104.345 13.295 104.575 ;
        RECT 13.625 104.345 15.585 104.575 ;
        RECT 17.255 104.275 19.215 104.575 ;
        RECT 19.545 104.275 21.505 104.575 ;
        RECT 23.175 104.275 25.135 104.575 ;
        RECT 25.465 104.275 27.425 104.575 ;
        RECT 29.095 104.275 31.055 104.575 ;
        RECT 31.385 104.275 33.345 104.575 ;
        RECT 35.015 104.275 36.975 104.575 ;
        RECT 37.305 104.275 39.265 104.575 ;
        RECT 40.935 104.275 42.895 104.575 ;
        RECT 43.225 104.275 45.185 104.575 ;
        RECT 46.855 104.275 48.815 104.575 ;
        RECT 49.145 104.275 51.105 104.575 ;
        RECT 52.775 104.275 54.735 104.575 ;
        RECT 55.065 104.275 57.025 104.575 ;
        RECT 58.695 104.275 60.655 104.575 ;
        RECT 60.985 104.275 62.945 104.575 ;
        RECT 64.615 104.345 66.575 104.575 ;
        RECT 66.905 104.345 68.865 104.575 ;
        RECT 69.585 103.885 70.175 104.780 ;
        RECT 8.665 102.705 70.175 103.885 ;
        RECT 71.775 123.695 114.165 124.285 ;
        RECT 71.775 103.885 72.365 123.695 ;
        RECT 72.805 122.800 77.615 123.695 ;
        RECT 79.005 123.005 80.965 123.305 ;
        RECT 81.295 123.005 83.255 123.305 ;
        RECT 84.925 123.005 86.885 123.305 ;
        RECT 87.215 123.005 89.175 123.305 ;
        RECT 90.845 123.005 95.095 123.305 ;
        RECT 96.765 123.005 98.725 123.305 ;
        RECT 99.055 123.005 101.015 123.305 ;
        RECT 102.685 123.005 104.645 123.305 ;
        RECT 104.975 123.005 106.935 123.305 ;
        RECT 72.805 114.800 73.035 122.800 ;
        RECT 75.095 114.800 75.325 122.800 ;
        RECT 77.385 114.800 77.615 122.800 ;
        RECT 78.725 120.650 78.955 122.800 ;
        RECT 78.490 119.950 79.190 120.650 ;
        RECT 78.725 114.800 78.955 119.950 ;
        RECT 81.015 119.150 81.245 122.800 ;
        RECT 83.305 120.650 83.535 122.800 ;
        RECT 83.070 119.950 83.770 120.650 ;
        RECT 80.780 118.450 81.480 119.150 ;
        RECT 81.015 114.800 81.245 118.450 ;
        RECT 83.305 114.800 83.535 119.950 ;
        RECT 84.645 116.150 84.875 122.800 ;
        RECT 86.935 117.650 87.165 122.800 ;
        RECT 86.700 116.950 87.400 117.650 ;
        RECT 84.410 115.450 85.110 116.150 ;
        RECT 84.645 114.800 84.875 115.450 ;
        RECT 86.935 114.800 87.165 116.950 ;
        RECT 89.225 116.150 89.455 122.800 ;
        RECT 90.565 122.150 90.795 122.800 ;
        RECT 90.330 121.450 91.030 122.150 ;
        RECT 88.990 115.450 89.690 116.150 ;
        RECT 89.225 114.800 89.455 115.450 ;
        RECT 90.565 114.800 90.795 121.450 ;
        RECT 92.855 114.800 93.085 123.005 ;
        RECT 108.325 122.800 113.135 123.695 ;
        RECT 95.145 122.150 95.375 122.800 ;
        RECT 94.910 121.450 95.610 122.150 ;
        RECT 95.145 114.800 95.375 121.450 ;
        RECT 96.485 116.150 96.715 122.800 ;
        RECT 98.775 117.650 99.005 122.800 ;
        RECT 98.540 116.950 99.240 117.650 ;
        RECT 96.250 115.450 96.950 116.150 ;
        RECT 96.485 114.800 96.715 115.450 ;
        RECT 98.775 114.800 99.005 116.950 ;
        RECT 101.065 116.150 101.295 122.800 ;
        RECT 102.405 120.650 102.635 122.800 ;
        RECT 102.170 119.950 102.870 120.650 ;
        RECT 100.830 115.450 101.530 116.150 ;
        RECT 101.065 114.800 101.295 115.450 ;
        RECT 102.405 114.800 102.635 119.950 ;
        RECT 104.695 119.150 104.925 122.800 ;
        RECT 106.985 120.650 107.215 122.800 ;
        RECT 106.750 119.950 107.450 120.650 ;
        RECT 104.460 118.450 105.160 119.150 ;
        RECT 104.695 114.800 104.925 118.450 ;
        RECT 106.985 114.800 107.215 119.950 ;
        RECT 108.325 114.800 108.555 122.800 ;
        RECT 110.615 114.800 110.845 122.800 ;
        RECT 112.905 114.800 113.135 122.800 ;
        RECT 73.085 114.365 75.045 114.595 ;
        RECT 75.375 114.365 77.335 114.595 ;
        RECT 79.005 114.295 80.965 114.595 ;
        RECT 81.295 114.295 83.255 114.595 ;
        RECT 84.925 114.295 86.885 114.595 ;
        RECT 87.215 114.295 89.175 114.595 ;
        RECT 90.845 114.295 92.805 114.595 ;
        RECT 93.135 114.295 95.095 114.595 ;
        RECT 96.765 114.295 98.725 114.595 ;
        RECT 99.055 114.295 101.015 114.595 ;
        RECT 102.685 114.295 104.645 114.595 ;
        RECT 104.975 114.295 106.935 114.595 ;
        RECT 108.605 114.365 110.565 114.595 ;
        RECT 110.895 114.365 112.855 114.595 ;
        RECT 73.085 112.985 75.045 113.215 ;
        RECT 75.375 112.985 77.335 113.215 ;
        RECT 79.005 112.985 80.965 113.285 ;
        RECT 81.295 112.985 83.255 113.285 ;
        RECT 84.925 112.985 86.885 113.285 ;
        RECT 87.215 112.985 89.175 113.285 ;
        RECT 90.845 112.985 92.805 113.285 ;
        RECT 93.135 112.985 95.095 113.285 ;
        RECT 96.765 112.985 98.725 113.285 ;
        RECT 99.055 112.985 101.015 113.285 ;
        RECT 102.685 112.985 104.645 113.285 ;
        RECT 104.975 112.985 106.935 113.285 ;
        RECT 108.605 112.985 110.565 113.215 ;
        RECT 110.895 112.985 112.855 113.215 ;
        RECT 72.805 104.780 73.035 112.780 ;
        RECT 75.095 104.780 75.325 112.780 ;
        RECT 77.385 104.780 77.615 112.780 ;
        RECT 78.725 107.630 78.955 112.780 ;
        RECT 81.015 109.130 81.245 112.780 ;
        RECT 80.780 108.430 81.480 109.130 ;
        RECT 78.490 106.930 79.190 107.630 ;
        RECT 78.725 104.780 78.955 106.930 ;
        RECT 81.015 104.780 81.245 108.430 ;
        RECT 83.305 107.630 83.535 112.780 ;
        RECT 84.645 112.130 84.875 112.780 ;
        RECT 84.410 111.430 85.110 112.130 ;
        RECT 83.070 106.930 83.770 107.630 ;
        RECT 83.305 104.780 83.535 106.930 ;
        RECT 84.645 104.780 84.875 111.430 ;
        RECT 86.935 110.630 87.165 112.780 ;
        RECT 89.225 112.130 89.455 112.780 ;
        RECT 88.990 111.430 89.690 112.130 ;
        RECT 86.700 109.930 87.400 110.630 ;
        RECT 86.935 104.780 87.165 109.930 ;
        RECT 89.225 104.780 89.455 111.430 ;
        RECT 90.565 106.130 90.795 112.780 ;
        RECT 90.330 105.430 91.030 106.130 ;
        RECT 90.565 104.780 90.795 105.430 ;
        RECT 72.805 103.885 77.615 104.780 ;
        RECT 92.855 104.575 93.085 112.780 ;
        RECT 95.145 106.130 95.375 112.780 ;
        RECT 96.485 112.130 96.715 112.780 ;
        RECT 96.250 111.430 96.950 112.130 ;
        RECT 94.910 105.430 95.610 106.130 ;
        RECT 95.145 104.780 95.375 105.430 ;
        RECT 96.485 104.780 96.715 111.430 ;
        RECT 98.775 110.630 99.005 112.780 ;
        RECT 101.065 112.130 101.295 112.780 ;
        RECT 100.830 111.430 101.530 112.130 ;
        RECT 98.540 109.930 99.240 110.630 ;
        RECT 98.775 104.780 99.005 109.930 ;
        RECT 101.065 104.780 101.295 111.430 ;
        RECT 102.405 107.630 102.635 112.780 ;
        RECT 104.695 109.130 104.925 112.780 ;
        RECT 104.460 108.430 105.160 109.130 ;
        RECT 102.170 106.930 102.870 107.630 ;
        RECT 102.405 104.780 102.635 106.930 ;
        RECT 104.695 104.780 104.925 108.430 ;
        RECT 106.985 107.630 107.215 112.780 ;
        RECT 106.750 106.930 107.450 107.630 ;
        RECT 106.985 104.780 107.215 106.930 ;
        RECT 108.325 104.780 108.555 112.780 ;
        RECT 110.615 104.780 110.845 112.780 ;
        RECT 112.905 104.780 113.135 112.780 ;
        RECT 79.005 104.275 80.965 104.575 ;
        RECT 81.295 104.275 83.255 104.575 ;
        RECT 84.925 104.275 86.885 104.575 ;
        RECT 87.215 104.275 89.175 104.575 ;
        RECT 90.845 104.275 95.095 104.575 ;
        RECT 96.765 104.275 98.725 104.575 ;
        RECT 99.055 104.275 101.015 104.575 ;
        RECT 102.685 104.275 104.645 104.575 ;
        RECT 104.975 104.275 106.935 104.575 ;
        RECT 108.325 103.885 113.135 104.780 ;
        RECT 113.575 103.885 114.165 123.695 ;
        RECT 128.935 123.505 135.120 124.285 ;
        RECT 138.080 128.380 145.960 128.970 ;
        RECT 138.080 124.680 138.670 128.380 ;
        RECT 139.205 127.290 139.435 127.530 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.205 125.530 139.435 125.690 ;
        RECT 140.495 125.530 140.725 128.380 ;
        RECT 143.725 127.920 144.425 127.990 ;
        RECT 143.595 127.690 144.555 127.920 ;
        RECT 141.785 127.290 142.015 127.530 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 143.315 126.865 143.545 127.530 ;
        RECT 143.280 126.165 143.580 126.865 ;
        RECT 141.785 125.530 142.015 125.690 ;
        RECT 143.315 125.370 143.545 126.165 ;
        RECT 139.390 125.140 143.545 125.370 ;
        RECT 144.605 124.680 144.835 127.530 ;
        RECT 145.370 124.680 145.960 128.380 ;
        RECT 138.080 124.090 145.960 124.680 ;
        RECT 71.775 102.705 114.165 103.885 ;
        RECT 115.905 122.915 135.120 123.505 ;
        RECT 115.905 122.475 116.495 122.915 ;
        RECT 115.905 122.245 118.390 122.475 ;
        RECT 115.905 114.185 117.185 122.245 ;
        RECT 118.595 114.235 118.825 122.195 ;
        RECT 119.975 118.645 120.205 122.195 ;
        RECT 120.410 122.010 121.410 122.710 ;
        RECT 121.615 118.645 121.845 122.195 ;
        RECT 119.975 117.075 121.845 118.645 ;
        RECT 115.905 113.955 118.390 114.185 ;
        RECT 115.905 112.845 116.495 113.955 ;
        RECT 115.905 112.615 118.390 112.845 ;
        RECT 115.905 104.555 117.185 112.615 ;
        RECT 118.595 104.605 118.825 112.565 ;
        RECT 119.975 109.685 120.205 117.075 ;
        RECT 121.615 114.235 121.845 117.075 ;
        RECT 122.995 118.645 123.225 122.195 ;
        RECT 123.430 122.010 124.430 122.710 ;
        RECT 128.345 122.475 135.120 122.915 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 126.450 122.245 135.120 122.475 ;
        RECT 124.635 118.645 124.865 122.195 ;
        RECT 122.995 117.075 124.865 118.645 ;
        RECT 122.995 114.235 123.225 117.075 ;
        RECT 120.410 112.615 121.410 114.185 ;
        RECT 123.430 112.615 124.430 114.185 ;
        RECT 121.615 109.685 121.845 112.565 ;
        RECT 119.975 108.115 121.845 109.685 ;
        RECT 119.975 104.605 120.205 108.115 ;
        RECT 115.905 104.325 118.390 104.555 ;
        RECT 115.905 103.885 116.495 104.325 ;
        RECT 120.410 104.090 121.410 104.790 ;
        RECT 121.615 104.605 121.845 108.115 ;
        RECT 122.995 109.685 123.225 112.565 ;
        RECT 124.635 109.685 124.865 117.075 ;
        RECT 126.015 114.235 126.245 122.195 ;
        RECT 127.655 114.185 135.120 122.245 ;
        RECT 126.450 113.955 135.120 114.185 ;
        RECT 128.345 112.845 135.120 113.955 ;
        RECT 126.450 112.615 135.120 112.845 ;
        RECT 122.995 108.115 124.865 109.685 ;
        RECT 122.995 104.605 123.225 108.115 ;
        RECT 123.430 104.090 124.430 104.790 ;
        RECT 124.635 104.605 124.865 108.115 ;
        RECT 126.015 104.605 126.245 112.565 ;
        RECT 127.655 107.765 135.120 112.615 ;
        RECT 136.295 108.925 142.995 109.515 ;
        RECT 127.655 104.835 138.400 107.765 ;
        RECT 127.655 104.555 135.710 104.835 ;
        RECT 126.450 104.325 135.710 104.555 ;
        RECT 128.345 103.885 135.710 104.325 ;
        RECT 115.905 102.705 135.710 103.885 ;
        RECT 8.665 102.115 135.710 102.705 ;
        RECT 136.295 102.495 138.400 104.255 ;
        RECT 8.665 44.835 10.615 102.115 ;
        RECT 4.100 42.225 10.615 44.835 ;
        RECT 11.055 101.425 29.605 102.115 ;
        RECT 11.055 93.015 11.285 101.425 ;
        RECT 13.345 93.015 13.575 101.425 ;
        RECT 15.635 93.015 15.865 101.425 ;
        RECT 17.925 93.015 18.155 101.425 ;
        RECT 20.215 93.015 20.445 101.425 ;
        RECT 22.505 93.015 22.735 101.425 ;
        RECT 24.795 93.015 25.025 101.425 ;
        RECT 27.085 93.015 27.315 101.425 ;
        RECT 29.375 93.015 29.605 101.425 ;
        RECT 30.715 101.425 49.265 102.115 ;
        RECT 30.715 93.220 30.945 101.425 ;
        RECT 33.005 93.220 33.235 101.425 ;
        RECT 35.295 93.220 35.525 101.425 ;
        RECT 37.585 93.220 37.815 101.425 ;
        RECT 39.875 93.220 40.105 101.425 ;
        RECT 42.165 93.220 42.395 101.425 ;
        RECT 44.455 93.220 44.685 101.425 ;
        RECT 46.745 93.220 46.975 101.425 ;
        RECT 49.035 93.220 49.265 101.425 ;
        RECT 50.375 101.425 68.925 102.115 ;
        RECT 50.375 93.220 50.605 101.425 ;
        RECT 52.665 93.220 52.895 101.425 ;
        RECT 54.955 93.220 55.185 101.425 ;
        RECT 57.245 93.220 57.475 101.425 ;
        RECT 59.535 93.220 59.765 101.425 ;
        RECT 61.825 93.220 62.055 101.425 ;
        RECT 64.115 93.220 64.345 101.425 ;
        RECT 66.405 93.220 66.635 101.425 ;
        RECT 68.695 93.220 68.925 101.425 ;
        RECT 70.035 101.425 88.585 102.115 ;
        RECT 70.035 93.220 70.265 101.425 ;
        RECT 72.325 93.220 72.555 101.425 ;
        RECT 74.615 93.220 74.845 101.425 ;
        RECT 76.905 93.220 77.135 101.425 ;
        RECT 79.195 93.220 79.425 101.425 ;
        RECT 81.485 93.220 81.715 101.425 ;
        RECT 83.775 93.220 84.005 101.425 ;
        RECT 86.065 93.220 86.295 101.425 ;
        RECT 88.355 93.220 88.585 101.425 ;
        RECT 89.695 101.425 108.245 102.115 ;
        RECT 89.695 93.220 89.925 101.425 ;
        RECT 91.985 93.220 92.215 101.425 ;
        RECT 94.275 93.220 94.505 101.425 ;
        RECT 96.565 93.220 96.795 101.425 ;
        RECT 98.855 93.220 99.085 101.425 ;
        RECT 101.145 93.220 101.375 101.425 ;
        RECT 103.435 93.220 103.665 101.425 ;
        RECT 105.725 93.220 105.955 101.425 ;
        RECT 108.015 93.220 108.245 101.425 ;
        RECT 109.355 101.425 127.905 102.115 ;
        RECT 109.355 93.015 109.585 101.425 ;
        RECT 111.645 93.015 111.875 101.425 ;
        RECT 113.935 93.015 114.165 101.425 ;
        RECT 116.225 93.015 116.455 101.425 ;
        RECT 118.515 93.015 118.745 101.425 ;
        RECT 120.805 93.015 121.035 101.425 ;
        RECT 123.095 93.015 123.325 101.425 ;
        RECT 125.385 93.015 125.615 101.425 ;
        RECT 127.675 93.015 127.905 101.425 ;
        RECT 11.055 91.405 29.605 93.015 ;
        RECT 30.995 92.785 32.955 93.015 ;
        RECT 33.285 92.785 35.245 93.015 ;
        RECT 35.575 92.785 37.535 93.015 ;
        RECT 37.865 92.785 39.825 93.015 ;
        RECT 40.155 92.785 42.115 93.015 ;
        RECT 42.445 92.785 44.405 93.015 ;
        RECT 44.735 92.785 46.695 93.015 ;
        RECT 47.025 92.785 48.985 93.015 ;
        RECT 50.655 92.785 52.615 93.015 ;
        RECT 52.945 92.785 54.905 93.015 ;
        RECT 55.235 92.785 57.195 93.015 ;
        RECT 57.525 92.785 59.485 93.015 ;
        RECT 59.815 92.785 61.775 93.015 ;
        RECT 62.105 92.785 64.065 93.015 ;
        RECT 64.395 92.785 66.355 93.015 ;
        RECT 66.685 92.785 68.645 93.015 ;
        RECT 70.315 92.785 72.275 93.015 ;
        RECT 72.605 92.785 74.565 93.015 ;
        RECT 74.895 92.785 76.855 93.015 ;
        RECT 77.185 92.785 79.145 93.015 ;
        RECT 79.475 92.785 81.435 93.015 ;
        RECT 81.765 92.785 83.725 93.015 ;
        RECT 84.055 92.785 86.015 93.015 ;
        RECT 86.345 92.785 88.305 93.015 ;
        RECT 89.975 92.785 91.935 93.015 ;
        RECT 92.265 92.785 94.225 93.015 ;
        RECT 94.555 92.785 96.515 93.015 ;
        RECT 96.845 92.785 98.805 93.015 ;
        RECT 99.135 92.785 101.095 93.015 ;
        RECT 101.425 92.785 103.385 93.015 ;
        RECT 103.715 92.785 105.675 93.015 ;
        RECT 106.005 92.785 107.965 93.015 ;
        RECT 30.995 91.405 32.955 91.635 ;
        RECT 11.055 82.995 11.285 91.405 ;
        RECT 13.345 82.995 13.575 91.405 ;
        RECT 15.635 82.995 15.865 91.405 ;
        RECT 17.925 82.995 18.155 91.405 ;
        RECT 20.215 82.995 20.445 91.405 ;
        RECT 22.505 82.995 22.735 91.405 ;
        RECT 24.795 82.995 25.025 91.405 ;
        RECT 27.085 82.995 27.315 91.405 ;
        RECT 29.375 82.995 29.605 91.405 ;
        RECT 33.285 91.345 35.245 91.875 ;
        RECT 35.575 91.345 37.535 91.875 ;
        RECT 37.865 91.405 39.825 91.635 ;
        RECT 40.155 91.405 42.115 91.635 ;
        RECT 42.445 91.345 44.405 91.875 ;
        RECT 44.735 91.345 46.695 91.875 ;
        RECT 47.025 91.405 48.985 91.635 ;
        RECT 50.655 91.345 52.615 91.875 ;
        RECT 52.945 91.405 54.905 91.635 ;
        RECT 55.235 91.405 57.195 91.635 ;
        RECT 57.525 91.345 59.485 91.875 ;
        RECT 59.815 91.345 61.775 91.875 ;
        RECT 62.105 91.405 64.065 91.635 ;
        RECT 64.395 91.405 66.355 91.635 ;
        RECT 66.685 91.345 68.645 91.875 ;
        RECT 70.315 91.345 72.275 91.875 ;
        RECT 72.605 91.405 74.565 91.635 ;
        RECT 74.895 91.405 76.855 91.635 ;
        RECT 77.185 91.345 79.145 91.875 ;
        RECT 79.475 91.345 81.435 91.875 ;
        RECT 81.765 91.405 83.725 91.635 ;
        RECT 84.055 91.405 86.015 91.635 ;
        RECT 86.345 91.345 88.305 91.875 ;
        RECT 89.975 91.405 91.935 91.635 ;
        RECT 92.265 91.345 94.225 91.875 ;
        RECT 94.555 91.345 96.515 91.875 ;
        RECT 96.845 91.405 98.805 91.635 ;
        RECT 99.135 91.405 101.095 91.635 ;
        RECT 101.425 91.345 103.385 91.875 ;
        RECT 103.715 91.345 105.675 91.875 ;
        RECT 106.005 91.405 107.965 91.635 ;
        RECT 109.355 91.405 127.905 93.015 ;
        RECT 30.715 84.590 30.945 91.200 ;
        RECT 33.005 88.540 33.235 91.200 ;
        RECT 35.295 91.090 35.525 91.200 ;
        RECT 35.260 89.690 35.560 91.090 ;
        RECT 32.970 85.740 33.270 88.540 ;
        RECT 30.680 83.190 30.980 84.590 ;
        RECT 33.005 83.200 33.235 85.740 ;
        RECT 35.295 83.200 35.525 89.690 ;
        RECT 37.585 88.540 37.815 91.200 ;
        RECT 37.550 85.740 37.850 88.540 ;
        RECT 37.585 83.200 37.815 85.740 ;
        RECT 39.875 84.590 40.105 91.200 ;
        RECT 42.165 88.540 42.395 91.200 ;
        RECT 44.455 91.090 44.685 91.200 ;
        RECT 44.420 89.690 44.720 91.090 ;
        RECT 42.130 85.740 42.430 88.540 ;
        RECT 39.840 83.190 40.140 84.590 ;
        RECT 42.165 83.200 42.395 85.740 ;
        RECT 44.455 83.200 44.685 89.690 ;
        RECT 46.745 88.540 46.975 91.200 ;
        RECT 46.710 85.740 47.010 88.540 ;
        RECT 46.745 83.200 46.975 85.740 ;
        RECT 49.035 84.590 49.265 91.200 ;
        RECT 50.375 91.090 50.605 91.200 ;
        RECT 50.340 89.690 50.640 91.090 ;
        RECT 49.000 83.190 49.300 84.590 ;
        RECT 50.375 83.200 50.605 89.690 ;
        RECT 52.665 88.540 52.895 91.200 ;
        RECT 52.630 85.740 52.930 88.540 ;
        RECT 52.665 83.200 52.895 85.740 ;
        RECT 54.955 84.590 55.185 91.200 ;
        RECT 57.245 88.540 57.475 91.200 ;
        RECT 59.535 91.090 59.765 91.200 ;
        RECT 59.500 89.690 59.800 91.090 ;
        RECT 57.210 85.740 57.510 88.540 ;
        RECT 54.920 83.190 55.220 84.590 ;
        RECT 57.245 83.200 57.475 85.740 ;
        RECT 59.535 83.200 59.765 89.690 ;
        RECT 61.825 88.540 62.055 91.200 ;
        RECT 61.790 85.740 62.090 88.540 ;
        RECT 61.825 83.200 62.055 85.740 ;
        RECT 64.115 84.590 64.345 91.200 ;
        RECT 66.405 88.540 66.635 91.200 ;
        RECT 68.695 91.090 68.925 91.200 ;
        RECT 70.035 91.090 70.265 91.200 ;
        RECT 68.660 89.690 68.960 91.090 ;
        RECT 70.000 89.690 70.300 91.090 ;
        RECT 66.370 85.740 66.670 88.540 ;
        RECT 64.080 83.190 64.380 84.590 ;
        RECT 66.405 83.200 66.635 85.740 ;
        RECT 68.695 83.200 68.925 89.690 ;
        RECT 70.035 83.200 70.265 89.690 ;
        RECT 72.325 88.540 72.555 91.200 ;
        RECT 72.290 85.740 72.590 88.540 ;
        RECT 72.325 83.200 72.555 85.740 ;
        RECT 74.615 84.590 74.845 91.200 ;
        RECT 76.905 88.540 77.135 91.200 ;
        RECT 79.195 91.090 79.425 91.200 ;
        RECT 79.160 89.690 79.460 91.090 ;
        RECT 76.870 85.740 77.170 88.540 ;
        RECT 74.580 83.190 74.880 84.590 ;
        RECT 76.905 83.200 77.135 85.740 ;
        RECT 79.195 83.200 79.425 89.690 ;
        RECT 81.485 88.540 81.715 91.200 ;
        RECT 81.450 85.740 81.750 88.540 ;
        RECT 81.485 83.200 81.715 85.740 ;
        RECT 83.775 84.590 84.005 91.200 ;
        RECT 86.065 88.540 86.295 91.200 ;
        RECT 88.355 91.090 88.585 91.200 ;
        RECT 88.320 89.690 88.620 91.090 ;
        RECT 86.030 85.740 86.330 88.540 ;
        RECT 83.740 83.190 84.040 84.590 ;
        RECT 86.065 83.200 86.295 85.740 ;
        RECT 88.355 83.200 88.585 89.690 ;
        RECT 89.695 84.590 89.925 91.200 ;
        RECT 91.985 88.540 92.215 91.200 ;
        RECT 94.275 91.090 94.505 91.200 ;
        RECT 94.240 89.690 94.540 91.090 ;
        RECT 91.950 85.740 92.250 88.540 ;
        RECT 89.660 83.190 89.960 84.590 ;
        RECT 91.985 83.200 92.215 85.740 ;
        RECT 94.275 83.200 94.505 89.690 ;
        RECT 96.565 88.540 96.795 91.200 ;
        RECT 96.530 85.740 96.830 88.540 ;
        RECT 96.565 83.200 96.795 85.740 ;
        RECT 98.855 84.590 99.085 91.200 ;
        RECT 101.145 88.540 101.375 91.200 ;
        RECT 103.435 91.090 103.665 91.200 ;
        RECT 103.400 89.690 103.700 91.090 ;
        RECT 101.110 85.740 101.410 88.540 ;
        RECT 98.820 83.190 99.120 84.590 ;
        RECT 101.145 83.200 101.375 85.740 ;
        RECT 103.435 83.200 103.665 89.690 ;
        RECT 105.725 88.540 105.955 91.200 ;
        RECT 105.690 85.740 105.990 88.540 ;
        RECT 105.725 83.200 105.955 85.740 ;
        RECT 108.015 84.590 108.245 91.200 ;
        RECT 107.980 83.190 108.280 84.590 ;
        RECT 109.355 82.995 109.585 91.405 ;
        RECT 111.645 82.995 111.875 91.405 ;
        RECT 113.935 82.995 114.165 91.405 ;
        RECT 116.225 82.995 116.455 91.405 ;
        RECT 118.515 82.995 118.745 91.405 ;
        RECT 120.805 82.995 121.035 91.405 ;
        RECT 123.095 82.995 123.325 91.405 ;
        RECT 125.385 82.995 125.615 91.405 ;
        RECT 127.675 82.995 127.905 91.405 ;
        RECT 11.055 81.385 29.605 82.995 ;
        RECT 30.995 82.405 32.955 82.995 ;
        RECT 33.285 82.765 35.245 82.995 ;
        RECT 35.575 82.765 37.535 82.995 ;
        RECT 37.865 82.405 39.825 82.995 ;
        RECT 40.155 82.405 42.115 82.995 ;
        RECT 42.445 82.765 44.405 82.995 ;
        RECT 44.735 82.765 46.695 82.995 ;
        RECT 47.025 82.405 48.985 82.995 ;
        RECT 50.655 82.765 52.615 82.995 ;
        RECT 52.945 82.405 54.905 82.995 ;
        RECT 55.235 82.405 57.195 82.995 ;
        RECT 57.525 82.765 59.485 82.995 ;
        RECT 59.815 82.765 61.775 82.995 ;
        RECT 62.105 82.405 64.065 82.995 ;
        RECT 64.395 82.405 66.355 82.995 ;
        RECT 66.685 82.765 68.645 82.995 ;
        RECT 70.315 82.765 72.275 82.995 ;
        RECT 72.605 82.405 74.565 82.995 ;
        RECT 74.895 82.405 76.855 82.995 ;
        RECT 77.185 82.765 79.145 82.995 ;
        RECT 79.475 82.765 81.435 82.995 ;
        RECT 81.765 82.405 83.725 82.995 ;
        RECT 84.055 82.405 86.015 82.995 ;
        RECT 86.345 82.765 88.305 82.995 ;
        RECT 89.975 82.405 91.935 82.995 ;
        RECT 92.265 82.765 94.225 82.995 ;
        RECT 94.555 82.765 96.515 82.995 ;
        RECT 96.845 82.405 98.805 82.995 ;
        RECT 99.135 82.405 101.095 82.995 ;
        RECT 101.425 82.765 103.385 82.995 ;
        RECT 103.715 82.765 105.675 82.995 ;
        RECT 106.005 82.405 107.965 82.995 ;
        RECT 30.995 81.385 32.955 81.615 ;
        RECT 11.055 72.975 11.285 81.385 ;
        RECT 13.345 72.975 13.575 81.385 ;
        RECT 15.635 72.975 15.865 81.385 ;
        RECT 17.925 72.975 18.155 81.385 ;
        RECT 20.215 72.975 20.445 81.385 ;
        RECT 22.505 72.975 22.735 81.385 ;
        RECT 24.795 72.975 25.025 81.385 ;
        RECT 27.085 72.975 27.315 81.385 ;
        RECT 29.375 72.975 29.605 81.385 ;
        RECT 33.285 81.325 35.245 81.855 ;
        RECT 35.575 81.325 37.535 81.855 ;
        RECT 37.865 81.385 39.825 81.615 ;
        RECT 40.155 81.385 42.115 81.615 ;
        RECT 42.445 81.325 44.405 81.855 ;
        RECT 44.735 81.325 46.695 81.855 ;
        RECT 47.025 81.385 48.985 81.615 ;
        RECT 50.655 81.325 52.615 81.855 ;
        RECT 52.945 81.385 54.905 81.615 ;
        RECT 55.235 81.385 57.195 81.615 ;
        RECT 57.525 81.325 59.485 81.855 ;
        RECT 59.815 81.325 61.775 81.855 ;
        RECT 62.105 81.385 64.065 81.615 ;
        RECT 64.395 81.385 66.355 81.615 ;
        RECT 66.685 81.325 68.645 81.855 ;
        RECT 70.315 81.325 72.275 81.855 ;
        RECT 72.605 81.385 74.565 81.615 ;
        RECT 74.895 81.385 76.855 81.615 ;
        RECT 77.185 81.325 79.145 81.855 ;
        RECT 79.475 81.325 81.435 81.855 ;
        RECT 81.765 81.385 83.725 81.615 ;
        RECT 84.055 81.385 86.015 81.615 ;
        RECT 86.345 81.325 88.305 81.855 ;
        RECT 89.975 81.385 91.935 81.615 ;
        RECT 92.265 81.325 94.225 81.855 ;
        RECT 94.555 81.325 96.515 81.855 ;
        RECT 96.845 81.385 98.805 81.615 ;
        RECT 99.135 81.385 101.095 81.615 ;
        RECT 101.425 81.325 103.385 81.855 ;
        RECT 103.715 81.325 105.675 81.855 ;
        RECT 106.005 81.385 107.965 81.615 ;
        RECT 109.355 81.385 127.905 82.995 ;
        RECT 30.715 81.070 30.945 81.180 ;
        RECT 30.680 79.670 30.980 81.070 ;
        RECT 30.715 73.180 30.945 79.670 ;
        RECT 33.005 78.520 33.235 81.180 ;
        RECT 32.970 75.720 33.270 78.520 ;
        RECT 33.005 73.180 33.235 75.720 ;
        RECT 35.295 74.570 35.525 81.180 ;
        RECT 37.585 78.520 37.815 81.180 ;
        RECT 39.875 81.070 40.105 81.180 ;
        RECT 39.840 79.670 40.140 81.070 ;
        RECT 37.550 75.720 37.850 78.520 ;
        RECT 35.260 73.170 35.560 74.570 ;
        RECT 37.585 73.180 37.815 75.720 ;
        RECT 39.875 73.180 40.105 79.670 ;
        RECT 42.165 78.520 42.395 81.180 ;
        RECT 42.130 75.720 42.430 78.520 ;
        RECT 42.165 73.180 42.395 75.720 ;
        RECT 44.455 74.570 44.685 81.180 ;
        RECT 46.745 78.520 46.975 81.180 ;
        RECT 49.035 81.070 49.265 81.180 ;
        RECT 49.000 79.670 49.300 81.070 ;
        RECT 46.710 75.720 47.010 78.520 ;
        RECT 44.420 73.170 44.720 74.570 ;
        RECT 46.745 73.180 46.975 75.720 ;
        RECT 49.035 73.180 49.265 79.670 ;
        RECT 50.375 74.570 50.605 81.180 ;
        RECT 52.665 78.520 52.895 81.180 ;
        RECT 54.955 81.070 55.185 81.180 ;
        RECT 54.920 79.670 55.220 81.070 ;
        RECT 52.630 75.720 52.930 78.520 ;
        RECT 50.340 73.170 50.640 74.570 ;
        RECT 52.665 73.180 52.895 75.720 ;
        RECT 54.955 73.180 55.185 79.670 ;
        RECT 57.245 78.520 57.475 81.180 ;
        RECT 57.210 75.720 57.510 78.520 ;
        RECT 57.245 73.180 57.475 75.720 ;
        RECT 59.535 74.570 59.765 81.180 ;
        RECT 61.825 78.520 62.055 81.180 ;
        RECT 64.115 81.070 64.345 81.180 ;
        RECT 64.080 79.670 64.380 81.070 ;
        RECT 61.790 75.720 62.090 78.520 ;
        RECT 59.500 73.170 59.800 74.570 ;
        RECT 61.825 73.180 62.055 75.720 ;
        RECT 64.115 73.180 64.345 79.670 ;
        RECT 66.405 78.520 66.635 81.180 ;
        RECT 66.370 75.720 66.670 78.520 ;
        RECT 66.405 73.180 66.635 75.720 ;
        RECT 68.695 74.570 68.925 81.180 ;
        RECT 70.035 74.570 70.265 81.180 ;
        RECT 72.325 78.520 72.555 81.180 ;
        RECT 74.615 81.070 74.845 81.180 ;
        RECT 74.580 79.670 74.880 81.070 ;
        RECT 72.290 75.720 72.590 78.520 ;
        RECT 68.660 73.170 68.960 74.570 ;
        RECT 70.000 73.170 70.300 74.570 ;
        RECT 72.325 73.180 72.555 75.720 ;
        RECT 74.615 73.180 74.845 79.670 ;
        RECT 76.905 78.520 77.135 81.180 ;
        RECT 76.870 75.720 77.170 78.520 ;
        RECT 76.905 73.180 77.135 75.720 ;
        RECT 79.195 74.570 79.425 81.180 ;
        RECT 81.485 78.520 81.715 81.180 ;
        RECT 83.775 81.070 84.005 81.180 ;
        RECT 83.740 79.670 84.040 81.070 ;
        RECT 81.450 75.720 81.750 78.520 ;
        RECT 79.160 73.170 79.460 74.570 ;
        RECT 81.485 73.180 81.715 75.720 ;
        RECT 83.775 73.180 84.005 79.670 ;
        RECT 86.065 78.520 86.295 81.180 ;
        RECT 86.030 75.720 86.330 78.520 ;
        RECT 86.065 73.180 86.295 75.720 ;
        RECT 88.355 74.570 88.585 81.180 ;
        RECT 89.695 81.070 89.925 81.180 ;
        RECT 89.660 79.670 89.960 81.070 ;
        RECT 88.320 73.170 88.620 74.570 ;
        RECT 89.695 73.180 89.925 79.670 ;
        RECT 91.985 78.520 92.215 81.180 ;
        RECT 91.950 75.720 92.250 78.520 ;
        RECT 91.985 73.180 92.215 75.720 ;
        RECT 94.275 74.570 94.505 81.180 ;
        RECT 96.565 78.520 96.795 81.180 ;
        RECT 98.855 81.070 99.085 81.180 ;
        RECT 98.820 79.670 99.120 81.070 ;
        RECT 96.530 75.720 96.830 78.520 ;
        RECT 94.240 73.170 94.540 74.570 ;
        RECT 96.565 73.180 96.795 75.720 ;
        RECT 98.855 73.180 99.085 79.670 ;
        RECT 101.145 78.520 101.375 81.180 ;
        RECT 101.110 75.720 101.410 78.520 ;
        RECT 101.145 73.180 101.375 75.720 ;
        RECT 103.435 74.570 103.665 81.180 ;
        RECT 105.725 78.520 105.955 81.180 ;
        RECT 108.015 81.070 108.245 81.180 ;
        RECT 107.980 79.670 108.280 81.070 ;
        RECT 105.690 75.720 105.990 78.520 ;
        RECT 103.400 73.170 103.700 74.570 ;
        RECT 105.725 73.180 105.955 75.720 ;
        RECT 108.015 73.180 108.245 79.670 ;
        RECT 109.355 72.975 109.585 81.385 ;
        RECT 111.645 72.975 111.875 81.385 ;
        RECT 113.935 72.975 114.165 81.385 ;
        RECT 116.225 72.975 116.455 81.385 ;
        RECT 118.515 72.975 118.745 81.385 ;
        RECT 120.805 72.975 121.035 81.385 ;
        RECT 123.095 72.975 123.325 81.385 ;
        RECT 125.385 72.975 125.615 81.385 ;
        RECT 127.675 72.975 127.905 81.385 ;
        RECT 11.055 71.365 29.605 72.975 ;
        RECT 30.995 72.385 32.955 72.975 ;
        RECT 33.285 72.745 35.245 72.975 ;
        RECT 35.575 72.745 37.535 72.975 ;
        RECT 37.865 72.385 39.825 72.975 ;
        RECT 40.155 72.385 42.115 72.975 ;
        RECT 42.445 72.745 44.405 72.975 ;
        RECT 44.735 72.745 46.695 72.975 ;
        RECT 47.025 72.385 48.985 72.975 ;
        RECT 50.655 72.745 52.615 72.975 ;
        RECT 52.945 72.385 54.905 72.975 ;
        RECT 55.235 72.385 57.195 72.975 ;
        RECT 57.525 72.745 59.485 72.975 ;
        RECT 59.815 72.745 61.775 72.975 ;
        RECT 62.105 72.385 64.065 72.975 ;
        RECT 64.395 72.385 66.355 72.975 ;
        RECT 66.685 72.745 68.645 72.975 ;
        RECT 70.315 72.745 72.275 72.975 ;
        RECT 72.605 72.385 74.565 72.975 ;
        RECT 74.895 72.385 76.855 72.975 ;
        RECT 77.185 72.745 79.145 72.975 ;
        RECT 79.475 72.745 81.435 72.975 ;
        RECT 81.765 72.385 83.725 72.975 ;
        RECT 84.055 72.385 86.015 72.975 ;
        RECT 86.345 72.745 88.305 72.975 ;
        RECT 89.975 72.385 91.935 72.975 ;
        RECT 92.265 72.745 94.225 72.975 ;
        RECT 94.555 72.745 96.515 72.975 ;
        RECT 96.845 72.385 98.805 72.975 ;
        RECT 99.135 72.385 101.095 72.975 ;
        RECT 101.425 72.745 103.385 72.975 ;
        RECT 103.715 72.745 105.675 72.975 ;
        RECT 106.005 72.385 107.965 72.975 ;
        RECT 11.055 62.955 11.285 71.365 ;
        RECT 13.345 62.955 13.575 71.365 ;
        RECT 15.635 62.955 15.865 71.365 ;
        RECT 17.925 62.955 18.155 71.365 ;
        RECT 20.215 62.955 20.445 71.365 ;
        RECT 22.505 62.955 22.735 71.365 ;
        RECT 24.795 62.955 25.025 71.365 ;
        RECT 27.085 62.955 27.315 71.365 ;
        RECT 29.375 62.955 29.605 71.365 ;
        RECT 30.995 71.305 32.955 71.835 ;
        RECT 33.285 71.365 35.245 71.595 ;
        RECT 35.575 71.365 37.535 71.595 ;
        RECT 37.865 71.305 39.825 71.835 ;
        RECT 40.155 71.305 42.115 71.835 ;
        RECT 42.445 71.365 44.405 71.595 ;
        RECT 44.735 71.365 46.695 71.595 ;
        RECT 47.025 71.305 48.985 71.835 ;
        RECT 50.655 71.365 52.615 71.595 ;
        RECT 52.945 71.305 54.905 71.835 ;
        RECT 55.235 71.305 57.195 71.835 ;
        RECT 57.525 71.365 59.485 71.595 ;
        RECT 59.815 71.365 61.775 71.595 ;
        RECT 62.105 71.305 64.065 71.835 ;
        RECT 64.395 71.305 66.355 71.835 ;
        RECT 66.685 71.365 68.645 71.595 ;
        RECT 70.315 71.365 72.275 71.595 ;
        RECT 72.605 71.305 74.565 71.835 ;
        RECT 74.895 71.305 76.855 71.835 ;
        RECT 77.185 71.365 79.145 71.595 ;
        RECT 79.475 71.365 81.435 71.595 ;
        RECT 81.765 71.305 83.725 71.835 ;
        RECT 84.055 71.305 86.015 71.835 ;
        RECT 86.345 71.365 88.305 71.595 ;
        RECT 89.975 71.305 91.935 71.835 ;
        RECT 92.265 71.365 94.225 71.595 ;
        RECT 94.555 71.365 96.515 71.595 ;
        RECT 96.845 71.305 98.805 71.835 ;
        RECT 99.135 71.305 101.095 71.835 ;
        RECT 101.425 71.365 103.385 71.595 ;
        RECT 103.715 71.365 105.675 71.595 ;
        RECT 106.005 71.305 107.965 71.835 ;
        RECT 109.355 71.365 127.905 72.975 ;
        RECT 30.715 71.050 30.945 71.160 ;
        RECT 30.680 69.650 30.980 71.050 ;
        RECT 30.715 63.160 30.945 69.650 ;
        RECT 33.005 68.500 33.235 71.160 ;
        RECT 32.970 65.700 33.270 68.500 ;
        RECT 33.005 63.160 33.235 65.700 ;
        RECT 35.295 64.550 35.525 71.160 ;
        RECT 37.585 68.500 37.815 71.160 ;
        RECT 39.875 71.050 40.105 71.160 ;
        RECT 39.840 69.650 40.140 71.050 ;
        RECT 37.550 65.700 37.850 68.500 ;
        RECT 35.260 63.150 35.560 64.550 ;
        RECT 37.585 63.160 37.815 65.700 ;
        RECT 39.875 63.160 40.105 69.650 ;
        RECT 42.165 68.500 42.395 71.160 ;
        RECT 42.130 65.700 42.430 68.500 ;
        RECT 42.165 63.160 42.395 65.700 ;
        RECT 44.455 64.550 44.685 71.160 ;
        RECT 46.745 68.500 46.975 71.160 ;
        RECT 49.035 71.050 49.265 71.160 ;
        RECT 49.000 69.650 49.300 71.050 ;
        RECT 46.710 65.700 47.010 68.500 ;
        RECT 44.420 63.150 44.720 64.550 ;
        RECT 46.745 63.160 46.975 65.700 ;
        RECT 49.035 63.160 49.265 69.650 ;
        RECT 50.375 64.550 50.605 71.160 ;
        RECT 52.665 68.500 52.895 71.160 ;
        RECT 54.955 71.050 55.185 71.160 ;
        RECT 54.920 69.650 55.220 71.050 ;
        RECT 52.630 65.700 52.930 68.500 ;
        RECT 50.340 63.150 50.640 64.550 ;
        RECT 52.665 63.160 52.895 65.700 ;
        RECT 54.955 63.160 55.185 69.650 ;
        RECT 57.245 68.500 57.475 71.160 ;
        RECT 57.210 65.700 57.510 68.500 ;
        RECT 57.245 63.160 57.475 65.700 ;
        RECT 59.535 64.550 59.765 71.160 ;
        RECT 61.825 68.500 62.055 71.160 ;
        RECT 64.115 71.050 64.345 71.160 ;
        RECT 64.080 69.650 64.380 71.050 ;
        RECT 61.790 65.700 62.090 68.500 ;
        RECT 59.500 63.150 59.800 64.550 ;
        RECT 61.825 63.160 62.055 65.700 ;
        RECT 64.115 63.160 64.345 69.650 ;
        RECT 66.405 68.500 66.635 71.160 ;
        RECT 66.370 65.700 66.670 68.500 ;
        RECT 66.405 63.160 66.635 65.700 ;
        RECT 68.695 64.550 68.925 71.160 ;
        RECT 70.035 64.550 70.265 71.160 ;
        RECT 72.325 68.500 72.555 71.160 ;
        RECT 74.615 71.050 74.845 71.160 ;
        RECT 74.580 69.650 74.880 71.050 ;
        RECT 72.290 65.700 72.590 68.500 ;
        RECT 68.660 63.150 68.960 64.550 ;
        RECT 70.000 63.150 70.300 64.550 ;
        RECT 72.325 63.160 72.555 65.700 ;
        RECT 74.615 63.160 74.845 69.650 ;
        RECT 76.905 68.500 77.135 71.160 ;
        RECT 76.870 65.700 77.170 68.500 ;
        RECT 76.905 63.160 77.135 65.700 ;
        RECT 79.195 64.550 79.425 71.160 ;
        RECT 81.485 68.500 81.715 71.160 ;
        RECT 83.775 71.050 84.005 71.160 ;
        RECT 83.740 69.650 84.040 71.050 ;
        RECT 81.450 65.700 81.750 68.500 ;
        RECT 79.160 63.150 79.460 64.550 ;
        RECT 81.485 63.160 81.715 65.700 ;
        RECT 83.775 63.160 84.005 69.650 ;
        RECT 86.065 68.500 86.295 71.160 ;
        RECT 86.030 65.700 86.330 68.500 ;
        RECT 86.065 63.160 86.295 65.700 ;
        RECT 88.355 64.550 88.585 71.160 ;
        RECT 89.695 71.050 89.925 71.160 ;
        RECT 89.660 69.650 89.960 71.050 ;
        RECT 88.320 63.150 88.620 64.550 ;
        RECT 89.695 63.160 89.925 69.650 ;
        RECT 91.985 68.500 92.215 71.160 ;
        RECT 91.950 65.700 92.250 68.500 ;
        RECT 91.985 63.160 92.215 65.700 ;
        RECT 94.275 64.550 94.505 71.160 ;
        RECT 96.565 68.500 96.795 71.160 ;
        RECT 98.855 71.050 99.085 71.160 ;
        RECT 98.820 69.650 99.120 71.050 ;
        RECT 96.530 65.700 96.830 68.500 ;
        RECT 94.240 63.150 94.540 64.550 ;
        RECT 96.565 63.160 96.795 65.700 ;
        RECT 98.855 63.160 99.085 69.650 ;
        RECT 101.145 68.500 101.375 71.160 ;
        RECT 101.110 65.700 101.410 68.500 ;
        RECT 101.145 63.160 101.375 65.700 ;
        RECT 103.435 64.550 103.665 71.160 ;
        RECT 105.725 68.500 105.955 71.160 ;
        RECT 108.015 71.050 108.245 71.160 ;
        RECT 107.980 69.650 108.280 71.050 ;
        RECT 105.690 65.700 105.990 68.500 ;
        RECT 103.400 63.150 103.700 64.550 ;
        RECT 105.725 63.160 105.955 65.700 ;
        RECT 108.015 63.160 108.245 69.650 ;
        RECT 109.355 62.955 109.585 71.365 ;
        RECT 111.645 62.955 111.875 71.365 ;
        RECT 113.935 62.955 114.165 71.365 ;
        RECT 116.225 62.955 116.455 71.365 ;
        RECT 118.515 62.955 118.745 71.365 ;
        RECT 120.805 62.955 121.035 71.365 ;
        RECT 123.095 62.955 123.325 71.365 ;
        RECT 125.385 62.955 125.615 71.365 ;
        RECT 127.675 62.955 127.905 71.365 ;
        RECT 11.055 61.345 29.605 62.955 ;
        RECT 30.995 62.725 32.955 62.955 ;
        RECT 33.285 62.365 35.245 62.955 ;
        RECT 35.575 62.365 37.535 62.955 ;
        RECT 37.865 62.725 39.825 62.955 ;
        RECT 40.155 62.725 42.115 62.955 ;
        RECT 42.445 62.365 44.405 62.955 ;
        RECT 44.735 62.365 46.695 62.955 ;
        RECT 47.025 62.725 48.985 62.955 ;
        RECT 50.655 62.365 52.615 62.955 ;
        RECT 52.945 62.725 54.905 62.955 ;
        RECT 55.235 62.725 57.195 62.955 ;
        RECT 57.525 62.365 59.485 62.955 ;
        RECT 59.815 62.365 61.775 62.955 ;
        RECT 62.105 62.725 64.065 62.955 ;
        RECT 64.395 62.725 66.355 62.955 ;
        RECT 66.685 62.365 68.645 62.955 ;
        RECT 70.315 62.365 72.275 62.955 ;
        RECT 72.605 62.725 74.565 62.955 ;
        RECT 74.895 62.725 76.855 62.955 ;
        RECT 77.185 62.365 79.145 62.955 ;
        RECT 79.475 62.365 81.435 62.955 ;
        RECT 81.765 62.725 83.725 62.955 ;
        RECT 84.055 62.725 86.015 62.955 ;
        RECT 86.345 62.365 88.305 62.955 ;
        RECT 89.975 62.725 91.935 62.955 ;
        RECT 92.265 62.365 94.225 62.955 ;
        RECT 94.555 62.365 96.515 62.955 ;
        RECT 96.845 62.725 98.805 62.955 ;
        RECT 99.135 62.725 101.095 62.955 ;
        RECT 101.425 62.365 103.385 62.955 ;
        RECT 103.715 62.365 105.675 62.955 ;
        RECT 106.005 62.725 107.965 62.955 ;
        RECT 11.055 52.935 11.285 61.345 ;
        RECT 13.345 52.935 13.575 61.345 ;
        RECT 15.635 52.935 15.865 61.345 ;
        RECT 17.925 52.935 18.155 61.345 ;
        RECT 20.215 52.935 20.445 61.345 ;
        RECT 22.505 52.935 22.735 61.345 ;
        RECT 24.795 52.935 25.025 61.345 ;
        RECT 27.085 52.935 27.315 61.345 ;
        RECT 29.375 52.935 29.605 61.345 ;
        RECT 30.995 61.285 32.955 61.815 ;
        RECT 33.285 61.345 35.245 61.575 ;
        RECT 35.575 61.345 37.535 61.575 ;
        RECT 37.865 61.285 39.825 61.815 ;
        RECT 40.155 61.285 42.115 61.815 ;
        RECT 42.445 61.345 44.405 61.575 ;
        RECT 44.735 61.345 46.695 61.575 ;
        RECT 47.025 61.285 48.985 61.815 ;
        RECT 50.655 61.345 52.615 61.575 ;
        RECT 52.945 61.285 54.905 61.815 ;
        RECT 55.235 61.285 57.195 61.815 ;
        RECT 57.525 61.345 59.485 61.575 ;
        RECT 59.815 61.345 61.775 61.575 ;
        RECT 62.105 61.285 64.065 61.815 ;
        RECT 64.395 61.285 66.355 61.815 ;
        RECT 66.685 61.345 68.645 61.575 ;
        RECT 70.315 61.345 72.275 61.575 ;
        RECT 72.605 61.285 74.565 61.815 ;
        RECT 74.895 61.285 76.855 61.815 ;
        RECT 77.185 61.345 79.145 61.575 ;
        RECT 79.475 61.345 81.435 61.575 ;
        RECT 81.765 61.285 83.725 61.815 ;
        RECT 84.055 61.285 86.015 61.815 ;
        RECT 86.345 61.345 88.305 61.575 ;
        RECT 89.975 61.285 91.935 61.815 ;
        RECT 92.265 61.345 94.225 61.575 ;
        RECT 94.555 61.345 96.515 61.575 ;
        RECT 96.845 61.285 98.805 61.815 ;
        RECT 99.135 61.285 101.095 61.815 ;
        RECT 101.425 61.345 103.385 61.575 ;
        RECT 103.715 61.345 105.675 61.575 ;
        RECT 106.005 61.285 107.965 61.815 ;
        RECT 109.355 61.345 127.905 62.955 ;
        RECT 30.715 54.530 30.945 61.140 ;
        RECT 33.005 58.480 33.235 61.140 ;
        RECT 35.295 61.030 35.525 61.140 ;
        RECT 35.260 59.630 35.560 61.030 ;
        RECT 32.970 55.680 33.270 58.480 ;
        RECT 30.680 53.130 30.980 54.530 ;
        RECT 33.005 53.140 33.235 55.680 ;
        RECT 35.295 53.140 35.525 59.630 ;
        RECT 37.585 58.480 37.815 61.140 ;
        RECT 37.550 55.680 37.850 58.480 ;
        RECT 37.585 53.140 37.815 55.680 ;
        RECT 39.875 54.530 40.105 61.140 ;
        RECT 42.165 58.480 42.395 61.140 ;
        RECT 44.455 61.030 44.685 61.140 ;
        RECT 44.420 59.630 44.720 61.030 ;
        RECT 42.130 55.680 42.430 58.480 ;
        RECT 39.840 53.130 40.140 54.530 ;
        RECT 42.165 53.140 42.395 55.680 ;
        RECT 44.455 53.140 44.685 59.630 ;
        RECT 46.745 58.480 46.975 61.140 ;
        RECT 46.710 55.680 47.010 58.480 ;
        RECT 46.745 53.140 46.975 55.680 ;
        RECT 49.035 54.530 49.265 61.140 ;
        RECT 50.375 61.030 50.605 61.140 ;
        RECT 50.340 59.630 50.640 61.030 ;
        RECT 49.000 53.130 49.300 54.530 ;
        RECT 50.375 53.140 50.605 59.630 ;
        RECT 52.665 58.480 52.895 61.140 ;
        RECT 52.630 55.680 52.930 58.480 ;
        RECT 52.665 53.140 52.895 55.680 ;
        RECT 54.955 54.530 55.185 61.140 ;
        RECT 57.245 58.480 57.475 61.140 ;
        RECT 59.535 61.030 59.765 61.140 ;
        RECT 59.500 59.630 59.800 61.030 ;
        RECT 57.210 55.680 57.510 58.480 ;
        RECT 54.920 53.130 55.220 54.530 ;
        RECT 57.245 53.140 57.475 55.680 ;
        RECT 59.535 53.140 59.765 59.630 ;
        RECT 61.825 58.480 62.055 61.140 ;
        RECT 61.790 55.680 62.090 58.480 ;
        RECT 61.825 53.140 62.055 55.680 ;
        RECT 64.115 54.530 64.345 61.140 ;
        RECT 66.405 58.480 66.635 61.140 ;
        RECT 68.695 61.030 68.925 61.140 ;
        RECT 70.035 61.030 70.265 61.140 ;
        RECT 68.660 59.630 68.960 61.030 ;
        RECT 70.000 59.630 70.300 61.030 ;
        RECT 66.370 55.680 66.670 58.480 ;
        RECT 64.080 53.130 64.380 54.530 ;
        RECT 66.405 53.140 66.635 55.680 ;
        RECT 68.695 53.140 68.925 59.630 ;
        RECT 70.035 53.140 70.265 59.630 ;
        RECT 72.325 58.480 72.555 61.140 ;
        RECT 72.290 55.680 72.590 58.480 ;
        RECT 72.325 53.140 72.555 55.680 ;
        RECT 74.615 54.530 74.845 61.140 ;
        RECT 76.905 58.480 77.135 61.140 ;
        RECT 79.195 61.030 79.425 61.140 ;
        RECT 79.160 59.630 79.460 61.030 ;
        RECT 76.870 55.680 77.170 58.480 ;
        RECT 74.580 53.130 74.880 54.530 ;
        RECT 76.905 53.140 77.135 55.680 ;
        RECT 79.195 53.140 79.425 59.630 ;
        RECT 81.485 58.480 81.715 61.140 ;
        RECT 81.450 55.680 81.750 58.480 ;
        RECT 81.485 53.140 81.715 55.680 ;
        RECT 83.775 54.530 84.005 61.140 ;
        RECT 86.065 58.480 86.295 61.140 ;
        RECT 88.355 61.030 88.585 61.140 ;
        RECT 88.320 59.630 88.620 61.030 ;
        RECT 86.030 55.680 86.330 58.480 ;
        RECT 83.740 53.130 84.040 54.530 ;
        RECT 86.065 53.140 86.295 55.680 ;
        RECT 88.355 53.140 88.585 59.630 ;
        RECT 89.695 54.530 89.925 61.140 ;
        RECT 91.985 58.480 92.215 61.140 ;
        RECT 94.275 61.030 94.505 61.140 ;
        RECT 94.240 59.630 94.540 61.030 ;
        RECT 91.950 55.680 92.250 58.480 ;
        RECT 89.660 53.130 89.960 54.530 ;
        RECT 91.985 53.140 92.215 55.680 ;
        RECT 94.275 53.140 94.505 59.630 ;
        RECT 96.565 58.480 96.795 61.140 ;
        RECT 96.530 55.680 96.830 58.480 ;
        RECT 96.565 53.140 96.795 55.680 ;
        RECT 98.855 54.530 99.085 61.140 ;
        RECT 101.145 58.480 101.375 61.140 ;
        RECT 103.435 61.030 103.665 61.140 ;
        RECT 103.400 59.630 103.700 61.030 ;
        RECT 101.110 55.680 101.410 58.480 ;
        RECT 98.820 53.130 99.120 54.530 ;
        RECT 101.145 53.140 101.375 55.680 ;
        RECT 103.435 53.140 103.665 59.630 ;
        RECT 105.725 58.480 105.955 61.140 ;
        RECT 105.690 55.680 105.990 58.480 ;
        RECT 105.725 53.140 105.955 55.680 ;
        RECT 108.015 54.530 108.245 61.140 ;
        RECT 107.980 53.130 108.280 54.530 ;
        RECT 109.355 52.935 109.585 61.345 ;
        RECT 111.645 52.935 111.875 61.345 ;
        RECT 113.935 52.935 114.165 61.345 ;
        RECT 116.225 52.935 116.455 61.345 ;
        RECT 118.515 52.935 118.745 61.345 ;
        RECT 120.805 52.935 121.035 61.345 ;
        RECT 123.095 52.935 123.325 61.345 ;
        RECT 125.385 52.935 125.615 61.345 ;
        RECT 127.675 52.935 127.905 61.345 ;
        RECT 11.055 51.325 29.605 52.935 ;
        RECT 30.995 52.705 32.955 52.935 ;
        RECT 33.285 52.345 35.245 52.935 ;
        RECT 35.575 52.345 37.535 52.935 ;
        RECT 37.865 52.705 39.825 52.935 ;
        RECT 40.155 52.705 42.115 52.935 ;
        RECT 42.445 52.345 44.405 52.935 ;
        RECT 44.735 52.345 46.695 52.935 ;
        RECT 47.025 52.705 48.985 52.935 ;
        RECT 50.655 52.345 52.615 52.935 ;
        RECT 52.945 52.705 54.905 52.935 ;
        RECT 55.235 52.705 57.195 52.935 ;
        RECT 57.525 52.345 59.485 52.935 ;
        RECT 59.815 52.345 61.775 52.935 ;
        RECT 62.105 52.705 64.065 52.935 ;
        RECT 64.395 52.705 66.355 52.935 ;
        RECT 66.685 52.345 68.645 52.935 ;
        RECT 70.315 52.345 72.275 52.935 ;
        RECT 72.605 52.705 74.565 52.935 ;
        RECT 74.895 52.705 76.855 52.935 ;
        RECT 77.185 52.345 79.145 52.935 ;
        RECT 79.475 52.345 81.435 52.935 ;
        RECT 81.765 52.705 83.725 52.935 ;
        RECT 84.055 52.705 86.015 52.935 ;
        RECT 86.345 52.345 88.305 52.935 ;
        RECT 89.975 52.705 91.935 52.935 ;
        RECT 92.265 52.345 94.225 52.935 ;
        RECT 94.555 52.345 96.515 52.935 ;
        RECT 96.845 52.705 98.805 52.935 ;
        RECT 99.135 52.705 101.095 52.935 ;
        RECT 101.425 52.345 103.385 52.935 ;
        RECT 103.715 52.345 105.675 52.935 ;
        RECT 106.005 52.705 107.965 52.935 ;
        RECT 30.995 51.325 32.955 51.555 ;
        RECT 33.285 51.325 35.245 51.555 ;
        RECT 35.575 51.325 37.535 51.555 ;
        RECT 37.865 51.325 39.825 51.555 ;
        RECT 40.155 51.325 42.115 51.555 ;
        RECT 42.445 51.325 44.405 51.555 ;
        RECT 44.735 51.325 46.695 51.555 ;
        RECT 47.025 51.325 48.985 51.555 ;
        RECT 50.655 51.325 52.615 51.555 ;
        RECT 52.945 51.325 54.905 51.555 ;
        RECT 55.235 51.325 57.195 51.555 ;
        RECT 57.525 51.325 59.485 51.555 ;
        RECT 59.815 51.325 61.775 51.555 ;
        RECT 62.105 51.325 64.065 51.555 ;
        RECT 64.395 51.325 66.355 51.555 ;
        RECT 66.685 51.325 68.645 51.555 ;
        RECT 70.315 51.325 72.275 51.555 ;
        RECT 72.605 51.325 74.565 51.555 ;
        RECT 74.895 51.325 76.855 51.555 ;
        RECT 77.185 51.325 79.145 51.555 ;
        RECT 79.475 51.325 81.435 51.555 ;
        RECT 81.765 51.325 83.725 51.555 ;
        RECT 84.055 51.325 86.015 51.555 ;
        RECT 86.345 51.325 88.305 51.555 ;
        RECT 89.975 51.325 91.935 51.555 ;
        RECT 92.265 51.325 94.225 51.555 ;
        RECT 94.555 51.325 96.515 51.555 ;
        RECT 96.845 51.325 98.805 51.555 ;
        RECT 99.135 51.325 101.095 51.555 ;
        RECT 101.425 51.325 103.385 51.555 ;
        RECT 103.715 51.325 105.675 51.555 ;
        RECT 106.005 51.325 107.965 51.555 ;
        RECT 109.355 51.325 127.905 52.935 ;
        RECT 11.055 42.915 11.285 51.325 ;
        RECT 13.345 42.915 13.575 51.325 ;
        RECT 15.635 42.915 15.865 51.325 ;
        RECT 17.925 42.915 18.155 51.325 ;
        RECT 20.215 42.915 20.445 51.325 ;
        RECT 22.505 42.915 22.735 51.325 ;
        RECT 24.795 42.915 25.025 51.325 ;
        RECT 27.085 42.915 27.315 51.325 ;
        RECT 29.375 42.915 29.605 51.325 ;
        RECT 11.055 42.225 29.605 42.915 ;
        RECT 30.715 42.915 30.945 51.120 ;
        RECT 33.005 42.915 33.235 51.120 ;
        RECT 35.295 42.915 35.525 51.120 ;
        RECT 37.585 42.915 37.815 51.120 ;
        RECT 39.875 42.915 40.105 51.120 ;
        RECT 42.165 42.915 42.395 51.120 ;
        RECT 44.455 42.915 44.685 51.120 ;
        RECT 46.745 42.915 46.975 51.120 ;
        RECT 49.035 42.915 49.265 51.120 ;
        RECT 30.715 42.225 49.265 42.915 ;
        RECT 50.375 42.915 50.605 51.120 ;
        RECT 52.665 42.915 52.895 51.120 ;
        RECT 54.955 42.915 55.185 51.120 ;
        RECT 57.245 42.915 57.475 51.120 ;
        RECT 59.535 42.915 59.765 51.120 ;
        RECT 61.825 42.915 62.055 51.120 ;
        RECT 64.115 42.915 64.345 51.120 ;
        RECT 66.405 42.915 66.635 51.120 ;
        RECT 68.695 42.915 68.925 51.120 ;
        RECT 50.375 42.225 68.925 42.915 ;
        RECT 70.035 42.915 70.265 51.120 ;
        RECT 72.325 42.915 72.555 51.120 ;
        RECT 74.615 42.915 74.845 51.120 ;
        RECT 76.905 42.915 77.135 51.120 ;
        RECT 79.195 42.915 79.425 51.120 ;
        RECT 81.485 42.915 81.715 51.120 ;
        RECT 83.775 42.915 84.005 51.120 ;
        RECT 86.065 42.915 86.295 51.120 ;
        RECT 88.355 42.915 88.585 51.120 ;
        RECT 70.035 42.225 88.585 42.915 ;
        RECT 89.695 42.915 89.925 51.120 ;
        RECT 91.985 42.915 92.215 51.120 ;
        RECT 94.275 42.915 94.505 51.120 ;
        RECT 96.565 42.915 96.795 51.120 ;
        RECT 98.855 42.915 99.085 51.120 ;
        RECT 101.145 42.915 101.375 51.120 ;
        RECT 103.435 42.915 103.665 51.120 ;
        RECT 105.725 42.915 105.955 51.120 ;
        RECT 108.015 42.915 108.245 51.120 ;
        RECT 89.695 42.225 108.245 42.915 ;
        RECT 109.355 42.915 109.585 51.325 ;
        RECT 111.645 42.915 111.875 51.325 ;
        RECT 113.935 42.915 114.165 51.325 ;
        RECT 116.225 42.915 116.455 51.325 ;
        RECT 118.515 42.915 118.745 51.325 ;
        RECT 120.805 42.915 121.035 51.325 ;
        RECT 123.095 42.915 123.325 51.325 ;
        RECT 125.385 42.915 125.615 51.325 ;
        RECT 127.675 42.915 127.905 51.325 ;
        RECT 109.355 42.225 127.905 42.915 ;
        RECT 128.345 42.225 135.710 102.115 ;
        RECT 136.295 100.155 138.400 101.915 ;
        RECT 136.295 97.815 138.400 99.575 ;
        RECT 136.295 95.475 138.400 97.235 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 141.695 93.725 142.995 108.925 ;
        RECT 149.570 107.765 155.900 137.690 ;
        RECT 235.765 109.725 236.085 109.785 ;
        RECT 261.065 109.725 261.385 109.785 ;
        RECT 235.765 109.585 261.385 109.725 ;
        RECT 235.765 109.525 236.085 109.585 ;
        RECT 261.065 109.525 261.385 109.585 ;
        RECT 242.665 109.385 242.985 109.445 ;
        RECT 282.225 109.385 282.545 109.445 ;
        RECT 242.665 109.245 282.545 109.385 ;
        RECT 242.665 109.185 242.985 109.245 ;
        RECT 282.225 109.185 282.545 109.245 ;
        RECT 245.425 109.045 245.745 109.105 ;
        RECT 289.125 109.045 289.445 109.105 ;
        RECT 245.425 108.905 289.445 109.045 ;
        RECT 245.425 108.845 245.745 108.905 ;
        RECT 289.125 108.845 289.445 108.905 ;
        RECT 246.345 108.705 246.665 108.765 ;
        RECT 228.495 108.565 246.665 108.705 ;
        RECT 215.985 108.365 216.305 108.425 ;
        RECT 221.505 108.365 221.825 108.425 ;
        RECT 215.985 108.225 221.825 108.365 ;
        RECT 215.985 108.165 216.305 108.225 ;
        RECT 221.505 108.165 221.825 108.225 ;
        RECT 214.145 108.025 214.465 108.085 ;
        RECT 228.495 108.025 228.635 108.565 ;
        RECT 246.345 108.505 246.665 108.565 ;
        RECT 252.785 108.705 253.105 108.765 ;
        RECT 292.345 108.705 292.665 108.765 ;
        RECT 252.785 108.565 292.665 108.705 ;
        RECT 252.785 108.505 253.105 108.565 ;
        RECT 292.345 108.505 292.665 108.565 ;
        RECT 228.865 108.365 229.185 108.425 ;
        RECT 252.325 108.365 252.645 108.425 ;
        RECT 272.565 108.365 272.885 108.425 ;
        RECT 304.765 108.365 305.085 108.425 ;
        RECT 228.865 108.225 252.645 108.365 ;
        RECT 228.865 108.165 229.185 108.225 ;
        RECT 252.325 108.165 252.645 108.225 ;
        RECT 257.015 108.225 305.085 108.365 ;
        RECT 214.145 107.885 228.635 108.025 ;
        RECT 238.985 108.025 239.305 108.085 ;
        RECT 256.465 108.025 256.785 108.085 ;
        RECT 238.985 107.885 256.785 108.025 ;
        RECT 214.145 107.825 214.465 107.885 ;
        RECT 238.985 107.825 239.305 107.885 ;
        RECT 256.465 107.825 256.785 107.885 ;
        RECT 146.290 104.835 155.900 107.765 ;
        RECT 169.525 107.685 169.845 107.745 ;
        RECT 187.005 107.685 187.325 107.745 ;
        RECT 169.525 107.545 187.325 107.685 ;
        RECT 169.525 107.485 169.845 107.545 ;
        RECT 187.005 107.485 187.325 107.545 ;
        RECT 204.945 107.685 205.265 107.745 ;
        RECT 216.905 107.685 217.225 107.745 ;
        RECT 253.245 107.685 253.565 107.745 ;
        RECT 257.015 107.685 257.155 108.225 ;
        RECT 272.565 108.165 272.885 108.225 ;
        RECT 304.765 108.165 305.085 108.225 ;
        RECT 271.645 108.025 271.965 108.085 ;
        RECT 307.985 108.025 308.305 108.085 ;
        RECT 271.645 107.885 308.305 108.025 ;
        RECT 271.645 107.825 271.965 107.885 ;
        RECT 307.985 107.825 308.305 107.885 ;
        RECT 204.945 107.545 217.225 107.685 ;
        RECT 204.945 107.485 205.265 107.545 ;
        RECT 216.905 107.485 217.225 107.545 ;
        RECT 221.365 107.545 257.155 107.685 ;
        RECT 262.905 107.685 263.225 107.745 ;
        RECT 275.785 107.685 276.105 107.745 ;
        RECT 262.905 107.545 276.105 107.685 ;
        RECT 178.265 107.345 178.585 107.405 ;
        RECT 197.585 107.345 197.905 107.405 ;
        RECT 208.625 107.345 208.945 107.405 ;
        RECT 221.365 107.345 221.505 107.545 ;
        RECT 253.245 107.485 253.565 107.545 ;
        RECT 262.905 107.485 263.225 107.545 ;
        RECT 275.785 107.485 276.105 107.545 ;
        RECT 178.265 107.205 221.505 107.345 ;
        RECT 244.965 107.345 245.285 107.405 ;
        RECT 248.185 107.345 248.505 107.405 ;
        RECT 257.385 107.345 257.705 107.405 ;
        RECT 244.965 107.205 257.705 107.345 ;
        RECT 178.265 107.145 178.585 107.205 ;
        RECT 197.585 107.145 197.905 107.205 ;
        RECT 208.625 107.145 208.945 107.205 ;
        RECT 244.965 107.145 245.285 107.205 ;
        RECT 248.185 107.145 248.505 107.205 ;
        RECT 257.385 107.145 257.705 107.205 ;
        RECT 260.605 107.345 260.925 107.405 ;
        RECT 273.485 107.345 273.805 107.405 ;
        RECT 260.605 107.205 273.805 107.345 ;
        RECT 260.605 107.145 260.925 107.205 ;
        RECT 273.485 107.145 273.805 107.205 ;
        RECT 279.005 107.345 279.325 107.405 ;
        RECT 283.145 107.345 283.465 107.405 ;
        RECT 279.005 107.205 283.465 107.345 ;
        RECT 279.005 107.145 279.325 107.205 ;
        RECT 283.145 107.145 283.465 107.205 ;
        RECT 289.125 107.345 289.445 107.405 ;
        RECT 303.385 107.345 303.705 107.405 ;
        RECT 289.125 107.205 303.705 107.345 ;
        RECT 289.125 107.145 289.445 107.205 ;
        RECT 303.385 107.145 303.705 107.205 ;
        RECT 187.005 107.005 187.325 107.065 ;
        RECT 196.205 107.005 196.525 107.065 ;
        RECT 187.005 106.865 196.525 107.005 ;
        RECT 187.005 106.805 187.325 106.865 ;
        RECT 196.205 106.805 196.525 106.865 ;
        RECT 216.905 107.005 217.225 107.065 ;
        RECT 229.785 107.005 230.105 107.065 ;
        RECT 216.905 106.865 230.105 107.005 ;
        RECT 216.905 106.805 217.225 106.865 ;
        RECT 229.785 106.805 230.105 106.865 ;
        RECT 242.205 107.005 242.525 107.065 ;
        RECT 255.545 107.005 255.865 107.065 ;
        RECT 242.205 106.865 255.865 107.005 ;
        RECT 242.205 106.805 242.525 106.865 ;
        RECT 255.545 106.805 255.865 106.865 ;
        RECT 256.005 107.005 256.325 107.065 ;
        RECT 260.145 107.005 260.465 107.065 ;
        RECT 256.005 106.865 260.465 107.005 ;
        RECT 256.005 106.805 256.325 106.865 ;
        RECT 260.145 106.805 260.465 106.865 ;
        RECT 261.065 107.005 261.385 107.065 ;
        RECT 271.645 107.005 271.965 107.065 ;
        RECT 261.065 106.865 271.965 107.005 ;
        RECT 261.065 106.805 261.385 106.865 ;
        RECT 271.645 106.805 271.965 106.865 ;
        RECT 272.105 107.005 272.425 107.065 ;
        RECT 282.685 107.005 283.005 107.065 ;
        RECT 272.105 106.865 283.005 107.005 ;
        RECT 272.105 106.805 272.425 106.865 ;
        RECT 282.685 106.805 283.005 106.865 ;
        RECT 292.805 107.005 293.125 107.065 ;
        RECT 307.065 107.005 307.385 107.065 ;
        RECT 292.805 106.865 307.385 107.005 ;
        RECT 292.805 106.805 293.125 106.865 ;
        RECT 307.065 106.805 307.385 106.865 ;
        RECT 162.095 106.185 311.135 106.665 ;
        RECT 164.020 105.985 164.310 106.030 ;
        RECT 173.205 105.985 173.525 106.045 ;
        RECT 164.020 105.845 173.525 105.985 ;
        RECT 164.020 105.800 164.310 105.845 ;
        RECT 173.205 105.785 173.525 105.845 ;
        RECT 181.500 105.985 181.790 106.030 ;
        RECT 189.305 105.985 189.625 106.045 ;
        RECT 181.500 105.845 189.625 105.985 ;
        RECT 181.500 105.800 181.790 105.845 ;
        RECT 189.305 105.785 189.625 105.845 ;
        RECT 189.765 105.985 190.085 106.045 ;
        RECT 191.160 105.985 191.450 106.030 ;
        RECT 194.380 105.985 194.670 106.030 ;
        RECT 198.505 105.985 198.825 106.045 ;
        RECT 189.765 105.845 192.295 105.985 ;
        RECT 189.765 105.785 190.085 105.845 ;
        RECT 191.160 105.800 191.450 105.845 ;
        RECT 177.805 105.645 178.125 105.705 ;
        RECT 170.075 105.505 178.125 105.645 ;
        RECT 164.465 105.305 164.785 105.365 ;
        RECT 164.940 105.305 165.230 105.350 ;
        RECT 164.465 105.165 165.230 105.305 ;
        RECT 164.465 105.105 164.785 105.165 ;
        RECT 164.940 105.120 165.230 105.165 ;
        RECT 166.780 105.305 167.070 105.350 ;
        RECT 167.225 105.305 167.545 105.365 ;
        RECT 166.780 105.165 167.545 105.305 ;
        RECT 166.780 105.120 167.070 105.165 ;
        RECT 167.225 105.105 167.545 105.165 ;
        RECT 168.620 105.305 168.910 105.350 ;
        RECT 169.065 105.305 169.385 105.365 ;
        RECT 168.620 105.165 169.385 105.305 ;
        RECT 168.620 105.120 168.910 105.165 ;
        RECT 169.065 105.105 169.385 105.165 ;
        RECT 170.075 104.965 170.215 105.505 ;
        RECT 177.805 105.445 178.125 105.505 ;
        RECT 181.025 105.645 181.345 105.705 ;
        RECT 191.605 105.645 191.925 105.705 ;
        RECT 181.025 105.505 182.635 105.645 ;
        RECT 181.025 105.445 181.345 105.505 ;
        RECT 170.460 105.305 170.750 105.350 ;
        RECT 172.760 105.305 173.050 105.350 ;
        RECT 173.665 105.305 173.985 105.365 ;
        RECT 182.495 105.350 182.635 105.505 ;
        RECT 187.555 105.505 191.925 105.645 ;
        RECT 192.155 105.645 192.295 105.845 ;
        RECT 194.380 105.845 198.825 105.985 ;
        RECT 194.380 105.800 194.670 105.845 ;
        RECT 198.505 105.785 198.825 105.845 ;
        RECT 199.900 105.985 200.190 106.030 ;
        RECT 207.705 105.985 208.025 106.045 ;
        RECT 212.320 105.985 212.610 106.030 ;
        RECT 199.900 105.845 208.025 105.985 ;
        RECT 199.900 105.800 200.190 105.845 ;
        RECT 207.705 105.785 208.025 105.845 ;
        RECT 208.255 105.845 209.315 105.985 ;
        RECT 208.255 105.645 208.395 105.845 ;
        RECT 192.155 105.505 208.395 105.645 ;
        RECT 177.360 105.305 177.650 105.350 ;
        RECT 180.580 105.305 180.870 105.350 ;
        RECT 170.460 105.165 173.985 105.305 ;
        RECT 170.460 105.120 170.750 105.165 ;
        RECT 172.760 105.120 173.050 105.165 ;
        RECT 173.665 105.105 173.985 105.165 ;
        RECT 174.215 105.165 177.115 105.305 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 146.290 101.325 148.395 103.085 ;
        RECT 146.290 98.985 148.395 100.745 ;
        RECT 146.290 96.645 148.395 98.405 ;
        RECT 146.290 94.305 148.395 96.065 ;
        RECT 136.295 91.965 138.400 93.725 ;
        RECT 141.695 93.135 148.395 93.725 ;
        RECT 146.290 91.965 148.395 92.555 ;
        RECT 136.295 90.795 143.395 91.385 ;
        RECT 136.295 89.625 138.400 90.215 ;
        RECT 146.290 89.625 148.395 91.385 ;
        RECT 136.295 87.285 138.400 89.045 ;
        RECT 146.290 88.455 148.395 89.045 ;
        RECT 146.290 87.285 148.395 87.875 ;
        RECT 136.295 86.115 138.400 86.705 ;
        RECT 136.295 84.945 138.400 85.535 ;
        RECT 146.290 84.945 148.395 86.705 ;
        RECT 136.295 82.605 138.400 84.365 ;
        RECT 146.290 83.775 148.395 84.365 ;
        RECT 146.290 82.605 148.395 83.195 ;
        RECT 136.295 81.435 141.260 82.025 ;
        RECT 143.790 81.435 148.395 82.025 ;
        RECT 136.295 80.265 138.400 80.855 ;
        RECT 136.295 79.095 138.400 79.685 ;
        RECT 136.295 76.755 138.400 78.515 ;
        RECT 136.295 75.585 138.400 76.175 ;
        RECT 136.295 74.415 138.400 75.005 ;
        RECT 136.295 72.075 138.400 73.835 ;
        RECT 136.295 70.905 138.400 71.495 ;
        RECT 136.295 69.735 138.400 70.325 ;
        RECT 136.295 67.395 138.400 69.155 ;
        RECT 136.295 66.225 138.400 66.815 ;
        RECT 136.295 65.055 138.400 65.645 ;
        RECT 136.295 62.715 138.400 64.475 ;
        RECT 143.790 62.135 145.190 81.435 ;
        RECT 146.290 79.095 148.395 80.855 ;
        RECT 146.290 77.925 148.395 78.515 ;
        RECT 146.290 76.755 148.395 77.345 ;
        RECT 146.290 74.415 148.395 76.175 ;
        RECT 146.290 73.245 148.395 73.835 ;
        RECT 146.290 72.075 148.395 72.665 ;
        RECT 146.290 69.735 148.395 71.495 ;
        RECT 146.290 68.565 148.395 69.155 ;
        RECT 146.290 67.395 148.395 67.985 ;
        RECT 146.290 65.055 148.395 66.815 ;
        RECT 146.290 63.885 148.395 64.475 ;
        RECT 146.290 62.715 148.395 63.305 ;
        RECT 136.295 61.545 140.910 62.135 ;
        RECT 143.790 61.545 148.395 62.135 ;
        RECT 136.295 60.375 138.400 60.965 ;
        RECT 136.295 59.205 138.400 59.795 ;
        RECT 136.295 56.865 138.400 58.625 ;
        RECT 136.295 55.695 138.400 56.285 ;
        RECT 136.295 54.525 138.400 55.115 ;
        RECT 136.295 52.185 138.400 53.945 ;
        RECT 136.295 51.015 138.400 51.605 ;
        RECT 136.295 49.845 138.400 50.435 ;
        RECT 136.295 47.505 138.400 49.265 ;
        RECT 136.295 46.335 138.400 46.925 ;
        RECT 136.295 45.165 138.400 45.755 ;
        RECT 136.295 42.825 138.400 44.585 ;
        RECT 139.510 42.245 140.910 61.545 ;
        RECT 146.290 59.205 148.395 60.965 ;
        RECT 146.290 58.035 148.395 58.625 ;
        RECT 146.290 56.865 148.395 57.455 ;
        RECT 146.290 54.525 148.395 56.285 ;
        RECT 146.290 53.355 148.395 53.945 ;
        RECT 146.290 52.185 148.395 52.775 ;
        RECT 146.290 49.845 148.395 51.605 ;
        RECT 146.290 48.675 148.395 49.265 ;
        RECT 146.290 47.505 148.395 48.095 ;
        RECT 146.290 45.165 148.395 46.925 ;
        RECT 146.290 43.995 148.395 44.585 ;
        RECT 146.290 42.825 148.395 43.415 ;
        RECT 4.100 41.635 135.710 42.225 ;
        RECT 136.295 41.655 140.910 42.245 ;
        RECT 143.435 41.655 148.395 42.245 ;
        RECT 4.100 4.900 4.900 41.635 ;
        RECT 7.065 39.040 130.565 39.630 ;
        RECT 7.065 36.430 10.615 39.040 ;
        RECT 8.665 9.480 10.615 36.430 ;
        RECT 11.115 38.350 20.505 38.580 ;
        RECT 22.015 38.350 30.845 38.650 ;
        RECT 32.635 38.350 41.465 38.650 ;
        RECT 43.255 38.350 52.085 38.650 ;
        RECT 53.875 38.350 62.705 38.650 ;
        RECT 64.215 38.350 73.605 38.580 ;
        RECT 11.115 34.890 11.345 38.350 ;
        RECT 13.405 34.890 13.635 38.190 ;
        RECT 15.695 34.890 15.925 38.350 ;
        RECT 17.985 34.890 18.215 38.190 ;
        RECT 20.275 34.890 20.505 38.350 ;
        RECT 11.020 33.490 11.345 34.890 ;
        RECT 13.370 33.490 13.670 34.890 ;
        RECT 15.660 33.490 15.960 34.890 ;
        RECT 17.950 33.490 18.250 34.890 ;
        RECT 20.240 33.490 20.540 34.890 ;
        RECT 11.115 30.030 11.345 33.490 ;
        RECT 13.405 30.190 13.635 33.490 ;
        RECT 15.695 30.030 15.925 33.490 ;
        RECT 17.985 30.190 18.215 33.490 ;
        RECT 20.275 30.030 20.505 33.490 ;
        RECT 21.735 32.890 21.965 38.190 ;
        RECT 24.025 34.890 24.255 38.190 ;
        RECT 26.315 36.890 26.545 38.190 ;
        RECT 26.280 35.490 26.580 36.890 ;
        RECT 23.990 33.490 24.290 34.890 ;
        RECT 21.700 31.490 22.000 32.890 ;
        RECT 21.735 30.190 21.965 31.490 ;
        RECT 24.025 30.190 24.255 33.490 ;
        RECT 26.315 30.190 26.545 35.490 ;
        RECT 28.605 34.890 28.835 38.190 ;
        RECT 28.570 33.490 28.870 34.890 ;
        RECT 28.605 30.190 28.835 33.490 ;
        RECT 30.895 32.890 31.125 38.190 ;
        RECT 32.355 36.890 32.585 38.190 ;
        RECT 32.320 35.490 32.620 36.890 ;
        RECT 30.860 31.490 31.160 32.890 ;
        RECT 30.895 30.190 31.125 31.490 ;
        RECT 32.355 30.190 32.585 35.490 ;
        RECT 34.645 34.890 34.875 38.190 ;
        RECT 34.610 33.490 34.910 34.890 ;
        RECT 34.645 30.190 34.875 33.490 ;
        RECT 36.935 32.890 37.165 38.190 ;
        RECT 39.225 34.890 39.455 38.190 ;
        RECT 41.515 36.890 41.745 38.190 ;
        RECT 41.480 35.490 41.780 36.890 ;
        RECT 39.190 33.490 39.490 34.890 ;
        RECT 36.900 31.490 37.200 32.890 ;
        RECT 36.935 30.190 37.165 31.490 ;
        RECT 39.225 30.190 39.455 33.490 ;
        RECT 41.515 30.190 41.745 35.490 ;
        RECT 42.975 32.890 43.205 38.190 ;
        RECT 45.265 34.890 45.495 38.190 ;
        RECT 47.555 36.890 47.785 38.190 ;
        RECT 47.520 35.490 47.820 36.890 ;
        RECT 45.230 33.490 45.530 34.890 ;
        RECT 42.940 31.490 43.240 32.890 ;
        RECT 42.975 30.190 43.205 31.490 ;
        RECT 45.265 30.190 45.495 33.490 ;
        RECT 47.555 30.190 47.785 35.490 ;
        RECT 49.845 34.890 50.075 38.190 ;
        RECT 49.810 33.490 50.110 34.890 ;
        RECT 49.845 30.190 50.075 33.490 ;
        RECT 52.135 32.890 52.365 38.190 ;
        RECT 53.595 36.890 53.825 38.190 ;
        RECT 53.560 35.490 53.860 36.890 ;
        RECT 52.100 31.490 52.400 32.890 ;
        RECT 52.135 30.190 52.365 31.490 ;
        RECT 53.595 30.190 53.825 35.490 ;
        RECT 55.885 34.890 56.115 38.190 ;
        RECT 55.850 33.490 56.150 34.890 ;
        RECT 55.885 30.190 56.115 33.490 ;
        RECT 58.175 32.890 58.405 38.190 ;
        RECT 60.465 34.890 60.695 38.190 ;
        RECT 62.755 36.890 62.985 38.190 ;
        RECT 62.720 35.490 63.020 36.890 ;
        RECT 60.430 33.490 60.730 34.890 ;
        RECT 58.140 31.490 58.440 32.890 ;
        RECT 58.175 30.190 58.405 31.490 ;
        RECT 60.465 30.190 60.695 33.490 ;
        RECT 62.755 30.190 62.985 35.490 ;
        RECT 64.215 34.890 64.445 38.350 ;
        RECT 66.505 34.890 66.735 38.190 ;
        RECT 68.795 34.890 69.025 38.350 ;
        RECT 71.085 34.890 71.315 38.190 ;
        RECT 73.375 34.890 73.605 38.350 ;
        RECT 64.180 33.490 64.480 34.890 ;
        RECT 66.470 33.490 66.770 34.890 ;
        RECT 68.760 33.490 69.060 34.890 ;
        RECT 71.050 33.490 71.350 34.890 ;
        RECT 73.340 33.490 73.640 34.890 ;
        RECT 64.215 30.030 64.445 33.490 ;
        RECT 66.505 30.190 66.735 33.490 ;
        RECT 68.795 30.030 69.025 33.490 ;
        RECT 71.085 30.190 71.315 33.490 ;
        RECT 73.375 30.030 73.605 33.490 ;
        RECT 11.115 29.800 20.505 30.030 ;
        RECT 22.015 29.730 30.845 30.030 ;
        RECT 32.635 29.730 41.465 30.030 ;
        RECT 43.255 29.730 52.085 30.030 ;
        RECT 53.875 29.730 62.705 30.030 ;
        RECT 64.215 29.800 73.605 30.030 ;
        RECT 11.115 28.420 20.505 28.650 ;
        RECT 22.015 28.420 30.845 28.720 ;
        RECT 32.635 28.650 41.465 28.720 ;
        RECT 43.255 28.650 52.085 28.720 ;
        RECT 32.355 28.420 41.745 28.650 ;
        RECT 11.115 24.960 11.345 28.420 ;
        RECT 13.405 24.960 13.635 28.260 ;
        RECT 15.695 24.960 15.925 28.420 ;
        RECT 17.985 24.960 18.215 28.260 ;
        RECT 20.275 24.960 20.505 28.420 ;
        RECT 21.735 26.960 21.965 28.260 ;
        RECT 21.700 25.560 22.000 26.960 ;
        RECT 11.020 23.560 11.345 24.960 ;
        RECT 13.370 23.560 13.670 24.960 ;
        RECT 15.660 23.560 15.960 24.960 ;
        RECT 17.950 23.560 18.250 24.960 ;
        RECT 20.240 23.560 20.540 24.960 ;
        RECT 11.115 20.100 11.345 23.560 ;
        RECT 13.405 20.260 13.635 23.560 ;
        RECT 15.695 20.100 15.925 23.560 ;
        RECT 17.985 20.260 18.215 23.560 ;
        RECT 20.275 20.100 20.505 23.560 ;
        RECT 21.735 20.260 21.965 25.560 ;
        RECT 24.025 24.960 24.255 28.260 ;
        RECT 23.990 23.560 24.290 24.960 ;
        RECT 24.025 20.260 24.255 23.560 ;
        RECT 26.315 22.960 26.545 28.260 ;
        RECT 28.605 24.960 28.835 28.260 ;
        RECT 30.895 26.960 31.125 28.260 ;
        RECT 30.860 25.560 31.160 26.960 ;
        RECT 28.570 23.560 28.870 24.960 ;
        RECT 26.280 21.560 26.580 22.960 ;
        RECT 26.315 20.260 26.545 21.560 ;
        RECT 28.605 20.260 28.835 23.560 ;
        RECT 30.895 20.260 31.125 25.560 ;
        RECT 32.355 20.100 32.585 28.420 ;
        RECT 34.645 24.960 34.875 28.260 ;
        RECT 34.610 23.560 34.910 24.960 ;
        RECT 34.645 20.260 34.875 23.560 ;
        RECT 36.935 20.100 37.165 28.420 ;
        RECT 39.225 24.960 39.455 28.260 ;
        RECT 39.190 23.560 39.490 24.960 ;
        RECT 39.225 20.260 39.455 23.560 ;
        RECT 41.515 20.100 41.745 28.420 ;
        RECT 11.115 19.870 20.505 20.100 ;
        RECT 22.015 19.800 30.845 20.100 ;
        RECT 32.355 19.870 41.745 20.100 ;
        RECT 42.975 28.420 52.365 28.650 ;
        RECT 53.875 28.420 62.705 28.720 ;
        RECT 64.215 28.420 73.605 28.650 ;
        RECT 42.975 20.100 43.205 28.420 ;
        RECT 45.265 24.960 45.495 28.260 ;
        RECT 45.230 23.560 45.530 24.960 ;
        RECT 45.265 20.260 45.495 23.560 ;
        RECT 47.555 20.100 47.785 28.420 ;
        RECT 49.845 24.960 50.075 28.260 ;
        RECT 49.810 23.560 50.110 24.960 ;
        RECT 49.845 20.260 50.075 23.560 ;
        RECT 52.135 20.100 52.365 28.420 ;
        RECT 53.595 22.960 53.825 28.260 ;
        RECT 55.885 24.960 56.115 28.260 ;
        RECT 58.175 26.960 58.405 28.260 ;
        RECT 58.140 25.560 58.440 26.960 ;
        RECT 55.850 23.560 56.150 24.960 ;
        RECT 53.560 21.560 53.860 22.960 ;
        RECT 53.595 20.260 53.825 21.560 ;
        RECT 55.885 20.260 56.115 23.560 ;
        RECT 58.175 20.260 58.405 25.560 ;
        RECT 60.465 24.960 60.695 28.260 ;
        RECT 60.430 23.560 60.730 24.960 ;
        RECT 60.465 20.260 60.695 23.560 ;
        RECT 62.755 22.960 62.985 28.260 ;
        RECT 64.215 24.960 64.445 28.420 ;
        RECT 66.505 24.960 66.735 28.260 ;
        RECT 68.795 24.960 69.025 28.420 ;
        RECT 71.085 24.960 71.315 28.260 ;
        RECT 73.375 24.960 73.605 28.420 ;
        RECT 64.180 23.560 64.480 24.960 ;
        RECT 66.470 23.560 66.770 24.960 ;
        RECT 68.760 23.560 69.060 24.960 ;
        RECT 71.050 23.560 71.350 24.960 ;
        RECT 73.340 23.560 73.640 24.960 ;
        RECT 62.720 21.560 63.020 22.960 ;
        RECT 62.755 20.260 62.985 21.560 ;
        RECT 64.215 20.100 64.445 23.560 ;
        RECT 66.505 20.260 66.735 23.560 ;
        RECT 68.795 20.100 69.025 23.560 ;
        RECT 71.085 20.260 71.315 23.560 ;
        RECT 73.375 20.100 73.605 23.560 ;
        RECT 42.975 19.870 52.365 20.100 ;
        RECT 32.635 19.800 41.465 19.870 ;
        RECT 43.255 19.800 52.085 19.870 ;
        RECT 53.875 19.800 62.705 20.100 ;
        RECT 64.215 19.870 73.605 20.100 ;
        RECT 11.115 18.490 20.505 18.720 ;
        RECT 22.015 18.490 30.845 18.790 ;
        RECT 32.635 18.490 41.465 18.790 ;
        RECT 43.255 18.490 52.085 18.790 ;
        RECT 53.875 18.490 62.705 18.790 ;
        RECT 64.215 18.490 73.605 18.720 ;
        RECT 11.115 15.030 11.345 18.490 ;
        RECT 13.405 15.030 13.635 18.330 ;
        RECT 15.695 15.030 15.925 18.490 ;
        RECT 17.985 15.030 18.215 18.330 ;
        RECT 20.275 15.030 20.505 18.490 ;
        RECT 11.020 13.630 11.345 15.030 ;
        RECT 13.370 13.630 13.670 15.030 ;
        RECT 15.660 13.630 15.960 15.030 ;
        RECT 17.950 13.630 18.250 15.030 ;
        RECT 20.240 13.630 20.540 15.030 ;
        RECT 11.115 10.170 11.345 13.630 ;
        RECT 13.405 10.330 13.635 13.630 ;
        RECT 15.695 10.170 15.925 13.630 ;
        RECT 17.985 10.330 18.215 13.630 ;
        RECT 20.275 10.170 20.505 13.630 ;
        RECT 21.735 13.030 21.965 18.330 ;
        RECT 24.025 15.030 24.255 18.330 ;
        RECT 26.315 17.030 26.545 18.330 ;
        RECT 26.280 15.630 26.580 17.030 ;
        RECT 23.990 13.630 24.290 15.030 ;
        RECT 21.700 11.630 22.000 13.030 ;
        RECT 21.735 10.330 21.965 11.630 ;
        RECT 24.025 10.330 24.255 13.630 ;
        RECT 26.315 10.330 26.545 15.630 ;
        RECT 28.605 15.030 28.835 18.330 ;
        RECT 28.570 13.630 28.870 15.030 ;
        RECT 28.605 10.330 28.835 13.630 ;
        RECT 30.895 13.030 31.125 18.330 ;
        RECT 32.355 17.030 32.585 18.330 ;
        RECT 32.320 15.630 32.620 17.030 ;
        RECT 30.860 11.630 31.160 13.030 ;
        RECT 30.895 10.330 31.125 11.630 ;
        RECT 32.355 10.330 32.585 15.630 ;
        RECT 34.645 15.030 34.875 18.330 ;
        RECT 34.610 13.630 34.910 15.030 ;
        RECT 34.645 10.330 34.875 13.630 ;
        RECT 36.935 13.030 37.165 18.330 ;
        RECT 39.225 15.030 39.455 18.330 ;
        RECT 41.515 17.030 41.745 18.330 ;
        RECT 41.480 15.630 41.780 17.030 ;
        RECT 39.190 13.630 39.490 15.030 ;
        RECT 36.900 11.630 37.200 13.030 ;
        RECT 36.935 10.330 37.165 11.630 ;
        RECT 39.225 10.330 39.455 13.630 ;
        RECT 41.515 10.330 41.745 15.630 ;
        RECT 42.975 13.030 43.205 18.330 ;
        RECT 45.265 15.030 45.495 18.330 ;
        RECT 47.555 17.030 47.785 18.330 ;
        RECT 47.520 15.630 47.820 17.030 ;
        RECT 45.230 13.630 45.530 15.030 ;
        RECT 42.940 11.630 43.240 13.030 ;
        RECT 42.975 10.330 43.205 11.630 ;
        RECT 45.265 10.330 45.495 13.630 ;
        RECT 47.555 10.330 47.785 15.630 ;
        RECT 49.845 15.030 50.075 18.330 ;
        RECT 49.810 13.630 50.110 15.030 ;
        RECT 49.845 10.330 50.075 13.630 ;
        RECT 52.135 13.030 52.365 18.330 ;
        RECT 53.595 17.030 53.825 18.330 ;
        RECT 53.560 15.630 53.860 17.030 ;
        RECT 52.100 11.630 52.400 13.030 ;
        RECT 52.135 10.330 52.365 11.630 ;
        RECT 53.595 10.330 53.825 15.630 ;
        RECT 55.885 15.030 56.115 18.330 ;
        RECT 55.850 13.630 56.150 15.030 ;
        RECT 55.885 10.330 56.115 13.630 ;
        RECT 58.175 13.030 58.405 18.330 ;
        RECT 60.465 15.030 60.695 18.330 ;
        RECT 62.755 17.030 62.985 18.330 ;
        RECT 62.720 15.630 63.020 17.030 ;
        RECT 60.430 13.630 60.730 15.030 ;
        RECT 58.140 11.630 58.440 13.030 ;
        RECT 58.175 10.330 58.405 11.630 ;
        RECT 60.465 10.330 60.695 13.630 ;
        RECT 62.755 10.330 62.985 15.630 ;
        RECT 64.215 15.030 64.445 18.490 ;
        RECT 66.505 15.030 66.735 18.330 ;
        RECT 68.795 15.030 69.025 18.490 ;
        RECT 71.085 15.030 71.315 18.330 ;
        RECT 73.375 15.030 73.605 18.490 ;
        RECT 64.180 13.630 64.480 15.030 ;
        RECT 66.470 13.630 66.770 15.030 ;
        RECT 68.760 13.630 69.060 15.030 ;
        RECT 71.050 13.630 71.350 15.030 ;
        RECT 73.340 13.630 73.640 15.030 ;
        RECT 64.215 10.170 64.445 13.630 ;
        RECT 66.505 10.330 66.735 13.630 ;
        RECT 68.795 10.170 69.025 13.630 ;
        RECT 71.085 10.330 71.315 13.630 ;
        RECT 73.375 10.170 73.605 13.630 ;
        RECT 11.115 9.940 20.505 10.170 ;
        RECT 22.015 9.870 30.845 10.170 ;
        RECT 32.635 9.870 41.465 10.170 ;
        RECT 43.255 9.870 52.085 10.170 ;
        RECT 53.875 9.870 62.705 10.170 ;
        RECT 64.215 9.940 73.605 10.170 ;
        RECT 74.105 9.480 80.255 39.040 ;
        RECT 81.035 38.350 82.995 38.580 ;
        RECT 83.325 38.350 85.285 38.580 ;
        RECT 87.075 38.350 89.035 38.700 ;
        RECT 89.365 38.350 91.325 38.700 ;
        RECT 93.115 38.350 97.365 38.700 ;
        RECT 99.155 38.350 101.115 38.700 ;
        RECT 101.445 38.350 103.405 38.700 ;
        RECT 105.195 38.350 107.155 38.700 ;
        RECT 107.485 38.350 109.445 38.700 ;
        RECT 111.235 38.350 115.485 38.700 ;
        RECT 117.275 38.350 119.235 38.700 ;
        RECT 119.565 38.350 121.525 38.700 ;
        RECT 123.315 38.350 125.275 38.580 ;
        RECT 125.605 38.350 127.565 38.580 ;
        RECT 80.755 30.190 80.985 38.190 ;
        RECT 83.045 30.190 83.275 38.190 ;
        RECT 85.335 30.190 85.565 38.190 ;
        RECT 86.795 35.995 87.025 38.190 ;
        RECT 86.560 35.295 87.260 35.995 ;
        RECT 86.795 30.190 87.025 35.295 ;
        RECT 89.085 34.495 89.315 38.190 ;
        RECT 91.375 35.995 91.605 38.190 ;
        RECT 92.835 37.495 93.065 38.190 ;
        RECT 92.600 36.795 93.300 37.495 ;
        RECT 91.140 35.295 91.840 35.995 ;
        RECT 88.850 33.795 89.550 34.495 ;
        RECT 89.085 30.190 89.315 33.795 ;
        RECT 91.375 30.190 91.605 35.295 ;
        RECT 92.835 30.190 93.065 36.795 ;
        RECT 95.125 30.190 95.355 38.350 ;
        RECT 97.415 37.495 97.645 38.190 ;
        RECT 97.180 36.795 97.880 37.495 ;
        RECT 97.415 30.190 97.645 36.795 ;
        RECT 98.875 31.495 99.105 38.190 ;
        RECT 101.165 32.995 101.395 38.190 ;
        RECT 100.930 32.295 101.630 32.995 ;
        RECT 98.640 30.795 99.340 31.495 ;
        RECT 98.875 30.190 99.105 30.795 ;
        RECT 101.165 30.190 101.395 32.295 ;
        RECT 103.455 31.495 103.685 38.190 ;
        RECT 104.915 31.495 105.145 38.190 ;
        RECT 107.205 32.995 107.435 38.190 ;
        RECT 106.970 32.295 107.670 32.995 ;
        RECT 103.220 30.795 103.920 31.495 ;
        RECT 104.680 30.795 105.380 31.495 ;
        RECT 103.455 30.190 103.685 30.795 ;
        RECT 104.915 30.190 105.145 30.795 ;
        RECT 107.205 30.190 107.435 32.295 ;
        RECT 109.495 31.495 109.725 38.190 ;
        RECT 110.955 37.495 111.185 38.190 ;
        RECT 110.720 36.795 111.420 37.495 ;
        RECT 109.260 30.795 109.960 31.495 ;
        RECT 109.495 30.190 109.725 30.795 ;
        RECT 110.955 30.190 111.185 36.795 ;
        RECT 113.245 30.190 113.475 38.350 ;
        RECT 115.535 37.495 115.765 38.190 ;
        RECT 115.300 36.795 116.000 37.495 ;
        RECT 115.535 30.190 115.765 36.795 ;
        RECT 116.995 35.995 117.225 38.190 ;
        RECT 116.760 35.295 117.460 35.995 ;
        RECT 116.995 30.190 117.225 35.295 ;
        RECT 119.285 34.495 119.515 38.190 ;
        RECT 121.575 35.995 121.805 38.190 ;
        RECT 121.340 35.295 122.040 35.995 ;
        RECT 119.050 33.795 119.750 34.495 ;
        RECT 119.285 30.190 119.515 33.795 ;
        RECT 121.575 30.190 121.805 35.295 ;
        RECT 123.035 30.190 123.265 38.190 ;
        RECT 125.325 30.190 125.555 38.190 ;
        RECT 127.615 30.190 127.845 38.190 ;
        RECT 81.035 29.800 82.995 30.030 ;
        RECT 83.325 29.800 85.285 30.030 ;
        RECT 87.075 29.680 89.035 30.030 ;
        RECT 89.365 29.680 91.325 30.030 ;
        RECT 93.115 29.680 95.075 30.030 ;
        RECT 95.405 29.680 97.365 30.030 ;
        RECT 99.155 29.680 101.115 30.030 ;
        RECT 101.445 29.680 103.405 30.030 ;
        RECT 105.195 29.680 107.155 30.030 ;
        RECT 107.485 29.680 109.445 30.030 ;
        RECT 111.235 29.680 113.195 30.030 ;
        RECT 113.525 29.680 115.485 30.030 ;
        RECT 117.275 29.680 119.235 30.030 ;
        RECT 119.565 29.680 121.525 30.030 ;
        RECT 123.315 29.800 125.275 30.030 ;
        RECT 125.605 29.800 127.565 30.030 ;
        RECT 81.035 28.420 82.995 28.650 ;
        RECT 83.325 28.420 85.285 28.650 ;
        RECT 87.075 28.420 89.035 28.770 ;
        RECT 89.365 28.420 91.325 28.770 ;
        RECT 93.115 28.420 95.075 28.770 ;
        RECT 95.405 28.420 97.365 28.770 ;
        RECT 99.155 28.420 101.115 28.770 ;
        RECT 101.445 28.420 103.405 28.770 ;
        RECT 105.195 28.420 107.155 28.770 ;
        RECT 107.485 28.420 109.445 28.770 ;
        RECT 111.235 28.420 113.195 28.770 ;
        RECT 113.525 28.420 115.485 28.770 ;
        RECT 117.275 28.420 119.235 28.770 ;
        RECT 119.565 28.420 121.525 28.770 ;
        RECT 123.315 28.420 125.275 28.650 ;
        RECT 125.605 28.420 127.565 28.650 ;
        RECT 80.755 20.260 80.985 28.260 ;
        RECT 83.045 20.260 83.275 28.260 ;
        RECT 85.335 20.260 85.565 28.260 ;
        RECT 86.795 23.065 87.025 28.260 ;
        RECT 89.085 24.565 89.315 28.260 ;
        RECT 88.850 23.865 89.550 24.565 ;
        RECT 86.560 22.365 87.260 23.065 ;
        RECT 86.795 20.260 87.025 22.365 ;
        RECT 89.085 20.260 89.315 23.865 ;
        RECT 91.375 23.065 91.605 28.260 ;
        RECT 91.140 22.365 91.840 23.065 ;
        RECT 91.375 20.260 91.605 22.365 ;
        RECT 92.835 21.565 93.065 28.260 ;
        RECT 92.600 20.865 93.300 21.565 ;
        RECT 92.835 20.260 93.065 20.865 ;
        RECT 95.125 20.100 95.355 28.260 ;
        RECT 97.415 21.565 97.645 28.260 ;
        RECT 98.875 27.565 99.105 28.260 ;
        RECT 98.640 26.865 99.340 27.565 ;
        RECT 97.180 20.865 97.880 21.565 ;
        RECT 97.415 20.260 97.645 20.865 ;
        RECT 98.875 20.260 99.105 26.865 ;
        RECT 101.165 26.065 101.395 28.260 ;
        RECT 103.455 27.565 103.685 28.260 ;
        RECT 104.915 27.565 105.145 28.260 ;
        RECT 103.220 26.865 103.920 27.565 ;
        RECT 104.680 26.865 105.380 27.565 ;
        RECT 100.930 25.365 101.630 26.065 ;
        RECT 101.165 20.260 101.395 25.365 ;
        RECT 103.455 20.260 103.685 26.865 ;
        RECT 104.915 20.260 105.145 26.865 ;
        RECT 107.205 26.065 107.435 28.260 ;
        RECT 109.495 27.565 109.725 28.260 ;
        RECT 109.260 26.865 109.960 27.565 ;
        RECT 106.970 25.365 107.670 26.065 ;
        RECT 107.205 20.260 107.435 25.365 ;
        RECT 109.495 20.260 109.725 26.865 ;
        RECT 110.955 21.565 111.185 28.260 ;
        RECT 110.720 20.865 111.420 21.565 ;
        RECT 110.955 20.260 111.185 20.865 ;
        RECT 113.245 20.100 113.475 28.260 ;
        RECT 115.535 21.565 115.765 28.260 ;
        RECT 116.995 23.065 117.225 28.260 ;
        RECT 119.285 24.565 119.515 28.260 ;
        RECT 119.050 23.865 119.750 24.565 ;
        RECT 116.760 22.365 117.460 23.065 ;
        RECT 115.300 20.865 116.000 21.565 ;
        RECT 115.535 20.260 115.765 20.865 ;
        RECT 116.995 20.260 117.225 22.365 ;
        RECT 119.285 20.260 119.515 23.865 ;
        RECT 121.575 23.065 121.805 28.260 ;
        RECT 121.340 22.365 122.040 23.065 ;
        RECT 121.575 20.260 121.805 22.365 ;
        RECT 123.035 20.260 123.265 28.260 ;
        RECT 125.325 20.260 125.555 28.260 ;
        RECT 127.615 20.260 127.845 28.260 ;
        RECT 81.035 19.870 82.995 20.100 ;
        RECT 83.325 19.870 85.285 20.100 ;
        RECT 87.075 19.750 89.035 20.100 ;
        RECT 89.365 19.750 91.325 20.100 ;
        RECT 93.115 19.750 97.365 20.100 ;
        RECT 99.155 19.750 101.115 20.100 ;
        RECT 101.445 19.750 103.405 20.100 ;
        RECT 105.195 19.750 107.155 20.100 ;
        RECT 107.485 19.750 109.445 20.100 ;
        RECT 111.235 19.750 115.485 20.100 ;
        RECT 117.275 19.750 119.235 20.100 ;
        RECT 119.565 19.750 121.525 20.100 ;
        RECT 123.315 19.870 125.275 20.100 ;
        RECT 125.605 19.870 127.565 20.100 ;
        RECT 81.035 18.490 82.995 18.720 ;
        RECT 83.325 18.490 85.285 18.720 ;
        RECT 87.075 18.490 89.035 18.720 ;
        RECT 89.365 18.490 91.325 18.720 ;
        RECT 93.115 18.490 95.075 18.720 ;
        RECT 95.405 18.490 97.365 18.720 ;
        RECT 99.155 18.490 101.115 18.720 ;
        RECT 101.445 18.490 103.405 18.720 ;
        RECT 105.195 18.490 107.155 18.720 ;
        RECT 107.485 18.490 109.445 18.720 ;
        RECT 111.235 18.490 113.195 18.720 ;
        RECT 113.525 18.490 115.485 18.720 ;
        RECT 117.275 18.490 119.235 18.720 ;
        RECT 119.565 18.490 121.525 18.720 ;
        RECT 123.315 18.490 125.275 18.720 ;
        RECT 125.605 18.490 127.565 18.720 ;
        RECT 80.755 10.330 80.985 18.330 ;
        RECT 83.045 10.330 83.275 18.330 ;
        RECT 85.335 10.330 85.565 18.330 ;
        RECT 86.795 10.330 87.025 18.330 ;
        RECT 89.085 10.330 89.315 18.330 ;
        RECT 91.375 10.330 91.605 18.330 ;
        RECT 92.835 10.330 93.065 18.330 ;
        RECT 95.125 10.330 95.355 18.330 ;
        RECT 97.415 10.330 97.645 18.330 ;
        RECT 98.875 10.330 99.105 18.330 ;
        RECT 101.165 10.330 101.395 18.330 ;
        RECT 103.455 10.330 103.685 18.330 ;
        RECT 104.915 10.330 105.145 18.330 ;
        RECT 107.205 10.330 107.435 18.330 ;
        RECT 109.495 10.330 109.725 18.330 ;
        RECT 110.955 10.330 111.185 18.330 ;
        RECT 113.245 10.330 113.475 18.330 ;
        RECT 115.535 10.330 115.765 18.330 ;
        RECT 116.995 10.330 117.225 18.330 ;
        RECT 119.285 10.330 119.515 18.330 ;
        RECT 121.575 10.330 121.805 18.330 ;
        RECT 123.035 10.330 123.265 18.330 ;
        RECT 125.325 10.330 125.555 18.330 ;
        RECT 127.615 10.330 127.845 18.330 ;
        RECT 81.035 9.940 82.995 10.170 ;
        RECT 83.325 9.940 85.285 10.170 ;
        RECT 87.075 9.940 89.035 10.170 ;
        RECT 89.365 9.940 91.325 10.170 ;
        RECT 93.115 9.940 95.075 10.170 ;
        RECT 95.405 9.940 97.365 10.170 ;
        RECT 99.155 9.940 101.115 10.170 ;
        RECT 101.445 9.940 103.405 10.170 ;
        RECT 105.195 9.940 107.155 10.170 ;
        RECT 107.485 9.940 109.445 10.170 ;
        RECT 111.235 9.940 113.195 10.170 ;
        RECT 113.525 9.940 115.485 10.170 ;
        RECT 117.275 9.940 119.235 10.170 ;
        RECT 119.565 9.940 121.525 10.170 ;
        RECT 123.315 9.940 125.275 10.170 ;
        RECT 125.605 9.940 127.565 10.170 ;
        RECT 128.345 9.480 130.565 39.040 ;
        RECT 8.665 8.890 130.565 9.480 ;
        RECT 7.065 5.690 130.565 8.890 ;
        RECT 135.120 18.845 135.710 41.635 ;
        RECT 136.295 40.485 138.400 41.075 ;
        RECT 136.295 39.315 138.400 39.905 ;
        RECT 146.290 39.315 148.395 41.075 ;
        RECT 136.295 36.975 138.400 38.735 ;
        RECT 146.290 38.145 148.395 38.735 ;
        RECT 146.290 36.975 148.395 37.565 ;
        RECT 136.295 35.805 138.400 36.395 ;
        RECT 136.295 34.635 138.400 35.225 ;
        RECT 146.290 34.635 148.395 36.395 ;
        RECT 136.295 32.295 138.400 34.055 ;
        RECT 146.290 33.465 148.395 34.055 ;
        RECT 143.640 32.295 148.395 32.885 ;
        RECT 136.295 31.125 138.400 31.715 ;
        RECT 136.295 29.955 141.055 30.545 ;
        RECT 146.290 29.955 148.395 31.715 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 136.295 26.445 138.400 28.205 ;
        RECT 146.290 27.615 148.395 29.375 ;
        RECT 136.295 24.105 138.400 25.865 ;
        RECT 146.290 25.275 148.395 27.035 ;
        RECT 136.295 21.765 138.400 23.525 ;
        RECT 146.290 22.935 148.395 24.695 ;
        RECT 136.295 19.425 138.400 21.185 ;
        RECT 146.290 20.595 148.395 22.355 ;
        RECT 141.295 19.425 148.395 20.015 ;
        RECT 148.980 18.845 155.900 104.835 ;
        RECT 167.315 104.825 170.215 104.965 ;
        RECT 167.315 104.625 167.455 104.825 ;
        RECT 173.205 104.765 173.525 105.025 ;
        RECT 174.215 105.010 174.355 105.165 ;
        RECT 174.140 104.780 174.430 105.010 ;
        RECT 175.505 104.765 175.825 105.025 ;
        RECT 167.700 104.625 167.990 104.670 ;
        RECT 175.595 104.625 175.735 104.765 ;
        RECT 167.315 104.485 167.990 104.625 ;
        RECT 167.700 104.440 167.990 104.485 ;
        RECT 169.155 104.485 175.735 104.625 ;
        RECT 176.975 104.625 177.115 105.165 ;
        RECT 177.360 105.165 182.175 105.305 ;
        RECT 177.360 105.120 177.650 105.165 ;
        RECT 180.580 105.120 180.870 105.165 ;
        RECT 177.805 104.765 178.125 105.025 ;
        RECT 178.280 104.780 178.570 105.010 ;
        RECT 178.355 104.625 178.495 104.780 ;
        RECT 179.645 104.625 179.965 104.685 ;
        RECT 176.975 104.485 179.965 104.625 ;
        RECT 165.860 104.285 166.150 104.330 ;
        RECT 169.155 104.285 169.295 104.485 ;
        RECT 179.645 104.425 179.965 104.485 ;
        RECT 165.860 104.145 169.295 104.285 ;
        RECT 165.860 104.100 166.150 104.145 ;
        RECT 169.525 104.085 169.845 104.345 ;
        RECT 169.985 104.285 170.305 104.345 ;
        RECT 170.920 104.285 171.210 104.330 ;
        RECT 169.985 104.145 171.210 104.285 ;
        RECT 169.985 104.085 170.305 104.145 ;
        RECT 170.920 104.100 171.210 104.145 ;
        RECT 175.505 104.085 175.825 104.345 ;
        RECT 175.965 104.285 176.285 104.345 ;
        RECT 182.035 104.285 182.175 105.165 ;
        RECT 182.420 105.120 182.710 105.350 ;
        RECT 184.245 105.105 184.565 105.365 ;
        RECT 185.165 105.305 185.485 105.365 ;
        RECT 186.100 105.305 186.390 105.350 ;
        RECT 185.165 105.165 186.390 105.305 ;
        RECT 185.165 105.105 185.485 105.165 ;
        RECT 186.100 105.120 186.390 105.165 ;
        RECT 187.555 104.965 187.695 105.505 ;
        RECT 191.605 105.445 191.925 105.505 ;
        RECT 208.625 105.445 208.945 105.705 ;
        RECT 209.175 105.645 209.315 105.845 ;
        RECT 212.320 105.845 215.295 105.985 ;
        RECT 212.320 105.800 212.610 105.845 ;
        RECT 215.155 105.645 215.295 105.845 ;
        RECT 215.985 105.785 216.305 106.045 ;
        RECT 218.300 105.985 218.590 106.030 ;
        RECT 223.805 105.985 224.125 106.045 ;
        RECT 218.300 105.845 224.125 105.985 ;
        RECT 218.300 105.800 218.590 105.845 ;
        RECT 223.805 105.785 224.125 105.845 ;
        RECT 225.200 105.985 225.490 106.030 ;
        RECT 228.405 105.985 228.725 106.045 ;
        RECT 225.200 105.845 228.725 105.985 ;
        RECT 225.200 105.800 225.490 105.845 ;
        RECT 228.405 105.785 228.725 105.845 ;
        RECT 230.705 105.985 231.025 106.045 ;
        RECT 231.640 105.985 231.930 106.030 ;
        RECT 230.705 105.845 231.930 105.985 ;
        RECT 230.705 105.785 231.025 105.845 ;
        RECT 231.640 105.800 231.930 105.845 ;
        RECT 233.005 105.985 233.325 106.045 ;
        RECT 233.940 105.985 234.230 106.030 ;
        RECT 233.005 105.845 234.230 105.985 ;
        RECT 233.005 105.785 233.325 105.845 ;
        RECT 233.940 105.800 234.230 105.845 ;
        RECT 235.305 105.985 235.625 106.045 ;
        RECT 236.240 105.985 236.530 106.030 ;
        RECT 235.305 105.845 236.530 105.985 ;
        RECT 235.305 105.785 235.625 105.845 ;
        RECT 236.240 105.800 236.530 105.845 ;
        RECT 237.605 105.985 237.925 106.045 ;
        RECT 238.080 105.985 238.370 106.030 ;
        RECT 237.605 105.845 238.370 105.985 ;
        RECT 237.605 105.785 237.925 105.845 ;
        RECT 238.080 105.800 238.370 105.845 ;
        RECT 242.220 105.985 242.510 106.030 ;
        RECT 242.665 105.985 242.985 106.045 ;
        RECT 242.220 105.845 242.985 105.985 ;
        RECT 242.220 105.800 242.510 105.845 ;
        RECT 219.205 105.645 219.525 105.705 ;
        RECT 209.175 105.505 213.915 105.645 ;
        RECT 215.155 105.505 219.525 105.645 ;
        RECT 190.700 105.305 190.990 105.350 ;
        RECT 190.700 105.165 193.215 105.305 ;
        RECT 190.700 105.120 190.990 105.165 ;
        RECT 183.415 104.825 187.695 104.965 ;
        RECT 192.080 104.965 192.370 105.010 ;
        RECT 192.525 104.965 192.845 105.025 ;
        RECT 192.080 104.825 192.845 104.965 ;
        RECT 193.075 104.965 193.215 105.165 ;
        RECT 193.445 105.105 193.765 105.365 ;
        RECT 194.825 105.305 195.145 105.365 ;
        RECT 195.300 105.305 195.590 105.350 ;
        RECT 194.825 105.165 195.590 105.305 ;
        RECT 194.825 105.105 195.145 105.165 ;
        RECT 195.300 105.120 195.590 105.165 ;
        RECT 195.745 105.305 196.065 105.365 ;
        RECT 197.140 105.305 197.430 105.350 ;
        RECT 195.745 105.165 197.430 105.305 ;
        RECT 195.745 105.105 196.065 105.165 ;
        RECT 197.140 105.120 197.430 105.165 ;
        RECT 198.965 105.105 199.285 105.365 ;
        RECT 202.660 105.305 202.950 105.350 ;
        RECT 204.485 105.305 204.805 105.365 ;
        RECT 202.660 105.165 204.805 105.305 ;
        RECT 202.660 105.120 202.950 105.165 ;
        RECT 204.485 105.105 204.805 105.165 ;
        RECT 205.880 105.305 206.170 105.350 ;
        RECT 207.705 105.305 208.025 105.365 ;
        RECT 205.880 105.165 208.025 105.305 ;
        RECT 205.880 105.120 206.170 105.165 ;
        RECT 207.705 105.105 208.025 105.165 ;
        RECT 208.180 105.305 208.470 105.350 ;
        RECT 211.845 105.305 212.165 105.365 ;
        RECT 208.180 105.165 212.165 105.305 ;
        RECT 208.180 105.120 208.470 105.165 ;
        RECT 211.845 105.105 212.165 105.165 ;
        RECT 213.240 105.120 213.530 105.350 ;
        RECT 200.345 104.965 200.665 105.025 ;
        RECT 205.405 104.965 205.725 105.025 ;
        RECT 193.075 104.825 200.665 104.965 ;
        RECT 183.415 104.670 183.555 104.825 ;
        RECT 192.080 104.780 192.370 104.825 ;
        RECT 192.525 104.765 192.845 104.825 ;
        RECT 200.345 104.765 200.665 104.825 ;
        RECT 201.815 104.825 205.725 104.965 ;
        RECT 183.340 104.440 183.630 104.670 ;
        RECT 185.180 104.625 185.470 104.670 ;
        RECT 193.905 104.625 194.225 104.685 ;
        RECT 185.180 104.485 194.225 104.625 ;
        RECT 185.180 104.440 185.470 104.485 ;
        RECT 193.905 104.425 194.225 104.485 ;
        RECT 196.220 104.625 196.510 104.670 ;
        RECT 200.805 104.625 201.125 104.685 ;
        RECT 196.220 104.485 201.125 104.625 ;
        RECT 196.220 104.440 196.510 104.485 ;
        RECT 200.805 104.425 201.125 104.485 ;
        RECT 186.545 104.285 186.865 104.345 ;
        RECT 175.965 104.145 186.865 104.285 ;
        RECT 175.965 104.085 176.285 104.145 ;
        RECT 186.545 104.085 186.865 104.145 ;
        RECT 187.005 104.085 187.325 104.345 ;
        RECT 188.860 104.285 189.150 104.330 ;
        RECT 189.305 104.285 189.625 104.345 ;
        RECT 188.860 104.145 189.625 104.285 ;
        RECT 188.860 104.100 189.150 104.145 ;
        RECT 189.305 104.085 189.625 104.145 ;
        RECT 191.145 104.285 191.465 104.345 ;
        RECT 193.445 104.285 193.765 104.345 ;
        RECT 191.145 104.145 193.765 104.285 ;
        RECT 191.145 104.085 191.465 104.145 ;
        RECT 193.445 104.085 193.765 104.145 ;
        RECT 198.060 104.285 198.350 104.330 ;
        RECT 201.815 104.285 201.955 104.825 ;
        RECT 205.405 104.765 205.725 104.825 ;
        RECT 209.560 104.965 209.850 105.010 ;
        RECT 209.560 104.825 212.995 104.965 ;
        RECT 209.560 104.780 209.850 104.825 ;
        RECT 203.580 104.625 203.870 104.670 ;
        RECT 212.305 104.625 212.625 104.685 ;
        RECT 203.580 104.485 212.625 104.625 ;
        RECT 203.580 104.440 203.870 104.485 ;
        RECT 212.305 104.425 212.625 104.485 ;
        RECT 198.060 104.145 201.955 104.285 ;
        RECT 198.060 104.100 198.350 104.145 ;
        RECT 204.945 104.085 205.265 104.345 ;
        RECT 205.865 104.285 206.185 104.345 ;
        RECT 206.340 104.285 206.630 104.330 ;
        RECT 205.865 104.145 206.630 104.285 ;
        RECT 212.855 104.285 212.995 104.825 ;
        RECT 213.315 104.625 213.455 105.120 ;
        RECT 213.775 104.965 213.915 105.505 ;
        RECT 219.205 105.445 219.525 105.505 ;
        RECT 221.060 105.645 221.350 105.690 ;
        RECT 227.040 105.645 227.330 105.690 ;
        RECT 242.295 105.645 242.435 105.800 ;
        RECT 242.665 105.785 242.985 105.845 ;
        RECT 251.405 105.985 251.725 106.045 ;
        RECT 263.380 105.985 263.670 106.030 ;
        RECT 251.405 105.845 263.670 105.985 ;
        RECT 251.405 105.785 251.725 105.845 ;
        RECT 263.380 105.800 263.670 105.845 ;
        RECT 266.140 105.800 266.430 106.030 ;
        RECT 246.805 105.645 247.125 105.705 ;
        RECT 253.705 105.645 254.025 105.705 ;
        RECT 266.215 105.645 266.355 105.800 ;
        RECT 273.485 105.785 273.805 106.045 ;
        RECT 275.785 105.785 276.105 106.045 ;
        RECT 279.020 105.800 279.310 106.030 ;
        RECT 221.060 105.505 227.330 105.645 ;
        RECT 221.060 105.460 221.350 105.505 ;
        RECT 227.040 105.460 227.330 105.505 ;
        RECT 232.175 105.505 242.435 105.645 ;
        RECT 242.755 105.505 245.655 105.645 ;
        RECT 216.905 105.105 217.225 105.365 ;
        RECT 217.365 105.105 217.685 105.365 ;
        RECT 221.520 105.305 221.810 105.350 ;
        RECT 226.120 105.305 226.410 105.350 ;
        RECT 228.865 105.305 229.185 105.365 ;
        RECT 232.175 105.305 232.315 105.505 ;
        RECT 217.915 105.165 225.875 105.305 ;
        RECT 217.915 104.965 218.055 105.165 ;
        RECT 221.520 105.120 221.810 105.165 ;
        RECT 213.775 104.825 218.055 104.965 ;
        RECT 221.045 104.965 221.365 105.025 ;
        RECT 221.980 104.965 222.270 105.010 ;
        RECT 221.045 104.825 222.270 104.965 ;
        RECT 225.735 104.965 225.875 105.165 ;
        RECT 226.120 105.165 229.185 105.305 ;
        RECT 226.120 105.120 226.410 105.165 ;
        RECT 228.865 105.105 229.185 105.165 ;
        RECT 229.415 105.165 232.315 105.305 ;
        RECT 229.415 104.965 229.555 105.165 ;
        RECT 232.560 105.120 232.850 105.350 ;
        RECT 234.385 105.305 234.705 105.365 ;
        RECT 234.860 105.305 235.150 105.350 ;
        RECT 234.385 105.165 235.150 105.305 ;
        RECT 225.735 104.825 229.555 104.965 ;
        RECT 221.045 104.765 221.365 104.825 ;
        RECT 221.980 104.780 222.270 104.825 ;
        RECT 229.785 104.765 230.105 105.025 ;
        RECT 232.635 104.965 232.775 105.120 ;
        RECT 234.385 105.105 234.705 105.165 ;
        RECT 234.860 105.120 235.150 105.165 ;
        RECT 235.305 105.305 235.625 105.365 ;
        RECT 237.160 105.305 237.450 105.350 ;
        RECT 235.305 105.165 237.450 105.305 ;
        RECT 235.305 105.105 235.625 105.165 ;
        RECT 237.160 105.120 237.450 105.165 ;
        RECT 238.985 105.105 239.305 105.365 ;
        RECT 242.755 105.350 242.895 105.505 ;
        RECT 242.680 105.120 242.970 105.350 ;
        RECT 244.965 105.105 245.285 105.365 ;
        RECT 245.515 105.305 245.655 105.505 ;
        RECT 246.805 105.505 253.475 105.645 ;
        RECT 246.805 105.445 247.125 105.505 ;
        RECT 248.200 105.305 248.490 105.350 ;
        RECT 245.515 105.165 248.490 105.305 ;
        RECT 253.335 105.305 253.475 105.505 ;
        RECT 253.705 105.505 266.355 105.645 ;
        RECT 267.505 105.645 267.825 105.705 ;
        RECT 279.095 105.645 279.235 105.800 ;
        RECT 282.685 105.785 283.005 106.045 ;
        RECT 283.145 105.985 283.465 106.045 ;
        RECT 288.220 105.985 288.510 106.030 ;
        RECT 283.145 105.845 288.510 105.985 ;
        RECT 283.145 105.785 283.465 105.845 ;
        RECT 288.220 105.800 288.510 105.845 ;
        RECT 291.900 105.800 292.190 106.030 ;
        RECT 297.405 105.985 297.725 106.045 ;
        RECT 308.920 105.985 309.210 106.030 ;
        RECT 297.405 105.845 309.210 105.985 ;
        RECT 267.505 105.505 279.235 105.645 ;
        RECT 281.305 105.645 281.625 105.705 ;
        RECT 291.975 105.645 292.115 105.800 ;
        RECT 297.405 105.785 297.725 105.845 ;
        RECT 308.920 105.800 309.210 105.845 ;
        RECT 281.305 105.505 292.115 105.645 ;
        RECT 298.320 105.645 298.970 105.690 ;
        RECT 299.245 105.645 299.565 105.705 ;
        RECT 301.920 105.645 302.210 105.690 ;
        RECT 309.825 105.645 310.145 105.705 ;
        RECT 298.320 105.505 302.210 105.645 ;
        RECT 253.705 105.445 254.025 105.505 ;
        RECT 267.505 105.445 267.825 105.505 ;
        RECT 281.305 105.445 281.625 105.505 ;
        RECT 298.320 105.460 298.970 105.505 ;
        RECT 299.245 105.445 299.565 105.505 ;
        RECT 301.620 105.460 302.210 105.505 ;
        RECT 305.775 105.505 310.145 105.645 ;
        RECT 253.335 105.165 257.155 105.305 ;
        RECT 248.200 105.120 248.490 105.165 ;
        RECT 238.525 104.965 238.845 105.025 ;
        RECT 232.635 104.825 238.845 104.965 ;
        RECT 238.525 104.765 238.845 104.825 ;
        RECT 243.600 104.965 243.890 105.010 ;
        RECT 249.565 104.965 249.885 105.025 ;
        RECT 243.600 104.825 249.885 104.965 ;
        RECT 243.600 104.780 243.890 104.825 ;
        RECT 249.565 104.765 249.885 104.825 ;
        RECT 250.945 104.765 251.265 105.025 ;
        RECT 255.085 104.965 255.405 105.025 ;
        RECT 256.480 104.965 256.770 105.010 ;
        RECT 255.085 104.825 256.770 104.965 ;
        RECT 257.015 104.965 257.155 105.165 ;
        RECT 257.385 105.105 257.705 105.365 ;
        RECT 260.605 105.105 260.925 105.365 ;
        RECT 262.460 105.305 262.750 105.350 ;
        RECT 263.365 105.305 263.685 105.365 ;
        RECT 262.460 105.165 263.685 105.305 ;
        RECT 262.460 105.120 262.750 105.165 ;
        RECT 263.365 105.105 263.685 105.165 ;
        RECT 264.300 105.305 264.590 105.350 ;
        RECT 264.745 105.305 265.065 105.365 ;
        RECT 264.300 105.165 265.065 105.305 ;
        RECT 264.300 105.120 264.590 105.165 ;
        RECT 264.745 105.105 265.065 105.165 ;
        RECT 267.060 105.120 267.350 105.350 ;
        RECT 268.900 105.305 269.190 105.350 ;
        RECT 267.595 105.165 269.190 105.305 ;
        RECT 257.015 104.825 261.755 104.965 ;
        RECT 255.085 104.765 255.405 104.825 ;
        RECT 256.480 104.780 256.770 104.825 ;
        RECT 228.865 104.625 229.185 104.685 ;
        RECT 244.965 104.625 245.285 104.685 ;
        RECT 261.615 104.670 261.755 104.825 ;
        RECT 259.700 104.625 259.990 104.670 ;
        RECT 213.315 104.485 241.055 104.625 ;
        RECT 228.865 104.425 229.185 104.485 ;
        RECT 215.065 104.285 215.385 104.345 ;
        RECT 212.855 104.145 215.385 104.285 ;
        RECT 205.865 104.085 206.185 104.145 ;
        RECT 206.340 104.100 206.630 104.145 ;
        RECT 215.065 104.085 215.385 104.145 ;
        RECT 219.220 104.285 219.510 104.330 ;
        RECT 219.665 104.285 219.985 104.345 ;
        RECT 219.220 104.145 219.985 104.285 ;
        RECT 219.220 104.100 219.510 104.145 ;
        RECT 219.665 104.085 219.985 104.145 ;
        RECT 234.385 104.285 234.705 104.345 ;
        RECT 237.145 104.285 237.465 104.345 ;
        RECT 234.385 104.145 237.465 104.285 ;
        RECT 234.385 104.085 234.705 104.145 ;
        RECT 237.145 104.085 237.465 104.145 ;
        RECT 238.065 104.285 238.385 104.345 ;
        RECT 240.380 104.285 240.670 104.330 ;
        RECT 238.065 104.145 240.670 104.285 ;
        RECT 240.915 104.285 241.055 104.485 ;
        RECT 244.965 104.485 259.990 104.625 ;
        RECT 244.965 104.425 245.285 104.485 ;
        RECT 259.700 104.440 259.990 104.485 ;
        RECT 261.540 104.440 261.830 104.670 ;
        RECT 267.135 104.625 267.275 105.120 ;
        RECT 267.595 105.025 267.735 105.165 ;
        RECT 268.900 105.120 269.190 105.165 ;
        RECT 269.805 105.305 270.125 105.365 ;
        RECT 274.420 105.305 274.710 105.350 ;
        RECT 269.805 105.165 274.710 105.305 ;
        RECT 269.805 105.105 270.125 105.165 ;
        RECT 274.420 105.120 274.710 105.165 ;
        RECT 274.880 105.120 275.170 105.350 ;
        RECT 279.465 105.305 279.785 105.365 ;
        RECT 279.940 105.305 280.230 105.350 ;
        RECT 279.465 105.165 280.230 105.305 ;
        RECT 267.505 104.765 267.825 105.025 ;
        RECT 267.965 104.965 268.285 105.025 ;
        RECT 269.360 104.965 269.650 105.010 ;
        RECT 274.955 104.965 275.095 105.120 ;
        RECT 279.465 105.105 279.785 105.165 ;
        RECT 279.940 105.120 280.230 105.165 ;
        RECT 281.765 105.105 282.085 105.365 ;
        RECT 283.620 105.305 283.910 105.350 ;
        RECT 284.985 105.305 285.305 105.365 ;
        RECT 283.620 105.165 285.305 105.305 ;
        RECT 283.620 105.120 283.910 105.165 ;
        RECT 284.985 105.105 285.305 105.165 ;
        RECT 285.460 105.305 285.750 105.350 ;
        RECT 286.825 105.305 287.145 105.365 ;
        RECT 285.460 105.165 287.145 105.305 ;
        RECT 285.460 105.120 285.750 105.165 ;
        RECT 286.825 105.105 287.145 105.165 ;
        RECT 287.300 105.120 287.590 105.350 ;
        RECT 267.965 104.825 275.095 104.965 ;
        RECT 276.705 104.965 277.025 105.025 ;
        RECT 276.705 104.825 286.595 104.965 ;
        RECT 267.965 104.765 268.285 104.825 ;
        RECT 269.360 104.780 269.650 104.825 ;
        RECT 276.705 104.765 277.025 104.825 ;
        RECT 270.265 104.625 270.585 104.685 ;
        RECT 286.455 104.670 286.595 104.825 ;
        RECT 280.860 104.625 281.150 104.670 ;
        RECT 284.540 104.625 284.830 104.670 ;
        RECT 267.135 104.485 269.805 104.625 ;
        RECT 247.265 104.285 247.585 104.345 ;
        RECT 240.915 104.145 247.585 104.285 ;
        RECT 238.065 104.085 238.385 104.145 ;
        RECT 240.380 104.100 240.670 104.145 ;
        RECT 247.265 104.085 247.585 104.145 ;
        RECT 247.725 104.085 248.045 104.345 ;
        RECT 253.720 104.285 254.010 104.330 ;
        RECT 254.625 104.285 254.945 104.345 ;
        RECT 253.720 104.145 254.945 104.285 ;
        RECT 253.720 104.100 254.010 104.145 ;
        RECT 254.625 104.085 254.945 104.145 ;
        RECT 255.545 104.285 255.865 104.345 ;
        RECT 258.320 104.285 258.610 104.330 ;
        RECT 255.545 104.145 258.610 104.285 ;
        RECT 255.545 104.085 255.865 104.145 ;
        RECT 258.320 104.100 258.610 104.145 ;
        RECT 260.145 104.285 260.465 104.345 ;
        RECT 267.980 104.285 268.270 104.330 ;
        RECT 260.145 104.145 268.270 104.285 ;
        RECT 269.665 104.285 269.805 104.485 ;
        RECT 270.265 104.485 281.150 104.625 ;
        RECT 270.265 104.425 270.585 104.485 ;
        RECT 280.860 104.440 281.150 104.485 ;
        RECT 281.395 104.485 284.830 104.625 ;
        RECT 270.725 104.285 271.045 104.345 ;
        RECT 269.665 104.145 271.045 104.285 ;
        RECT 260.145 104.085 260.465 104.145 ;
        RECT 267.980 104.100 268.270 104.145 ;
        RECT 270.725 104.085 271.045 104.145 ;
        RECT 272.580 104.285 272.870 104.330 ;
        RECT 273.025 104.285 273.345 104.345 ;
        RECT 272.580 104.145 273.345 104.285 ;
        RECT 272.580 104.100 272.870 104.145 ;
        RECT 273.025 104.085 273.345 104.145 ;
        RECT 274.405 104.285 274.725 104.345 ;
        RECT 281.395 104.285 281.535 104.485 ;
        RECT 284.540 104.440 284.830 104.485 ;
        RECT 286.380 104.440 286.670 104.670 ;
        RECT 287.375 104.625 287.515 105.120 ;
        RECT 289.125 105.105 289.445 105.365 ;
        RECT 292.345 105.305 292.665 105.365 ;
        RECT 292.820 105.305 293.110 105.350 ;
        RECT 294.185 105.305 294.505 105.365 ;
        RECT 292.345 105.165 294.505 105.305 ;
        RECT 292.345 105.105 292.665 105.165 ;
        RECT 292.820 105.120 293.110 105.165 ;
        RECT 294.185 105.105 294.505 105.165 ;
        RECT 295.125 105.305 295.415 105.350 ;
        RECT 296.960 105.305 297.250 105.350 ;
        RECT 300.540 105.305 300.830 105.350 ;
        RECT 295.125 105.165 300.830 105.305 ;
        RECT 295.125 105.120 295.415 105.165 ;
        RECT 296.960 105.120 297.250 105.165 ;
        RECT 300.540 105.120 300.830 105.165 ;
        RECT 301.620 105.145 301.910 105.460 ;
        RECT 304.320 105.305 304.610 105.350 ;
        RECT 305.775 105.305 305.915 105.505 ;
        RECT 309.825 105.445 310.145 105.505 ;
        RECT 304.320 105.165 305.915 105.305 ;
        RECT 304.320 105.120 304.610 105.165 ;
        RECT 306.160 105.120 306.450 105.350 ;
        RECT 288.665 104.965 288.985 105.025 ;
        RECT 294.660 104.965 294.950 105.010 ;
        RECT 288.665 104.825 294.950 104.965 ;
        RECT 288.665 104.765 288.985 104.825 ;
        RECT 294.660 104.780 294.950 104.825 ;
        RECT 296.025 104.765 296.345 105.025 ;
        RECT 303.845 104.965 304.165 105.025 ;
        RECT 306.235 104.965 306.375 105.120 ;
        RECT 307.985 105.105 308.305 105.365 ;
        RECT 303.845 104.825 306.375 104.965 ;
        RECT 303.845 104.765 304.165 104.825 ;
        RECT 291.885 104.625 292.205 104.685 ;
        RECT 287.375 104.485 292.205 104.625 ;
        RECT 291.885 104.425 292.205 104.485 ;
        RECT 295.530 104.625 295.820 104.670 ;
        RECT 297.420 104.625 297.710 104.670 ;
        RECT 300.540 104.625 300.830 104.670 ;
        RECT 305.240 104.625 305.530 104.670 ;
        RECT 295.530 104.485 300.830 104.625 ;
        RECT 295.530 104.440 295.820 104.485 ;
        RECT 297.420 104.440 297.710 104.485 ;
        RECT 300.540 104.440 300.830 104.485 ;
        RECT 301.175 104.485 305.530 104.625 ;
        RECT 274.405 104.145 281.535 104.285 ;
        RECT 290.505 104.285 290.825 104.345 ;
        RECT 301.175 104.285 301.315 104.485 ;
        RECT 305.240 104.440 305.530 104.485 ;
        RECT 307.065 104.425 307.385 104.685 ;
        RECT 290.505 104.145 301.315 104.285 ;
        RECT 274.405 104.085 274.725 104.145 ;
        RECT 290.505 104.085 290.825 104.145 ;
        RECT 303.385 104.085 303.705 104.345 ;
        RECT 162.095 103.465 311.135 103.945 ;
        RECT 167.175 103.265 167.465 103.310 ;
        RECT 175.505 103.265 175.825 103.325 ;
        RECT 167.175 103.125 175.825 103.265 ;
        RECT 167.175 103.080 167.465 103.125 ;
        RECT 175.505 103.065 175.825 103.125 ;
        RECT 178.215 103.265 178.505 103.310 ;
        RECT 195.300 103.265 195.590 103.310 ;
        RECT 178.215 103.125 195.590 103.265 ;
        RECT 178.215 103.080 178.505 103.125 ;
        RECT 195.300 103.080 195.590 103.125 ;
        RECT 202.200 103.265 202.490 103.310 ;
        RECT 203.105 103.265 203.425 103.325 ;
        RECT 202.200 103.125 203.425 103.265 ;
        RECT 202.200 103.080 202.490 103.125 ;
        RECT 203.105 103.065 203.425 103.125 ;
        RECT 207.705 103.265 208.025 103.325 ;
        RECT 215.065 103.265 215.385 103.325 ;
        RECT 221.045 103.265 221.365 103.325 ;
        RECT 241.285 103.265 241.605 103.325 ;
        RECT 245.900 103.265 246.190 103.310 ;
        RECT 207.705 103.125 214.835 103.265 ;
        RECT 207.705 103.065 208.025 103.125 ;
        RECT 166.730 102.925 167.020 102.970 ;
        RECT 168.620 102.925 168.910 102.970 ;
        RECT 171.740 102.925 172.030 102.970 ;
        RECT 166.730 102.785 172.030 102.925 ;
        RECT 166.730 102.740 167.020 102.785 ;
        RECT 168.620 102.740 168.910 102.785 ;
        RECT 171.740 102.740 172.030 102.785 ;
        RECT 174.600 102.925 174.890 102.970 ;
        RECT 175.965 102.925 176.285 102.985 ;
        RECT 174.600 102.785 176.285 102.925 ;
        RECT 174.600 102.740 174.890 102.785 ;
        RECT 175.965 102.725 176.285 102.785 ;
        RECT 177.770 102.925 178.060 102.970 ;
        RECT 179.660 102.925 179.950 102.970 ;
        RECT 182.780 102.925 183.070 102.970 ;
        RECT 177.770 102.785 183.070 102.925 ;
        RECT 177.770 102.740 178.060 102.785 ;
        RECT 179.660 102.740 179.950 102.785 ;
        RECT 182.780 102.740 183.070 102.785 ;
        RECT 185.640 102.925 185.930 102.970 ;
        RECT 186.970 102.925 187.260 102.970 ;
        RECT 188.860 102.925 189.150 102.970 ;
        RECT 191.980 102.925 192.270 102.970 ;
        RECT 185.640 102.785 186.775 102.925 ;
        RECT 185.640 102.740 185.930 102.785 ;
        RECT 176.900 102.585 177.190 102.630 ;
        RECT 186.085 102.585 186.405 102.645 ;
        RECT 165.935 102.445 186.405 102.585 ;
        RECT 186.635 102.585 186.775 102.785 ;
        RECT 186.970 102.785 192.270 102.925 ;
        RECT 186.970 102.740 187.260 102.785 ;
        RECT 188.860 102.740 189.150 102.785 ;
        RECT 191.980 102.740 192.270 102.785 ;
        RECT 192.525 102.925 192.845 102.985 ;
        RECT 203.990 102.925 204.280 102.970 ;
        RECT 205.880 102.925 206.170 102.970 ;
        RECT 209.000 102.925 209.290 102.970 ;
        RECT 192.525 102.785 198.275 102.925 ;
        RECT 192.525 102.725 192.845 102.785 ;
        RECT 198.135 102.630 198.275 102.785 ;
        RECT 203.990 102.785 209.290 102.925 ;
        RECT 214.695 102.925 214.835 103.125 ;
        RECT 215.065 103.125 230.015 103.265 ;
        RECT 215.065 103.065 215.385 103.125 ;
        RECT 221.045 103.065 221.365 103.125 ;
        RECT 216.445 102.925 216.765 102.985 ;
        RECT 214.695 102.785 216.765 102.925 ;
        RECT 203.990 102.740 204.280 102.785 ;
        RECT 205.880 102.740 206.170 102.785 ;
        RECT 209.000 102.740 209.290 102.785 ;
        RECT 216.445 102.725 216.765 102.785 ;
        RECT 218.250 102.925 218.540 102.970 ;
        RECT 220.140 102.925 220.430 102.970 ;
        RECT 223.260 102.925 223.550 102.970 ;
        RECT 218.250 102.785 223.550 102.925 ;
        RECT 218.250 102.740 218.540 102.785 ;
        RECT 220.140 102.740 220.430 102.785 ;
        RECT 223.260 102.740 223.550 102.785 ;
        RECT 227.040 102.740 227.330 102.970 ;
        RECT 186.635 102.445 197.355 102.585 ;
        RECT 165.385 102.045 165.705 102.305 ;
        RECT 165.935 102.290 166.075 102.445 ;
        RECT 176.900 102.400 177.190 102.445 ;
        RECT 186.085 102.385 186.405 102.445 ;
        RECT 165.860 102.060 166.150 102.290 ;
        RECT 166.325 102.245 166.615 102.290 ;
        RECT 168.160 102.245 168.450 102.290 ;
        RECT 171.740 102.245 172.030 102.290 ;
        RECT 166.325 102.105 172.030 102.245 ;
        RECT 166.325 102.060 166.615 102.105 ;
        RECT 168.160 102.060 168.450 102.105 ;
        RECT 171.740 102.060 172.030 102.105 ;
        RECT 165.935 101.905 166.075 102.060 ;
        RECT 166.765 101.905 167.085 101.965 ;
        RECT 172.820 101.950 173.110 102.265 ;
        RECT 177.365 102.245 177.655 102.290 ;
        RECT 179.200 102.245 179.490 102.290 ;
        RECT 182.780 102.245 183.070 102.290 ;
        RECT 177.365 102.105 183.070 102.245 ;
        RECT 177.365 102.060 177.655 102.105 ;
        RECT 179.200 102.060 179.490 102.105 ;
        RECT 182.780 102.060 183.070 102.105 ;
        RECT 165.935 101.765 167.085 101.905 ;
        RECT 166.765 101.705 167.085 101.765 ;
        RECT 169.520 101.905 170.170 101.950 ;
        RECT 172.820 101.905 173.410 101.950 ;
        RECT 174.125 101.905 174.445 101.965 ;
        RECT 183.860 101.950 184.150 102.265 ;
        RECT 186.565 102.245 186.855 102.290 ;
        RECT 188.400 102.245 188.690 102.290 ;
        RECT 191.980 102.245 192.270 102.290 ;
        RECT 186.565 102.105 192.270 102.245 ;
        RECT 186.565 102.060 186.855 102.105 ;
        RECT 188.400 102.060 188.690 102.105 ;
        RECT 191.980 102.060 192.270 102.105 ;
        RECT 193.060 102.245 193.350 102.265 ;
        RECT 196.205 102.245 196.525 102.305 ;
        RECT 197.215 102.290 197.355 102.445 ;
        RECT 198.060 102.400 198.350 102.630 ;
        RECT 203.120 102.585 203.410 102.630 ;
        RECT 210.465 102.585 210.785 102.645 ;
        RECT 203.120 102.445 210.785 102.585 ;
        RECT 203.120 102.400 203.410 102.445 ;
        RECT 210.465 102.385 210.785 102.445 ;
        RECT 210.925 102.585 211.245 102.645 ;
        RECT 214.145 102.585 214.465 102.645 ;
        RECT 214.620 102.585 214.910 102.630 ;
        RECT 210.925 102.445 214.910 102.585 ;
        RECT 210.925 102.385 211.245 102.445 ;
        RECT 214.145 102.385 214.465 102.445 ;
        RECT 214.620 102.400 214.910 102.445 ;
        RECT 215.065 102.385 215.385 102.645 ;
        RECT 218.760 102.585 219.050 102.630 ;
        RECT 227.115 102.585 227.255 102.740 ;
        RECT 229.875 102.630 230.015 103.125 ;
        RECT 241.285 103.125 246.190 103.265 ;
        RECT 241.285 103.065 241.605 103.125 ;
        RECT 245.900 103.080 246.190 103.125 ;
        RECT 246.345 103.265 246.665 103.325 ;
        RECT 250.945 103.265 251.265 103.325 ;
        RECT 246.345 103.125 251.265 103.265 ;
        RECT 246.345 103.065 246.665 103.125 ;
        RECT 250.945 103.065 251.265 103.125 ;
        RECT 255.085 103.265 255.405 103.325 ;
        RECT 260.605 103.265 260.925 103.325 ;
        RECT 261.540 103.265 261.830 103.310 ;
        RECT 255.085 103.125 261.830 103.265 ;
        RECT 255.085 103.065 255.405 103.125 ;
        RECT 260.605 103.065 260.925 103.125 ;
        RECT 261.540 103.080 261.830 103.125 ;
        RECT 265.205 103.265 265.525 103.325 ;
        RECT 275.800 103.265 276.090 103.310 ;
        RECT 284.985 103.265 285.305 103.325 ;
        RECT 265.205 103.125 276.090 103.265 ;
        RECT 265.205 103.065 265.525 103.125 ;
        RECT 275.800 103.080 276.090 103.125 ;
        RECT 278.635 103.125 285.305 103.265 ;
        RECT 231.640 102.740 231.930 102.970 ;
        RECT 237.570 102.925 237.860 102.970 ;
        RECT 239.460 102.925 239.750 102.970 ;
        RECT 242.580 102.925 242.870 102.970 ;
        RECT 250.500 102.925 250.790 102.970 ;
        RECT 237.570 102.785 242.870 102.925 ;
        RECT 237.570 102.740 237.860 102.785 ;
        RECT 239.460 102.740 239.750 102.785 ;
        RECT 242.580 102.740 242.870 102.785 ;
        RECT 245.515 102.785 250.790 102.925 ;
        RECT 218.760 102.445 227.255 102.585 ;
        RECT 218.760 102.400 219.050 102.445 ;
        RECT 229.800 102.400 230.090 102.630 ;
        RECT 193.060 102.105 196.525 102.245 ;
        RECT 169.520 101.765 174.445 101.905 ;
        RECT 169.520 101.720 170.170 101.765 ;
        RECT 173.120 101.720 173.410 101.765 ;
        RECT 174.125 101.705 174.445 101.765 ;
        RECT 180.560 101.905 181.210 101.950 ;
        RECT 183.860 101.905 184.450 101.950 ;
        RECT 180.560 101.765 184.935 101.905 ;
        RECT 180.560 101.720 181.210 101.765 ;
        RECT 184.160 101.720 184.450 101.765 ;
        RECT 164.480 101.565 164.770 101.610 ;
        RECT 168.605 101.565 168.925 101.625 ;
        RECT 164.480 101.425 168.925 101.565 ;
        RECT 184.795 101.565 184.935 101.765 ;
        RECT 187.465 101.705 187.785 101.965 ;
        RECT 193.060 101.950 193.350 102.105 ;
        RECT 196.205 102.045 196.525 102.105 ;
        RECT 197.140 102.245 197.430 102.290 ;
        RECT 198.965 102.245 199.285 102.305 ;
        RECT 197.140 102.105 199.285 102.245 ;
        RECT 197.140 102.060 197.430 102.105 ;
        RECT 198.965 102.045 199.285 102.105 ;
        RECT 200.345 102.245 200.665 102.305 ;
        RECT 201.280 102.245 201.570 102.290 ;
        RECT 200.345 102.105 201.570 102.245 ;
        RECT 200.345 102.045 200.665 102.105 ;
        RECT 201.280 102.060 201.570 102.105 ;
        RECT 203.585 102.245 203.875 102.290 ;
        RECT 205.420 102.245 205.710 102.290 ;
        RECT 209.000 102.245 209.290 102.290 ;
        RECT 203.585 102.105 209.290 102.245 ;
        RECT 203.585 102.060 203.875 102.105 ;
        RECT 205.420 102.060 205.710 102.105 ;
        RECT 209.000 102.060 209.290 102.105 ;
        RECT 189.760 101.905 190.410 101.950 ;
        RECT 193.060 101.905 193.650 101.950 ;
        RECT 189.760 101.765 193.650 101.905 ;
        RECT 189.760 101.720 190.410 101.765 ;
        RECT 193.360 101.720 193.650 101.765 ;
        RECT 193.995 101.765 197.355 101.905 ;
        RECT 188.845 101.565 189.165 101.625 ;
        RECT 193.995 101.565 194.135 101.765 ;
        RECT 197.215 101.625 197.355 101.765 ;
        RECT 197.585 101.705 197.905 101.965 ;
        RECT 184.795 101.425 194.135 101.565 ;
        RECT 194.840 101.565 195.130 101.610 ;
        RECT 195.285 101.565 195.605 101.625 ;
        RECT 194.840 101.425 195.605 101.565 ;
        RECT 164.480 101.380 164.770 101.425 ;
        RECT 168.605 101.365 168.925 101.425 ;
        RECT 188.845 101.365 189.165 101.425 ;
        RECT 194.840 101.380 195.130 101.425 ;
        RECT 195.285 101.365 195.605 101.425 ;
        RECT 197.125 101.365 197.445 101.625 ;
        RECT 199.055 101.565 199.195 102.045 ;
        RECT 204.500 101.905 204.790 101.950 ;
        RECT 205.865 101.905 206.185 101.965 ;
        RECT 204.500 101.765 206.185 101.905 ;
        RECT 204.500 101.720 204.790 101.765 ;
        RECT 205.865 101.705 206.185 101.765 ;
        RECT 206.780 101.905 207.430 101.950 ;
        RECT 207.705 101.905 208.025 101.965 ;
        RECT 210.080 101.950 210.370 102.265 ;
        RECT 210.555 102.245 210.695 102.385 ;
        RECT 217.380 102.245 217.670 102.290 ;
        RECT 210.555 102.105 217.670 102.245 ;
        RECT 217.380 102.060 217.670 102.105 ;
        RECT 217.845 102.245 218.135 102.290 ;
        RECT 219.680 102.245 219.970 102.290 ;
        RECT 223.260 102.245 223.550 102.290 ;
        RECT 217.845 102.105 223.550 102.245 ;
        RECT 217.845 102.060 218.135 102.105 ;
        RECT 219.680 102.060 219.970 102.105 ;
        RECT 223.260 102.060 223.550 102.105 ;
        RECT 210.080 101.905 210.670 101.950 ;
        RECT 221.040 101.905 221.690 101.950 ;
        RECT 223.805 101.905 224.125 101.965 ;
        RECT 224.340 101.950 224.630 102.265 ;
        RECT 226.105 102.245 226.425 102.305 ;
        RECT 231.715 102.245 231.855 102.740 ;
        RECT 238.065 102.385 238.385 102.645 ;
        RECT 239.905 102.585 240.225 102.645 ;
        RECT 245.515 102.585 245.655 102.785 ;
        RECT 250.500 102.740 250.790 102.785 ;
        RECT 239.905 102.445 245.655 102.585 ;
        RECT 247.725 102.585 248.045 102.645 ;
        RECT 248.200 102.585 248.490 102.630 ;
        RECT 247.725 102.445 248.490 102.585 ;
        RECT 239.905 102.385 240.225 102.445 ;
        RECT 247.725 102.385 248.045 102.445 ;
        RECT 248.200 102.400 248.490 102.445 ;
        RECT 248.660 102.585 248.950 102.630 ;
        RECT 249.565 102.585 249.885 102.645 ;
        RECT 248.660 102.445 249.885 102.585 ;
        RECT 248.660 102.400 248.950 102.445 ;
        RECT 249.565 102.385 249.885 102.445 ;
        RECT 226.105 102.105 231.855 102.245 ;
        RECT 226.105 102.045 226.425 102.105 ;
        RECT 232.545 102.045 232.865 102.305 ;
        RECT 236.700 102.060 236.990 102.290 ;
        RECT 237.165 102.245 237.455 102.290 ;
        RECT 239.000 102.245 239.290 102.290 ;
        RECT 242.580 102.245 242.870 102.290 ;
        RECT 237.165 102.105 242.870 102.245 ;
        RECT 237.165 102.060 237.455 102.105 ;
        RECT 239.000 102.060 239.290 102.105 ;
        RECT 242.580 102.060 242.870 102.105 ;
        RECT 243.660 102.245 243.950 102.265 ;
        RECT 246.345 102.245 246.665 102.305 ;
        RECT 250.025 102.245 250.345 102.305 ;
        RECT 243.660 102.105 250.345 102.245 ;
        RECT 251.030 102.245 251.170 103.065 ;
        RECT 253.670 102.925 253.960 102.970 ;
        RECT 255.560 102.925 255.850 102.970 ;
        RECT 258.680 102.925 258.970 102.970 ;
        RECT 253.670 102.785 258.970 102.925 ;
        RECT 253.670 102.740 253.960 102.785 ;
        RECT 255.560 102.740 255.850 102.785 ;
        RECT 258.680 102.740 258.970 102.785 ;
        RECT 262.870 102.925 263.160 102.970 ;
        RECT 264.760 102.925 265.050 102.970 ;
        RECT 267.880 102.925 268.170 102.970 ;
        RECT 262.870 102.785 268.170 102.925 ;
        RECT 262.870 102.740 263.160 102.785 ;
        RECT 264.760 102.740 265.050 102.785 ;
        RECT 267.880 102.740 268.170 102.785 ;
        RECT 268.425 102.925 268.745 102.985 ;
        RECT 278.635 102.970 278.775 103.125 ;
        RECT 284.985 103.065 285.305 103.125 ;
        RECT 291.885 103.265 292.205 103.325 ;
        RECT 295.565 103.265 295.885 103.325 ;
        RECT 291.885 103.125 295.885 103.265 ;
        RECT 291.885 103.065 292.205 103.125 ;
        RECT 295.565 103.065 295.885 103.125 ;
        RECT 296.025 103.265 296.345 103.325 ;
        RECT 304.320 103.265 304.610 103.310 ;
        RECT 296.025 103.125 304.610 103.265 ;
        RECT 296.025 103.065 296.345 103.125 ;
        RECT 304.320 103.080 304.610 103.125 ;
        RECT 278.560 102.925 278.850 102.970 ;
        RECT 268.425 102.785 278.850 102.925 ;
        RECT 268.425 102.725 268.745 102.785 ;
        RECT 278.560 102.740 278.850 102.785 ;
        RECT 281.420 102.925 281.710 102.970 ;
        RECT 284.540 102.925 284.830 102.970 ;
        RECT 286.430 102.925 286.720 102.970 ;
        RECT 281.420 102.785 286.720 102.925 ;
        RECT 281.420 102.740 281.710 102.785 ;
        RECT 284.540 102.740 284.830 102.785 ;
        RECT 286.430 102.740 286.720 102.785 ;
        RECT 289.550 102.925 289.840 102.970 ;
        RECT 291.440 102.925 291.730 102.970 ;
        RECT 294.560 102.925 294.850 102.970 ;
        RECT 289.550 102.785 294.850 102.925 ;
        RECT 289.550 102.740 289.840 102.785 ;
        RECT 291.440 102.740 291.730 102.785 ;
        RECT 294.560 102.740 294.850 102.785 ;
        RECT 295.105 102.925 295.425 102.985 ;
        RECT 302.940 102.925 303.230 102.970 ;
        RECT 295.105 102.785 303.230 102.925 ;
        RECT 295.105 102.725 295.425 102.785 ;
        RECT 302.940 102.740 303.230 102.785 ;
        RECT 252.800 102.585 253.090 102.630 ;
        RECT 262.000 102.585 262.290 102.630 ;
        RECT 266.125 102.585 266.445 102.645 ;
        RECT 252.800 102.445 266.445 102.585 ;
        RECT 252.800 102.400 253.090 102.445 ;
        RECT 262.000 102.400 262.290 102.445 ;
        RECT 251.420 102.245 251.710 102.290 ;
        RECT 251.030 102.105 251.710 102.245 ;
        RECT 224.340 101.905 224.930 101.950 ;
        RECT 232.635 101.905 232.775 102.045 ;
        RECT 206.780 101.765 210.670 101.905 ;
        RECT 206.780 101.720 207.430 101.765 ;
        RECT 207.705 101.705 208.025 101.765 ;
        RECT 210.380 101.720 210.670 101.765 ;
        RECT 211.935 101.765 220.815 101.905 ;
        RECT 211.935 101.625 212.075 101.765 ;
        RECT 208.165 101.565 208.485 101.625 ;
        RECT 199.055 101.425 208.485 101.565 ;
        RECT 208.165 101.365 208.485 101.425 ;
        RECT 211.845 101.365 212.165 101.625 ;
        RECT 212.305 101.365 212.625 101.625 ;
        RECT 214.145 101.365 214.465 101.625 ;
        RECT 220.675 101.565 220.815 101.765 ;
        RECT 221.040 101.765 224.930 101.905 ;
        RECT 221.040 101.720 221.690 101.765 ;
        RECT 223.805 101.705 224.125 101.765 ;
        RECT 224.640 101.720 224.930 101.765 ;
        RECT 225.275 101.765 232.775 101.905 ;
        RECT 236.775 101.905 236.915 102.060 ;
        RECT 243.660 101.950 243.950 102.105 ;
        RECT 246.345 102.045 246.665 102.105 ;
        RECT 250.025 102.045 250.345 102.105 ;
        RECT 251.420 102.060 251.710 102.105 ;
        RECT 240.360 101.905 241.010 101.950 ;
        RECT 243.660 101.905 244.250 101.950 ;
        RECT 252.875 101.905 253.015 102.400 ;
        RECT 266.125 102.385 266.445 102.445 ;
        RECT 272.105 102.385 272.425 102.645 ;
        RECT 272.565 102.385 272.885 102.645 ;
        RECT 279.005 102.585 279.325 102.645 ;
        RECT 287.300 102.585 287.590 102.630 ;
        RECT 288.665 102.585 288.985 102.645 ;
        RECT 279.005 102.445 288.985 102.585 ;
        RECT 279.005 102.385 279.325 102.445 ;
        RECT 287.300 102.400 287.590 102.445 ;
        RECT 288.665 102.385 288.985 102.445 ;
        RECT 293.265 102.585 293.585 102.645 ;
        RECT 301.100 102.585 301.390 102.630 ;
        RECT 307.080 102.585 307.370 102.630 ;
        RECT 293.265 102.445 307.370 102.585 ;
        RECT 293.265 102.385 293.585 102.445 ;
        RECT 301.100 102.400 301.390 102.445 ;
        RECT 307.080 102.400 307.370 102.445 ;
        RECT 253.265 102.245 253.555 102.290 ;
        RECT 255.100 102.245 255.390 102.290 ;
        RECT 258.680 102.245 258.970 102.290 ;
        RECT 253.265 102.105 258.970 102.245 ;
        RECT 253.265 102.060 253.555 102.105 ;
        RECT 255.100 102.060 255.390 102.105 ;
        RECT 258.680 102.060 258.970 102.105 ;
        RECT 236.775 101.765 240.135 101.905 ;
        RECT 225.275 101.565 225.415 101.765 ;
        RECT 239.995 101.625 240.135 101.765 ;
        RECT 240.360 101.765 244.250 101.905 ;
        RECT 240.360 101.720 241.010 101.765 ;
        RECT 243.960 101.720 244.250 101.765 ;
        RECT 244.595 101.765 253.015 101.905 ;
        RECT 220.675 101.425 225.415 101.565 ;
        RECT 226.120 101.565 226.410 101.610 ;
        RECT 228.865 101.565 229.185 101.625 ;
        RECT 226.120 101.425 229.185 101.565 ;
        RECT 226.120 101.380 226.410 101.425 ;
        RECT 228.865 101.365 229.185 101.425 ;
        RECT 229.325 101.365 229.645 101.625 ;
        RECT 239.905 101.565 240.225 101.625 ;
        RECT 244.595 101.565 244.735 101.765 ;
        RECT 254.165 101.705 254.485 101.965 ;
        RECT 259.760 101.950 260.050 102.265 ;
        RECT 262.465 102.245 262.755 102.290 ;
        RECT 264.300 102.245 264.590 102.290 ;
        RECT 267.880 102.245 268.170 102.290 ;
        RECT 262.465 102.105 268.170 102.245 ;
        RECT 262.465 102.060 262.755 102.105 ;
        RECT 264.300 102.060 264.590 102.105 ;
        RECT 267.880 102.060 268.170 102.105 ;
        RECT 256.460 101.905 257.110 101.950 ;
        RECT 259.760 101.905 260.350 101.950 ;
        RECT 256.095 101.765 260.350 101.905 ;
        RECT 239.905 101.425 244.735 101.565 ;
        RECT 245.440 101.565 245.730 101.610 ;
        RECT 245.885 101.565 246.205 101.625 ;
        RECT 245.440 101.425 246.205 101.565 ;
        RECT 239.905 101.365 240.225 101.425 ;
        RECT 245.440 101.380 245.730 101.425 ;
        RECT 245.885 101.365 246.205 101.425 ;
        RECT 246.805 101.565 247.125 101.625 ;
        RECT 247.740 101.565 248.030 101.610 ;
        RECT 248.645 101.565 248.965 101.625 ;
        RECT 246.805 101.425 248.965 101.565 ;
        RECT 246.805 101.365 247.125 101.425 ;
        RECT 247.740 101.380 248.030 101.425 ;
        RECT 248.645 101.365 248.965 101.425 ;
        RECT 250.025 101.565 250.345 101.625 ;
        RECT 256.095 101.565 256.235 101.765 ;
        RECT 256.460 101.720 257.110 101.765 ;
        RECT 260.060 101.720 260.350 101.765 ;
        RECT 260.605 101.905 260.925 101.965 ;
        RECT 265.665 101.950 265.985 101.965 ;
        RECT 268.960 101.950 269.250 102.265 ;
        RECT 273.025 102.045 273.345 102.305 ;
        RECT 276.720 102.245 277.010 102.290 ;
        RECT 276.720 102.105 279.695 102.245 ;
        RECT 276.720 102.060 277.010 102.105 ;
        RECT 263.380 101.905 263.670 101.950 ;
        RECT 265.660 101.905 266.310 101.950 ;
        RECT 268.960 101.905 269.550 101.950 ;
        RECT 277.625 101.905 277.945 101.965 ;
        RECT 260.605 101.765 263.670 101.905 ;
        RECT 260.605 101.705 260.925 101.765 ;
        RECT 263.380 101.720 263.670 101.765 ;
        RECT 263.915 101.765 269.550 101.905 ;
        RECT 263.915 101.565 264.055 101.765 ;
        RECT 265.660 101.720 266.310 101.765 ;
        RECT 269.260 101.720 269.550 101.765 ;
        RECT 270.815 101.765 277.945 101.905 ;
        RECT 265.665 101.705 265.985 101.720 ;
        RECT 250.025 101.425 264.055 101.565 ;
        RECT 269.805 101.565 270.125 101.625 ;
        RECT 270.815 101.610 270.955 101.765 ;
        RECT 277.625 101.705 277.945 101.765 ;
        RECT 270.740 101.565 271.030 101.610 ;
        RECT 269.805 101.425 271.030 101.565 ;
        RECT 250.025 101.365 250.345 101.425 ;
        RECT 269.805 101.365 270.125 101.425 ;
        RECT 270.740 101.380 271.030 101.425 ;
        RECT 274.865 101.365 275.185 101.625 ;
        RECT 279.555 101.565 279.695 102.105 ;
        RECT 280.340 101.950 280.630 102.265 ;
        RECT 281.420 102.245 281.710 102.290 ;
        RECT 285.000 102.245 285.290 102.290 ;
        RECT 286.835 102.245 287.125 102.290 ;
        RECT 281.420 102.105 287.125 102.245 ;
        RECT 281.420 102.060 281.710 102.105 ;
        RECT 285.000 102.060 285.290 102.105 ;
        RECT 286.835 102.060 287.125 102.105 ;
        RECT 289.145 102.245 289.435 102.290 ;
        RECT 290.980 102.245 291.270 102.290 ;
        RECT 294.560 102.245 294.850 102.290 ;
        RECT 289.145 102.105 294.850 102.245 ;
        RECT 289.145 102.060 289.435 102.105 ;
        RECT 290.980 102.060 291.270 102.105 ;
        RECT 294.560 102.060 294.850 102.105 ;
        RECT 280.040 101.905 280.630 101.950 ;
        RECT 282.685 101.905 283.005 101.965 ;
        RECT 283.280 101.905 283.930 101.950 ;
        RECT 280.040 101.765 283.930 101.905 ;
        RECT 280.040 101.720 280.330 101.765 ;
        RECT 282.685 101.705 283.005 101.765 ;
        RECT 283.280 101.720 283.930 101.765 ;
        RECT 285.905 101.705 286.225 101.965 ;
        RECT 290.045 101.705 290.365 101.965 ;
        RECT 290.505 101.905 290.825 101.965 ;
        RECT 295.640 101.950 295.930 102.265 ;
        RECT 296.485 102.245 296.805 102.305 ;
        RECT 302.020 102.245 302.310 102.290 ;
        RECT 296.485 102.105 302.310 102.245 ;
        RECT 296.485 102.045 296.805 102.105 ;
        RECT 302.020 102.060 302.310 102.105 ;
        RECT 303.385 102.245 303.705 102.305 ;
        RECT 306.160 102.245 306.450 102.290 ;
        RECT 303.385 102.105 306.450 102.245 ;
        RECT 303.385 102.045 303.705 102.105 ;
        RECT 306.160 102.060 306.450 102.105 ;
        RECT 292.340 101.905 292.990 101.950 ;
        RECT 295.640 101.905 296.230 101.950 ;
        RECT 296.945 101.905 297.265 101.965 ;
        RECT 299.720 101.905 300.010 101.950 ;
        RECT 290.505 101.765 296.230 101.905 ;
        RECT 290.505 101.705 290.825 101.765 ;
        RECT 292.340 101.720 292.990 101.765 ;
        RECT 295.940 101.720 296.230 101.765 ;
        RECT 296.575 101.765 300.010 101.905 ;
        RECT 280.845 101.565 281.165 101.625 ;
        RECT 279.555 101.425 281.165 101.565 ;
        RECT 280.845 101.365 281.165 101.425 ;
        RECT 294.185 101.565 294.505 101.625 ;
        RECT 296.575 101.565 296.715 101.765 ;
        RECT 296.945 101.705 297.265 101.765 ;
        RECT 299.720 101.720 300.010 101.765 ;
        RECT 300.180 101.905 300.470 101.950 ;
        RECT 304.765 101.905 305.085 101.965 ;
        RECT 300.180 101.765 305.085 101.905 ;
        RECT 300.180 101.720 300.470 101.765 ;
        RECT 304.765 101.705 305.085 101.765 ;
        RECT 294.185 101.425 296.715 101.565 ;
        RECT 294.185 101.365 294.505 101.425 ;
        RECT 297.405 101.365 297.725 101.625 ;
        RECT 297.865 101.365 298.185 101.625 ;
        RECT 306.145 101.565 306.465 101.625 ;
        RECT 306.620 101.565 306.910 101.610 ;
        RECT 306.145 101.425 306.910 101.565 ;
        RECT 306.145 101.365 306.465 101.425 ;
        RECT 306.620 101.380 306.910 101.425 ;
        RECT 162.095 100.745 311.135 101.225 ;
        RECT 164.005 100.345 164.325 100.605 ;
        RECT 166.305 100.345 166.625 100.605 ;
        RECT 180.105 100.545 180.425 100.605 ;
        RECT 181.040 100.545 181.330 100.590 ;
        RECT 180.105 100.405 181.330 100.545 ;
        RECT 180.105 100.345 180.425 100.405 ;
        RECT 181.040 100.360 181.330 100.405 ;
        RECT 182.865 100.545 183.185 100.605 ;
        RECT 183.340 100.545 183.630 100.590 ;
        RECT 182.865 100.405 183.630 100.545 ;
        RECT 182.865 100.345 183.185 100.405 ;
        RECT 183.340 100.360 183.630 100.405 ;
        RECT 184.705 100.545 185.025 100.605 ;
        RECT 185.640 100.545 185.930 100.590 ;
        RECT 184.705 100.405 185.930 100.545 ;
        RECT 184.705 100.345 185.025 100.405 ;
        RECT 185.640 100.360 185.930 100.405 ;
        RECT 197.140 100.545 197.430 100.590 ;
        RECT 200.345 100.545 200.665 100.605 ;
        RECT 212.305 100.545 212.625 100.605 ;
        RECT 197.140 100.405 200.665 100.545 ;
        RECT 197.140 100.360 197.430 100.405 ;
        RECT 200.345 100.345 200.665 100.405 ;
        RECT 210.095 100.405 212.625 100.545 ;
        RECT 168.620 100.205 168.910 100.250 ;
        RECT 169.985 100.205 170.305 100.265 ;
        RECT 168.620 100.065 170.305 100.205 ;
        RECT 168.620 100.020 168.910 100.065 ;
        RECT 169.985 100.005 170.305 100.065 ;
        RECT 170.900 100.205 171.550 100.250 ;
        RECT 174.500 100.205 174.790 100.250 ;
        RECT 170.900 100.065 174.790 100.205 ;
        RECT 170.900 100.020 171.550 100.065 ;
        RECT 174.200 100.020 174.790 100.065 ;
        RECT 186.085 100.205 186.405 100.265 ;
        RECT 189.305 100.205 189.625 100.265 ;
        RECT 189.780 100.205 190.070 100.250 ;
        RECT 186.085 100.065 188.615 100.205 ;
        RECT 174.200 99.925 174.490 100.020 ;
        RECT 186.085 100.005 186.405 100.065 ;
        RECT 164.925 99.665 165.245 99.925 ;
        RECT 165.385 99.665 165.705 99.925 ;
        RECT 166.765 99.865 167.085 99.925 ;
        RECT 167.240 99.865 167.530 99.910 ;
        RECT 166.765 99.725 167.530 99.865 ;
        RECT 166.765 99.665 167.085 99.725 ;
        RECT 167.240 99.680 167.530 99.725 ;
        RECT 167.705 99.865 167.995 99.910 ;
        RECT 169.540 99.865 169.830 99.910 ;
        RECT 173.120 99.865 173.410 99.910 ;
        RECT 167.705 99.725 173.410 99.865 ;
        RECT 167.705 99.680 167.995 99.725 ;
        RECT 169.540 99.680 169.830 99.725 ;
        RECT 173.120 99.680 173.410 99.725 ;
        RECT 174.125 99.705 174.490 99.925 ;
        RECT 178.280 99.865 178.570 99.910 ;
        RECT 180.105 99.865 180.425 99.925 ;
        RECT 181.960 99.865 182.250 99.910 ;
        RECT 182.865 99.865 183.185 99.925 ;
        RECT 178.280 99.725 181.715 99.865 ;
        RECT 174.125 99.665 174.445 99.705 ;
        RECT 178.280 99.680 178.570 99.725 ;
        RECT 180.105 99.665 180.425 99.725 ;
        RECT 175.965 99.325 176.285 99.585 ;
        RECT 178.740 99.340 179.030 99.570 ;
        RECT 168.110 99.185 168.400 99.230 ;
        RECT 170.000 99.185 170.290 99.230 ;
        RECT 173.120 99.185 173.410 99.230 ;
        RECT 168.110 99.045 173.410 99.185 ;
        RECT 168.110 99.000 168.400 99.045 ;
        RECT 170.000 99.000 170.290 99.045 ;
        RECT 173.120 99.000 173.410 99.045 ;
        RECT 176.425 98.645 176.745 98.905 ;
        RECT 178.815 98.845 178.955 99.340 ;
        RECT 179.645 99.325 179.965 99.585 ;
        RECT 181.575 99.185 181.715 99.725 ;
        RECT 181.960 99.725 183.185 99.865 ;
        RECT 181.960 99.680 182.250 99.725 ;
        RECT 182.865 99.665 183.185 99.725 ;
        RECT 183.785 99.865 184.105 99.925 ;
        RECT 184.260 99.865 184.550 99.910 ;
        RECT 183.785 99.725 184.550 99.865 ;
        RECT 183.785 99.665 184.105 99.725 ;
        RECT 184.260 99.680 184.550 99.725 ;
        RECT 186.545 99.665 186.865 99.925 ;
        RECT 188.475 99.910 188.615 100.065 ;
        RECT 189.305 100.065 190.070 100.205 ;
        RECT 189.305 100.005 189.625 100.065 ;
        RECT 189.780 100.020 190.070 100.065 ;
        RECT 192.060 100.205 192.710 100.250 ;
        RECT 195.660 100.205 195.950 100.250 ;
        RECT 196.205 100.205 196.525 100.265 ;
        RECT 198.045 100.205 198.365 100.265 ;
        RECT 207.705 100.250 208.025 100.265 ;
        RECT 210.095 100.250 210.235 100.405 ;
        RECT 212.305 100.345 212.625 100.405 ;
        RECT 214.605 100.545 214.925 100.605 ;
        RECT 215.540 100.545 215.830 100.590 ;
        RECT 214.605 100.405 215.830 100.545 ;
        RECT 214.605 100.345 214.925 100.405 ;
        RECT 215.540 100.360 215.830 100.405 ;
        RECT 219.665 100.345 219.985 100.605 ;
        RECT 226.120 100.545 226.410 100.590 ;
        RECT 229.785 100.545 230.105 100.605 ;
        RECT 226.120 100.405 230.105 100.545 ;
        RECT 226.120 100.360 226.410 100.405 ;
        RECT 229.785 100.345 230.105 100.405 ;
        RECT 232.545 100.545 232.865 100.605 ;
        RECT 250.485 100.545 250.805 100.605 ;
        RECT 232.545 100.405 250.805 100.545 ;
        RECT 232.545 100.345 232.865 100.405 ;
        RECT 250.485 100.345 250.805 100.405 ;
        RECT 252.340 100.545 252.630 100.590 ;
        RECT 254.165 100.545 254.485 100.605 ;
        RECT 252.340 100.405 254.485 100.545 ;
        RECT 252.340 100.360 252.630 100.405 ;
        RECT 254.165 100.345 254.485 100.405 ;
        RECT 254.625 100.345 254.945 100.605 ;
        RECT 259.225 100.545 259.545 100.605 ;
        RECT 255.865 100.405 259.545 100.545 ;
        RECT 192.060 100.065 198.365 100.205 ;
        RECT 192.060 100.020 192.710 100.065 ;
        RECT 195.360 100.020 195.950 100.065 ;
        RECT 188.400 99.680 188.690 99.910 ;
        RECT 188.865 99.865 189.155 99.910 ;
        RECT 190.700 99.865 190.990 99.910 ;
        RECT 194.280 99.865 194.570 99.910 ;
        RECT 188.865 99.725 194.570 99.865 ;
        RECT 188.865 99.680 189.155 99.725 ;
        RECT 190.700 99.680 190.990 99.725 ;
        RECT 194.280 99.680 194.570 99.725 ;
        RECT 195.360 99.705 195.650 100.020 ;
        RECT 196.205 100.005 196.525 100.065 ;
        RECT 198.045 100.005 198.365 100.065 ;
        RECT 204.140 100.205 204.430 100.250 ;
        RECT 207.380 100.205 208.030 100.250 ;
        RECT 204.140 100.065 208.030 100.205 ;
        RECT 204.140 100.020 204.730 100.065 ;
        RECT 207.380 100.020 208.030 100.065 ;
        RECT 210.020 100.020 210.310 100.250 ;
        RECT 210.465 100.205 210.785 100.265 ;
        RECT 218.760 100.205 219.050 100.250 ;
        RECT 219.755 100.205 219.895 100.345 ;
        RECT 221.045 100.250 221.365 100.265 ;
        RECT 210.465 100.065 211.615 100.205 ;
        RECT 204.440 99.705 204.730 100.020 ;
        RECT 207.705 100.005 208.025 100.020 ;
        RECT 210.465 100.005 210.785 100.065 ;
        RECT 211.475 99.910 211.615 100.065 ;
        RECT 218.760 100.065 219.895 100.205 ;
        RECT 221.040 100.205 221.690 100.250 ;
        RECT 224.640 100.205 224.930 100.250 ;
        RECT 221.040 100.065 224.930 100.205 ;
        RECT 218.760 100.020 219.050 100.065 ;
        RECT 221.040 100.020 221.690 100.065 ;
        RECT 224.340 100.020 224.930 100.065 ;
        RECT 221.045 100.005 221.365 100.020 ;
        RECT 205.520 99.865 205.810 99.910 ;
        RECT 209.100 99.865 209.390 99.910 ;
        RECT 210.935 99.865 211.225 99.910 ;
        RECT 205.520 99.725 211.225 99.865 ;
        RECT 205.520 99.680 205.810 99.725 ;
        RECT 209.100 99.680 209.390 99.725 ;
        RECT 210.935 99.680 211.225 99.725 ;
        RECT 211.400 99.680 211.690 99.910 ;
        RECT 213.240 99.865 213.530 99.910 ;
        RECT 213.685 99.865 214.005 99.925 ;
        RECT 213.240 99.725 214.005 99.865 ;
        RECT 213.240 99.680 213.530 99.725 ;
        RECT 192.985 99.525 193.305 99.585 ;
        RECT 211.475 99.525 211.615 99.680 ;
        RECT 213.685 99.665 214.005 99.725 ;
        RECT 215.525 99.865 215.845 99.925 ;
        RECT 216.460 99.865 216.750 99.910 ;
        RECT 215.525 99.725 216.750 99.865 ;
        RECT 215.525 99.665 215.845 99.725 ;
        RECT 216.460 99.680 216.750 99.725 ;
        RECT 217.845 99.865 218.135 99.910 ;
        RECT 219.680 99.865 219.970 99.910 ;
        RECT 223.260 99.865 223.550 99.910 ;
        RECT 217.845 99.725 223.550 99.865 ;
        RECT 217.845 99.680 218.135 99.725 ;
        RECT 219.680 99.680 219.970 99.725 ;
        RECT 223.260 99.680 223.550 99.725 ;
        RECT 224.340 99.705 224.630 100.020 ;
        RECT 241.285 100.005 241.605 100.265 ;
        RECT 243.580 100.205 244.230 100.250 ;
        RECT 246.345 100.205 246.665 100.265 ;
        RECT 247.180 100.205 247.470 100.250 ;
        RECT 252.785 100.205 253.105 100.265 ;
        RECT 255.865 100.205 256.005 100.405 ;
        RECT 259.225 100.345 259.545 100.405 ;
        RECT 260.145 100.545 260.465 100.605 ;
        RECT 262.000 100.545 262.290 100.590 ;
        RECT 260.145 100.405 262.290 100.545 ;
        RECT 260.145 100.345 260.465 100.405 ;
        RECT 262.000 100.360 262.290 100.405 ;
        RECT 262.920 100.360 263.210 100.590 ;
        RECT 265.665 100.545 265.985 100.605 ;
        RECT 284.525 100.545 284.845 100.605 ;
        RECT 265.665 100.405 271.415 100.545 ;
        RECT 243.580 100.065 247.470 100.205 ;
        RECT 243.580 100.020 244.230 100.065 ;
        RECT 246.345 100.005 246.665 100.065 ;
        RECT 246.880 100.020 247.470 100.065 ;
        RECT 249.195 100.065 253.105 100.205 ;
        RECT 226.105 99.865 226.425 99.925 ;
        RECT 227.960 99.865 228.250 99.910 ;
        RECT 226.105 99.725 228.250 99.865 ;
        RECT 226.105 99.665 226.425 99.725 ;
        RECT 227.960 99.680 228.250 99.725 ;
        RECT 228.405 99.865 228.725 99.925 ;
        RECT 230.245 99.910 230.565 99.925 ;
        RECT 228.405 99.725 228.920 99.865 ;
        RECT 228.405 99.665 228.725 99.725 ;
        RECT 229.340 99.680 229.630 99.910 ;
        RECT 229.800 99.680 230.090 99.910 ;
        RECT 230.245 99.865 230.575 99.910 ;
        RECT 230.245 99.725 230.760 99.865 ;
        RECT 230.245 99.680 230.575 99.725 ;
        RECT 217.380 99.525 217.670 99.570 ;
        RECT 229.415 99.525 229.555 99.680 ;
        RECT 192.985 99.385 211.155 99.525 ;
        RECT 211.475 99.385 217.670 99.525 ;
        RECT 192.985 99.325 193.305 99.385 ;
        RECT 186.545 99.185 186.865 99.245 ;
        RECT 181.575 99.045 186.865 99.185 ;
        RECT 186.545 98.985 186.865 99.045 ;
        RECT 189.270 99.185 189.560 99.230 ;
        RECT 191.160 99.185 191.450 99.230 ;
        RECT 194.280 99.185 194.570 99.230 ;
        RECT 205.520 99.185 205.810 99.230 ;
        RECT 208.640 99.185 208.930 99.230 ;
        RECT 210.530 99.185 210.820 99.230 ;
        RECT 189.270 99.045 194.570 99.185 ;
        RECT 189.270 99.000 189.560 99.045 ;
        RECT 191.160 99.000 191.450 99.045 ;
        RECT 194.280 99.000 194.570 99.045 ;
        RECT 194.915 99.045 205.175 99.185 ;
        RECT 187.925 98.845 188.245 98.905 ;
        RECT 189.765 98.845 190.085 98.905 ;
        RECT 178.815 98.705 190.085 98.845 ;
        RECT 187.925 98.645 188.245 98.705 ;
        RECT 189.765 98.645 190.085 98.705 ;
        RECT 193.445 98.845 193.765 98.905 ;
        RECT 194.915 98.845 195.055 99.045 ;
        RECT 193.445 98.705 195.055 98.845 ;
        RECT 202.660 98.845 202.950 98.890 ;
        RECT 204.485 98.845 204.805 98.905 ;
        RECT 202.660 98.705 204.805 98.845 ;
        RECT 205.035 98.845 205.175 99.045 ;
        RECT 205.520 99.045 210.820 99.185 ;
        RECT 211.015 99.185 211.155 99.385 ;
        RECT 217.380 99.340 217.670 99.385 ;
        RECT 217.915 99.385 229.555 99.525 ;
        RECT 229.875 99.525 230.015 99.680 ;
        RECT 230.245 99.665 230.565 99.680 ;
        RECT 239.905 99.665 240.225 99.925 ;
        RECT 240.385 99.865 240.675 99.910 ;
        RECT 242.220 99.865 242.510 99.910 ;
        RECT 245.800 99.865 246.090 99.910 ;
        RECT 240.385 99.725 246.090 99.865 ;
        RECT 240.385 99.680 240.675 99.725 ;
        RECT 242.220 99.680 242.510 99.725 ;
        RECT 245.800 99.680 246.090 99.725 ;
        RECT 246.880 99.705 247.170 100.020 ;
        RECT 247.725 99.865 248.045 99.925 ;
        RECT 249.195 99.910 249.335 100.065 ;
        RECT 252.785 100.005 253.105 100.065 ;
        RECT 253.335 100.065 256.005 100.205 ;
        RECT 256.465 100.205 256.785 100.265 ;
        RECT 259.685 100.205 260.005 100.265 ;
        RECT 262.995 100.205 263.135 100.360 ;
        RECT 265.665 100.345 265.985 100.405 ;
        RECT 256.465 100.065 258.535 100.205 ;
        RECT 249.120 99.865 249.410 99.910 ;
        RECT 247.725 99.725 249.410 99.865 ;
        RECT 247.725 99.665 248.045 99.725 ;
        RECT 249.120 99.680 249.410 99.725 ;
        RECT 250.025 99.665 250.345 99.925 ;
        RECT 250.485 99.665 250.805 99.925 ;
        RECT 250.945 99.865 251.265 99.925 ;
        RECT 253.335 99.865 253.475 100.065 ;
        RECT 256.465 100.005 256.785 100.065 ;
        RECT 250.945 99.725 253.475 99.865 ;
        RECT 250.945 99.665 251.265 99.725 ;
        RECT 254.165 99.665 254.485 99.925 ;
        RECT 256.925 99.865 257.245 99.925 ;
        RECT 257.860 99.865 258.150 99.910 ;
        RECT 256.925 99.725 258.150 99.865 ;
        RECT 258.395 99.865 258.535 100.065 ;
        RECT 259.685 100.065 263.135 100.205 ;
        RECT 267.160 100.205 267.450 100.250 ;
        RECT 270.400 100.205 271.050 100.250 ;
        RECT 271.275 100.205 271.415 100.405 ;
        RECT 272.655 100.405 284.845 100.545 ;
        RECT 272.655 100.205 272.795 100.405 ;
        RECT 284.525 100.345 284.845 100.405 ;
        RECT 285.905 100.545 286.225 100.605 ;
        RECT 287.760 100.545 288.050 100.590 ;
        RECT 285.905 100.405 288.050 100.545 ;
        RECT 285.905 100.345 286.225 100.405 ;
        RECT 287.760 100.360 288.050 100.405 ;
        RECT 288.205 100.545 288.525 100.605 ;
        RECT 292.360 100.545 292.650 100.590 ;
        RECT 298.325 100.545 298.645 100.605 ;
        RECT 288.205 100.405 292.650 100.545 ;
        RECT 288.205 100.345 288.525 100.405 ;
        RECT 292.360 100.360 292.650 100.405 ;
        RECT 292.895 100.405 298.645 100.545 ;
        RECT 267.160 100.065 272.795 100.205 ;
        RECT 273.040 100.205 273.330 100.250 ;
        RECT 274.865 100.205 275.185 100.265 ;
        RECT 273.040 100.065 275.185 100.205 ;
        RECT 259.685 100.005 260.005 100.065 ;
        RECT 267.160 100.020 267.750 100.065 ;
        RECT 270.400 100.020 271.050 100.065 ;
        RECT 273.040 100.020 273.330 100.065 ;
        RECT 260.160 99.865 260.450 99.910 ;
        RECT 260.605 99.865 260.925 99.925 ;
        RECT 258.395 99.725 259.915 99.865 ;
        RECT 256.925 99.665 257.245 99.725 ;
        RECT 257.860 99.680 258.150 99.725 ;
        RECT 259.775 99.585 259.915 99.725 ;
        RECT 260.160 99.725 260.925 99.865 ;
        RECT 260.160 99.680 260.450 99.725 ;
        RECT 260.605 99.665 260.925 99.725 ;
        RECT 263.840 99.865 264.130 99.910 ;
        RECT 264.285 99.865 264.605 99.925 ;
        RECT 263.840 99.725 264.605 99.865 ;
        RECT 263.840 99.680 264.130 99.725 ;
        RECT 264.285 99.665 264.605 99.725 ;
        RECT 267.460 99.705 267.750 100.020 ;
        RECT 274.865 100.005 275.185 100.065 ;
        RECT 278.540 100.205 279.190 100.250 ;
        RECT 282.140 100.205 282.430 100.250 ;
        RECT 282.685 100.205 283.005 100.265 ;
        RECT 290.505 100.205 290.825 100.265 ;
        RECT 278.540 100.065 290.825 100.205 ;
        RECT 278.540 100.020 279.190 100.065 ;
        RECT 281.840 100.020 282.430 100.065 ;
        RECT 268.540 99.865 268.830 99.910 ;
        RECT 272.120 99.865 272.410 99.910 ;
        RECT 273.955 99.865 274.245 99.910 ;
        RECT 268.540 99.725 274.245 99.865 ;
        RECT 268.540 99.680 268.830 99.725 ;
        RECT 272.120 99.680 272.410 99.725 ;
        RECT 273.955 99.680 274.245 99.725 ;
        RECT 275.345 99.865 275.635 99.910 ;
        RECT 277.180 99.865 277.470 99.910 ;
        RECT 280.760 99.865 281.050 99.910 ;
        RECT 275.345 99.725 281.050 99.865 ;
        RECT 275.345 99.680 275.635 99.725 ;
        RECT 277.180 99.680 277.470 99.725 ;
        RECT 280.760 99.680 281.050 99.725 ;
        RECT 281.840 99.705 282.130 100.020 ;
        RECT 282.685 100.005 283.005 100.065 ;
        RECT 290.505 100.005 290.825 100.065 ;
        RECT 283.145 99.865 283.465 99.925 ;
        RECT 284.985 99.865 285.305 99.925 ;
        RECT 285.920 99.865 286.210 99.910 ;
        RECT 283.145 99.725 284.755 99.865 ;
        RECT 283.145 99.665 283.465 99.725 ;
        RECT 244.045 99.525 244.365 99.585 ;
        RECT 248.185 99.525 248.505 99.585 ;
        RECT 248.660 99.525 248.950 99.570 ;
        RECT 229.875 99.385 231.855 99.525 ;
        RECT 213.225 99.185 213.545 99.245 ;
        RECT 217.915 99.185 218.055 99.385 ;
        RECT 211.015 99.045 212.995 99.185 ;
        RECT 205.520 99.000 205.810 99.045 ;
        RECT 208.640 99.000 208.930 99.045 ;
        RECT 210.530 99.000 210.820 99.045 ;
        RECT 209.545 98.845 209.865 98.905 ;
        RECT 205.035 98.705 209.865 98.845 ;
        RECT 193.445 98.645 193.765 98.705 ;
        RECT 202.660 98.660 202.950 98.705 ;
        RECT 204.485 98.645 204.805 98.705 ;
        RECT 209.545 98.645 209.865 98.705 ;
        RECT 210.005 98.845 210.325 98.905 ;
        RECT 212.320 98.845 212.610 98.890 ;
        RECT 210.005 98.705 212.610 98.845 ;
        RECT 212.855 98.845 212.995 99.045 ;
        RECT 213.225 99.045 218.055 99.185 ;
        RECT 218.250 99.185 218.540 99.230 ;
        RECT 220.140 99.185 220.430 99.230 ;
        RECT 223.260 99.185 223.550 99.230 ;
        RECT 218.250 99.045 223.550 99.185 ;
        RECT 213.225 98.985 213.545 99.045 ;
        RECT 218.250 99.000 218.540 99.045 ;
        RECT 220.140 99.000 220.430 99.045 ;
        RECT 223.260 99.000 223.550 99.045 ;
        RECT 229.325 98.845 229.645 98.905 ;
        RECT 212.855 98.705 229.645 98.845 ;
        RECT 210.005 98.645 210.325 98.705 ;
        RECT 212.320 98.660 212.610 98.705 ;
        RECT 229.325 98.645 229.645 98.705 ;
        RECT 231.165 98.645 231.485 98.905 ;
        RECT 231.715 98.845 231.855 99.385 ;
        RECT 244.045 99.385 248.950 99.525 ;
        RECT 244.045 99.325 244.365 99.385 ;
        RECT 248.185 99.325 248.505 99.385 ;
        RECT 248.660 99.340 248.950 99.385 ;
        RECT 249.565 99.525 249.885 99.585 ;
        RECT 255.100 99.525 255.390 99.570 ;
        RECT 255.545 99.525 255.865 99.585 ;
        RECT 258.780 99.525 259.070 99.570 ;
        RECT 249.565 99.385 259.070 99.525 ;
        RECT 249.565 99.325 249.885 99.385 ;
        RECT 255.100 99.340 255.390 99.385 ;
        RECT 255.545 99.325 255.865 99.385 ;
        RECT 258.780 99.340 259.070 99.385 ;
        RECT 259.685 99.525 260.005 99.585 ;
        RECT 269.805 99.525 270.125 99.585 ;
        RECT 259.685 99.385 270.125 99.525 ;
        RECT 259.685 99.325 260.005 99.385 ;
        RECT 269.805 99.325 270.125 99.385 ;
        RECT 274.420 99.525 274.710 99.570 ;
        RECT 274.880 99.525 275.170 99.570 ;
        RECT 274.420 99.385 275.170 99.525 ;
        RECT 274.420 99.340 274.710 99.385 ;
        RECT 274.880 99.340 275.170 99.385 ;
        RECT 240.790 99.185 241.080 99.230 ;
        RECT 242.680 99.185 242.970 99.230 ;
        RECT 245.800 99.185 246.090 99.230 ;
        RECT 240.790 99.045 246.090 99.185 ;
        RECT 240.790 99.000 241.080 99.045 ;
        RECT 242.680 99.000 242.970 99.045 ;
        RECT 245.800 99.000 246.090 99.045 ;
        RECT 249.105 99.185 249.425 99.245 ;
        RECT 256.940 99.185 257.230 99.230 ;
        RECT 249.105 99.045 257.230 99.185 ;
        RECT 249.105 98.985 249.425 99.045 ;
        RECT 256.940 99.000 257.230 99.045 ;
        RECT 268.540 99.185 268.830 99.230 ;
        RECT 271.660 99.185 271.950 99.230 ;
        RECT 273.550 99.185 273.840 99.230 ;
        RECT 268.540 99.045 273.840 99.185 ;
        RECT 268.540 99.000 268.830 99.045 ;
        RECT 271.660 99.000 271.950 99.045 ;
        RECT 273.550 99.000 273.840 99.045 ;
        RECT 244.965 98.845 245.285 98.905 ;
        RECT 231.715 98.705 245.285 98.845 ;
        RECT 244.965 98.645 245.285 98.705 ;
        RECT 251.880 98.845 252.170 98.890 ;
        RECT 256.005 98.845 256.325 98.905 ;
        RECT 251.880 98.705 256.325 98.845 ;
        RECT 251.880 98.660 252.170 98.705 ;
        RECT 256.005 98.645 256.325 98.705 ;
        RECT 259.225 98.845 259.545 98.905 ;
        RECT 263.825 98.845 264.145 98.905 ;
        RECT 259.225 98.705 264.145 98.845 ;
        RECT 259.225 98.645 259.545 98.705 ;
        RECT 263.825 98.645 264.145 98.705 ;
        RECT 265.665 98.845 265.985 98.905 ;
        RECT 267.965 98.845 268.285 98.905 ;
        RECT 265.665 98.705 268.285 98.845 ;
        RECT 274.955 98.845 275.095 99.340 ;
        RECT 276.245 99.325 276.565 99.585 ;
        RECT 283.605 99.325 283.925 99.585 ;
        RECT 284.615 99.570 284.755 99.725 ;
        RECT 284.985 99.725 286.210 99.865 ;
        RECT 284.985 99.665 285.305 99.725 ;
        RECT 285.920 99.680 286.210 99.725 ;
        RECT 288.205 99.665 288.525 99.925 ;
        RECT 291.425 99.665 291.745 99.925 ;
        RECT 284.540 99.340 284.830 99.570 ;
        RECT 285.445 99.325 285.765 99.585 ;
        RECT 275.750 99.185 276.040 99.230 ;
        RECT 277.640 99.185 277.930 99.230 ;
        RECT 280.760 99.185 281.050 99.230 ;
        RECT 275.750 99.045 281.050 99.185 ;
        RECT 283.695 99.185 283.835 99.325 ;
        RECT 289.140 99.185 289.430 99.230 ;
        RECT 283.695 99.045 289.430 99.185 ;
        RECT 275.750 99.000 276.040 99.045 ;
        RECT 277.640 99.000 277.930 99.045 ;
        RECT 280.760 99.000 281.050 99.045 ;
        RECT 289.140 99.000 289.430 99.045 ;
        RECT 279.005 98.845 279.325 98.905 ;
        RECT 274.955 98.705 279.325 98.845 ;
        RECT 265.665 98.645 265.985 98.705 ;
        RECT 267.965 98.645 268.285 98.705 ;
        RECT 279.005 98.645 279.325 98.705 ;
        RECT 281.765 98.845 282.085 98.905 ;
        RECT 283.620 98.845 283.910 98.890 ;
        RECT 281.765 98.705 283.910 98.845 ;
        RECT 281.765 98.645 282.085 98.705 ;
        RECT 283.620 98.660 283.910 98.705 ;
        RECT 284.525 98.845 284.845 98.905 ;
        RECT 292.895 98.845 293.035 100.405 ;
        RECT 298.325 100.345 298.645 100.405 ;
        RECT 299.705 100.545 300.025 100.605 ;
        RECT 302.925 100.545 303.245 100.605 ;
        RECT 303.400 100.545 303.690 100.590 ;
        RECT 299.705 100.405 301.775 100.545 ;
        RECT 299.705 100.345 300.025 100.405 ;
        RECT 294.645 100.205 294.965 100.265 ;
        RECT 293.815 100.065 294.965 100.205 ;
        RECT 293.815 99.910 293.955 100.065 ;
        RECT 294.645 100.005 294.965 100.065 ;
        RECT 297.400 100.205 298.050 100.250 ;
        RECT 301.000 100.205 301.290 100.250 ;
        RECT 297.400 100.065 301.290 100.205 ;
        RECT 301.635 100.205 301.775 100.405 ;
        RECT 302.925 100.405 303.690 100.545 ;
        RECT 302.925 100.345 303.245 100.405 ;
        RECT 303.400 100.360 303.690 100.405 ;
        RECT 304.305 100.545 304.625 100.605 ;
        RECT 305.700 100.545 305.990 100.590 ;
        RECT 304.305 100.405 305.990 100.545 ;
        RECT 304.305 100.345 304.625 100.405 ;
        RECT 305.700 100.360 305.990 100.405 ;
        RECT 306.605 100.545 306.925 100.605 ;
        RECT 308.000 100.545 308.290 100.590 ;
        RECT 306.605 100.405 308.290 100.545 ;
        RECT 306.605 100.345 306.925 100.405 ;
        RECT 308.000 100.360 308.290 100.405 ;
        RECT 301.635 100.065 304.995 100.205 ;
        RECT 297.400 100.020 298.050 100.065 ;
        RECT 300.700 100.020 301.290 100.065 ;
        RECT 293.740 99.680 294.030 99.910 ;
        RECT 294.205 99.865 294.495 99.910 ;
        RECT 296.040 99.865 296.330 99.910 ;
        RECT 299.620 99.865 299.910 99.910 ;
        RECT 294.205 99.725 299.910 99.865 ;
        RECT 294.205 99.680 294.495 99.725 ;
        RECT 296.040 99.680 296.330 99.725 ;
        RECT 299.620 99.680 299.910 99.725 ;
        RECT 300.700 99.865 300.990 100.020 ;
        RECT 302.925 99.865 303.245 99.925 ;
        RECT 304.855 99.910 304.995 100.065 ;
        RECT 300.700 99.725 303.245 99.865 ;
        RECT 300.700 99.705 300.990 99.725 ;
        RECT 295.120 99.525 295.410 99.570 ;
        RECT 297.865 99.525 298.185 99.585 ;
        RECT 295.120 99.385 298.185 99.525 ;
        RECT 295.120 99.340 295.410 99.385 ;
        RECT 297.865 99.325 298.185 99.385 ;
        RECT 298.325 99.525 298.645 99.585 ;
        RECT 300.715 99.525 300.855 99.705 ;
        RECT 302.925 99.665 303.245 99.725 ;
        RECT 304.320 99.680 304.610 99.910 ;
        RECT 304.780 99.680 305.070 99.910 ;
        RECT 305.685 99.865 306.005 99.925 ;
        RECT 307.080 99.865 307.370 99.910 ;
        RECT 305.685 99.725 307.370 99.865 ;
        RECT 298.325 99.385 300.855 99.525 ;
        RECT 304.395 99.525 304.535 99.680 ;
        RECT 305.685 99.665 306.005 99.725 ;
        RECT 307.080 99.680 307.370 99.725 ;
        RECT 305.225 99.525 305.545 99.585 ;
        RECT 304.395 99.385 305.545 99.525 ;
        RECT 298.325 99.325 298.645 99.385 ;
        RECT 305.225 99.325 305.545 99.385 ;
        RECT 294.610 99.185 294.900 99.230 ;
        RECT 296.500 99.185 296.790 99.230 ;
        RECT 299.620 99.185 299.910 99.230 ;
        RECT 294.610 99.045 299.910 99.185 ;
        RECT 294.610 99.000 294.900 99.045 ;
        RECT 296.500 99.000 296.790 99.045 ;
        RECT 299.620 99.000 299.910 99.045 ;
        RECT 284.525 98.705 293.035 98.845 ;
        RECT 296.945 98.845 297.265 98.905 ;
        RECT 302.480 98.845 302.770 98.890 ;
        RECT 296.945 98.705 302.770 98.845 ;
        RECT 284.525 98.645 284.845 98.705 ;
        RECT 296.945 98.645 297.265 98.705 ;
        RECT 302.480 98.660 302.770 98.705 ;
        RECT 162.095 98.025 311.135 98.505 ;
        RECT 167.175 97.825 167.465 97.870 ;
        RECT 176.425 97.825 176.745 97.885 ;
        RECT 167.175 97.685 176.745 97.825 ;
        RECT 167.175 97.640 167.465 97.685 ;
        RECT 176.425 97.625 176.745 97.685 ;
        RECT 187.465 97.825 187.785 97.885 ;
        RECT 193.460 97.825 193.750 97.870 ;
        RECT 187.465 97.685 193.750 97.825 ;
        RECT 187.465 97.625 187.785 97.685 ;
        RECT 193.460 97.640 193.750 97.685 ;
        RECT 195.745 97.825 196.065 97.885 ;
        RECT 210.925 97.825 211.245 97.885 ;
        RECT 195.745 97.685 211.245 97.825 ;
        RECT 195.745 97.625 196.065 97.685 ;
        RECT 210.925 97.625 211.245 97.685 ;
        RECT 211.860 97.825 212.150 97.870 ;
        RECT 214.145 97.825 214.465 97.885 ;
        RECT 211.860 97.685 214.465 97.825 ;
        RECT 211.860 97.640 212.150 97.685 ;
        RECT 214.145 97.625 214.465 97.685 ;
        RECT 220.125 97.825 220.445 97.885 ;
        RECT 220.600 97.825 220.890 97.870 ;
        RECT 220.125 97.685 220.890 97.825 ;
        RECT 220.125 97.625 220.445 97.685 ;
        RECT 220.600 97.640 220.890 97.685 ;
        RECT 226.105 97.625 226.425 97.885 ;
        RECT 229.325 97.825 229.645 97.885 ;
        RECT 255.545 97.825 255.865 97.885 ;
        RECT 257.860 97.825 258.150 97.870 ;
        RECT 229.325 97.685 244.735 97.825 ;
        RECT 229.325 97.625 229.645 97.685 ;
        RECT 166.730 97.485 167.020 97.530 ;
        RECT 168.620 97.485 168.910 97.530 ;
        RECT 171.740 97.485 172.030 97.530 ;
        RECT 174.585 97.485 174.905 97.545 ;
        RECT 185.130 97.485 185.420 97.530 ;
        RECT 187.020 97.485 187.310 97.530 ;
        RECT 190.140 97.485 190.430 97.530 ;
        RECT 222.440 97.485 222.730 97.530 ;
        RECT 166.730 97.345 172.030 97.485 ;
        RECT 166.730 97.300 167.020 97.345 ;
        RECT 168.620 97.300 168.910 97.345 ;
        RECT 171.740 97.300 172.030 97.345 ;
        RECT 173.065 97.345 184.475 97.485 ;
        RECT 165.860 97.145 166.150 97.190 ;
        RECT 173.065 97.145 173.205 97.345 ;
        RECT 174.585 97.285 174.905 97.345 ;
        RECT 165.860 97.005 173.205 97.145 ;
        RECT 178.740 97.145 179.030 97.190 ;
        RECT 179.645 97.145 179.965 97.205 ;
        RECT 184.335 97.190 184.475 97.345 ;
        RECT 185.130 97.345 190.430 97.485 ;
        RECT 185.130 97.300 185.420 97.345 ;
        RECT 187.020 97.300 187.310 97.345 ;
        RECT 190.140 97.300 190.430 97.345 ;
        RECT 190.775 97.345 207.015 97.485 ;
        RECT 181.500 97.145 181.790 97.190 ;
        RECT 178.740 97.005 181.790 97.145 ;
        RECT 165.860 96.960 166.150 97.005 ;
        RECT 178.740 96.960 179.030 97.005 ;
        RECT 179.645 96.945 179.965 97.005 ;
        RECT 181.500 96.960 181.790 97.005 ;
        RECT 184.260 96.960 184.550 97.190 ;
        RECT 187.465 97.145 187.785 97.205 ;
        RECT 190.775 97.145 190.915 97.345 ;
        RECT 187.465 97.005 190.915 97.145 ;
        RECT 192.525 97.145 192.845 97.205 ;
        RECT 196.220 97.145 196.510 97.190 ;
        RECT 198.045 97.145 198.365 97.205 ;
        RECT 192.525 97.005 196.510 97.145 ;
        RECT 187.465 96.945 187.785 97.005 ;
        RECT 192.525 96.945 192.845 97.005 ;
        RECT 196.220 96.960 196.510 97.005 ;
        RECT 196.755 97.005 198.365 97.145 ;
        RECT 164.940 96.620 165.230 96.850 ;
        RECT 166.325 96.805 166.615 96.850 ;
        RECT 168.160 96.805 168.450 96.850 ;
        RECT 171.740 96.805 172.030 96.850 ;
        RECT 166.325 96.665 172.030 96.805 ;
        RECT 166.325 96.620 166.615 96.665 ;
        RECT 168.160 96.620 168.450 96.665 ;
        RECT 171.740 96.620 172.030 96.665 ;
        RECT 165.015 96.465 165.155 96.620 ;
        RECT 168.605 96.465 168.925 96.525 ;
        RECT 172.820 96.510 173.110 96.825 ;
        RECT 182.405 96.605 182.725 96.865 ;
        RECT 183.325 96.605 183.645 96.865 ;
        RECT 183.800 96.620 184.090 96.850 ;
        RECT 184.725 96.805 185.015 96.850 ;
        RECT 186.560 96.805 186.850 96.850 ;
        RECT 190.140 96.805 190.430 96.850 ;
        RECT 184.725 96.665 190.430 96.805 ;
        RECT 184.725 96.620 185.015 96.665 ;
        RECT 186.560 96.620 186.850 96.665 ;
        RECT 190.140 96.620 190.430 96.665 ;
        RECT 165.015 96.325 168.925 96.465 ;
        RECT 168.605 96.265 168.925 96.325 ;
        RECT 169.520 96.465 170.170 96.510 ;
        RECT 172.820 96.465 173.410 96.510 ;
        RECT 174.125 96.465 174.445 96.525 ;
        RECT 180.105 96.465 180.425 96.525 ;
        RECT 169.520 96.325 174.445 96.465 ;
        RECT 169.520 96.280 170.170 96.325 ;
        RECT 173.120 96.280 173.410 96.325 ;
        RECT 174.125 96.265 174.445 96.325 ;
        RECT 174.675 96.325 180.425 96.465 ;
        RECT 183.875 96.465 184.015 96.620 ;
        RECT 185.165 96.465 185.485 96.525 ;
        RECT 183.875 96.325 185.485 96.465 ;
        RECT 164.020 96.125 164.310 96.170 ;
        RECT 170.905 96.125 171.225 96.185 ;
        RECT 174.675 96.170 174.815 96.325 ;
        RECT 180.105 96.265 180.425 96.325 ;
        RECT 185.165 96.265 185.485 96.325 ;
        RECT 185.625 96.265 185.945 96.525 ;
        RECT 191.220 96.510 191.510 96.825 ;
        RECT 195.745 96.605 196.065 96.865 ;
        RECT 187.920 96.465 188.570 96.510 ;
        RECT 191.220 96.465 191.810 96.510 ;
        RECT 196.755 96.465 196.895 97.005 ;
        RECT 198.045 96.945 198.365 97.005 ;
        RECT 197.125 96.805 197.445 96.865 ;
        RECT 199.440 96.805 199.730 96.850 ;
        RECT 197.125 96.665 199.730 96.805 ;
        RECT 197.125 96.605 197.445 96.665 ;
        RECT 199.440 96.620 199.730 96.665 ;
        RECT 203.565 96.605 203.885 96.865 ;
        RECT 204.960 96.805 205.250 96.850 ;
        RECT 205.865 96.805 206.185 96.865 ;
        RECT 204.960 96.665 206.185 96.805 ;
        RECT 204.960 96.620 205.250 96.665 ;
        RECT 205.865 96.605 206.185 96.665 ;
        RECT 206.325 96.605 206.645 96.865 ;
        RECT 206.875 96.850 207.015 97.345 ;
        RECT 222.440 97.345 224.495 97.485 ;
        RECT 222.440 97.300 222.730 97.345 ;
        RECT 211.845 97.145 212.165 97.205 ;
        RECT 208.255 97.005 212.165 97.145 ;
        RECT 208.255 96.850 208.395 97.005 ;
        RECT 211.845 96.945 212.165 97.005 ;
        RECT 224.355 97.145 224.495 97.345 ;
        RECT 243.125 97.285 243.445 97.545 ;
        RECT 232.545 97.145 232.865 97.205 ;
        RECT 224.355 97.005 232.865 97.145 ;
        RECT 206.800 96.805 207.090 96.850 ;
        RECT 206.800 96.665 207.935 96.805 ;
        RECT 206.800 96.620 207.090 96.665 ;
        RECT 187.920 96.325 196.895 96.465 ;
        RECT 204.485 96.465 204.805 96.525 ;
        RECT 204.485 96.325 206.555 96.465 ;
        RECT 187.920 96.280 188.570 96.325 ;
        RECT 191.520 96.280 191.810 96.325 ;
        RECT 164.020 95.985 171.225 96.125 ;
        RECT 164.020 95.940 164.310 95.985 ;
        RECT 170.905 95.925 171.225 95.985 ;
        RECT 174.600 95.940 174.890 96.170 ;
        RECT 175.505 95.925 175.825 96.185 ;
        RECT 177.345 95.925 177.665 96.185 ;
        RECT 177.820 96.125 178.110 96.170 ;
        RECT 186.085 96.125 186.405 96.185 ;
        RECT 177.820 95.985 186.405 96.125 ;
        RECT 177.820 95.940 178.110 95.985 ;
        RECT 186.085 95.925 186.405 95.985 ;
        RECT 187.465 96.125 187.785 96.185 ;
        RECT 192.155 96.125 192.295 96.325 ;
        RECT 204.485 96.265 204.805 96.325 ;
        RECT 187.465 95.985 192.295 96.125 ;
        RECT 193.000 96.125 193.290 96.170 ;
        RECT 193.905 96.125 194.225 96.185 ;
        RECT 193.000 95.985 194.225 96.125 ;
        RECT 187.465 95.925 187.785 95.985 ;
        RECT 193.000 95.940 193.290 95.985 ;
        RECT 193.905 95.925 194.225 95.985 ;
        RECT 195.285 95.925 195.605 96.185 ;
        RECT 198.505 96.125 198.825 96.185 ;
        RECT 202.660 96.125 202.950 96.170 ;
        RECT 198.505 95.985 202.950 96.125 ;
        RECT 198.505 95.925 198.825 95.985 ;
        RECT 202.660 95.940 202.950 95.985 ;
        RECT 205.405 95.925 205.725 96.185 ;
        RECT 206.415 96.125 206.555 96.325 ;
        RECT 207.245 96.265 207.565 96.525 ;
        RECT 207.795 96.465 207.935 96.665 ;
        RECT 208.180 96.620 208.470 96.850 ;
        RECT 209.100 96.620 209.390 96.850 ;
        RECT 209.545 96.805 209.865 96.865 ;
        RECT 221.505 96.805 221.825 96.865 ;
        RECT 209.545 96.665 221.825 96.805 ;
        RECT 208.625 96.465 208.945 96.525 ;
        RECT 207.795 96.325 208.945 96.465 ;
        RECT 208.625 96.265 208.945 96.325 ;
        RECT 209.175 96.465 209.315 96.620 ;
        RECT 209.545 96.605 209.865 96.665 ;
        RECT 221.505 96.605 221.825 96.665 ;
        RECT 222.885 96.605 223.205 96.865 ;
        RECT 224.355 96.850 224.495 97.005 ;
        RECT 232.545 96.945 232.865 97.005 ;
        RECT 244.595 97.145 244.735 97.685 ;
        RECT 255.545 97.685 258.150 97.825 ;
        RECT 255.545 97.625 255.865 97.685 ;
        RECT 257.860 97.640 258.150 97.685 ;
        RECT 276.245 97.825 276.565 97.885 ;
        RECT 277.640 97.825 277.930 97.870 ;
        RECT 276.245 97.685 277.930 97.825 ;
        RECT 276.245 97.625 276.565 97.685 ;
        RECT 277.640 97.640 277.930 97.685 ;
        RECT 282.225 97.825 282.545 97.885 ;
        RECT 286.365 97.825 286.685 97.885 ;
        RECT 289.140 97.825 289.430 97.870 ;
        RECT 282.225 97.685 286.135 97.825 ;
        RECT 282.225 97.625 282.545 97.685 ;
        RECT 259.685 97.485 260.005 97.545 ;
        RECT 279.890 97.485 280.180 97.530 ;
        RECT 281.780 97.485 282.070 97.530 ;
        RECT 284.900 97.485 285.190 97.530 ;
        RECT 254.715 97.345 260.005 97.485 ;
        RECT 244.595 97.005 248.900 97.145 ;
        RECT 223.360 96.620 223.650 96.850 ;
        RECT 224.280 96.620 224.570 96.850 ;
        RECT 225.200 96.805 225.490 96.850 ;
        RECT 225.645 96.805 225.965 96.865 ;
        RECT 225.200 96.665 225.965 96.805 ;
        RECT 225.200 96.620 225.490 96.665 ;
        RECT 216.905 96.465 217.225 96.525 ;
        RECT 223.435 96.465 223.575 96.620 ;
        RECT 225.645 96.605 225.965 96.665 ;
        RECT 226.565 96.805 226.885 96.865 ;
        RECT 227.730 96.805 228.020 96.850 ;
        RECT 226.565 96.665 228.020 96.805 ;
        RECT 226.565 96.605 226.885 96.665 ;
        RECT 227.730 96.620 228.020 96.665 ;
        RECT 228.405 96.605 228.725 96.865 ;
        RECT 229.795 96.620 230.085 96.850 ;
        RECT 230.260 96.805 230.550 96.850 ;
        RECT 241.285 96.805 241.605 96.865 ;
        RECT 230.260 96.665 241.605 96.805 ;
        RECT 230.260 96.620 230.550 96.665 ;
        RECT 209.175 96.325 223.575 96.465 ;
        RECT 224.740 96.465 225.030 96.510 ;
        RECT 224.740 96.325 228.635 96.465 ;
        RECT 209.175 96.125 209.315 96.325 ;
        RECT 216.905 96.265 217.225 96.325 ;
        RECT 224.740 96.280 225.030 96.325 ;
        RECT 206.415 95.985 209.315 96.125 ;
        RECT 210.005 96.125 210.325 96.185 ;
        RECT 213.225 96.125 213.545 96.185 ;
        RECT 210.005 95.985 213.545 96.125 ;
        RECT 210.005 95.925 210.325 95.985 ;
        RECT 213.225 95.925 213.545 95.985 ;
        RECT 227.025 95.925 227.345 96.185 ;
        RECT 228.495 96.125 228.635 96.325 ;
        RECT 228.865 96.265 229.185 96.525 ;
        RECT 229.875 96.465 230.015 96.620 ;
        RECT 241.285 96.605 241.605 96.665 ;
        RECT 241.745 96.805 242.065 96.865 ;
        RECT 244.060 96.805 244.350 96.850 ;
        RECT 241.745 96.665 244.350 96.805 ;
        RECT 244.595 96.805 244.735 97.005 ;
        RECT 244.980 96.805 245.270 96.850 ;
        RECT 244.595 96.665 245.270 96.805 ;
        RECT 241.745 96.605 242.065 96.665 ;
        RECT 244.060 96.620 244.350 96.665 ;
        RECT 244.980 96.620 245.270 96.665 ;
        RECT 245.425 96.805 245.745 96.865 ;
        RECT 245.900 96.805 246.190 96.850 ;
        RECT 245.425 96.665 246.190 96.805 ;
        RECT 245.425 96.605 245.745 96.665 ;
        RECT 245.900 96.620 246.190 96.665 ;
        RECT 246.345 96.605 246.665 96.865 ;
        RECT 247.100 96.805 247.390 96.850 ;
        RECT 247.100 96.620 247.495 96.805 ;
        RECT 235.765 96.465 236.085 96.525 ;
        RECT 229.875 96.325 236.085 96.465 ;
        RECT 229.875 96.125 230.015 96.325 ;
        RECT 235.765 96.265 236.085 96.325 ;
        RECT 244.505 96.265 244.825 96.525 ;
        RECT 228.495 95.985 230.015 96.125 ;
        RECT 247.355 96.125 247.495 96.620 ;
        RECT 248.185 96.605 248.505 96.865 ;
        RECT 248.760 96.850 248.900 97.005 ;
        RECT 248.685 96.620 248.975 96.850 ;
        RECT 253.695 96.805 253.985 96.850 ;
        RECT 254.715 96.805 254.855 97.345 ;
        RECT 259.685 97.285 260.005 97.345 ;
        RECT 278.635 97.345 279.695 97.485 ;
        RECT 272.105 97.145 272.425 97.205 ;
        RECT 274.420 97.145 274.710 97.190 ;
        RECT 277.165 97.145 277.485 97.205 ;
        RECT 272.105 97.005 277.485 97.145 ;
        RECT 272.105 96.945 272.425 97.005 ;
        RECT 274.420 96.960 274.710 97.005 ;
        RECT 277.165 96.945 277.485 97.005 ;
        RECT 255.545 96.805 255.865 96.865 ;
        RECT 253.695 96.665 254.855 96.805 ;
        RECT 255.350 96.665 255.865 96.805 ;
        RECT 253.695 96.620 253.985 96.665 ;
        RECT 255.545 96.605 255.865 96.665 ;
        RECT 256.005 96.605 256.325 96.865 ;
        RECT 257.385 96.805 257.705 96.865 ;
        RECT 259.240 96.805 259.530 96.850 ;
        RECT 259.685 96.805 260.005 96.865 ;
        RECT 257.385 96.665 257.900 96.805 ;
        RECT 259.240 96.665 260.005 96.805 ;
        RECT 257.385 96.605 257.705 96.665 ;
        RECT 259.240 96.620 259.530 96.665 ;
        RECT 259.685 96.605 260.005 96.665 ;
        RECT 260.145 96.605 260.465 96.865 ;
        RECT 260.605 96.805 260.925 96.865 ;
        RECT 267.505 96.805 267.825 96.865 ;
        RECT 269.345 96.805 269.665 96.865 ;
        RECT 275.800 96.805 276.090 96.850 ;
        RECT 260.605 96.665 266.355 96.805 ;
        RECT 260.605 96.605 260.925 96.665 ;
        RECT 247.725 96.265 248.045 96.525 ;
        RECT 254.165 96.465 254.485 96.525 ;
        RECT 249.195 96.325 254.485 96.465 ;
        RECT 249.195 96.125 249.335 96.325 ;
        RECT 254.165 96.265 254.485 96.325 ;
        RECT 254.640 96.280 254.930 96.510 ;
        RECT 255.635 96.465 255.775 96.605 ;
        RECT 265.665 96.465 265.985 96.525 ;
        RECT 255.635 96.325 265.985 96.465 ;
        RECT 266.215 96.465 266.355 96.665 ;
        RECT 267.505 96.665 276.090 96.805 ;
        RECT 267.505 96.605 267.825 96.665 ;
        RECT 269.345 96.605 269.665 96.665 ;
        RECT 275.800 96.620 276.090 96.665 ;
        RECT 275.340 96.465 275.630 96.510 ;
        RECT 278.635 96.465 278.775 97.345 ;
        RECT 279.005 96.945 279.325 97.205 ;
        RECT 279.555 97.145 279.695 97.345 ;
        RECT 279.890 97.345 285.190 97.485 ;
        RECT 285.995 97.485 286.135 97.685 ;
        RECT 286.365 97.685 289.430 97.825 ;
        RECT 286.365 97.625 286.685 97.685 ;
        RECT 289.140 97.640 289.430 97.685 ;
        RECT 290.045 97.625 290.365 97.885 ;
        RECT 303.400 97.825 303.690 97.870 ;
        RECT 307.985 97.825 308.305 97.885 ;
        RECT 303.400 97.685 308.305 97.825 ;
        RECT 303.400 97.640 303.690 97.685 ;
        RECT 295.530 97.485 295.820 97.530 ;
        RECT 297.420 97.485 297.710 97.530 ;
        RECT 300.540 97.485 300.830 97.530 ;
        RECT 285.995 97.345 292.575 97.485 ;
        RECT 279.890 97.300 280.180 97.345 ;
        RECT 281.780 97.300 282.070 97.345 ;
        RECT 284.900 97.300 285.190 97.345 ;
        RECT 292.435 97.205 292.575 97.345 ;
        RECT 295.530 97.345 300.830 97.485 ;
        RECT 295.530 97.300 295.820 97.345 ;
        RECT 297.420 97.300 297.710 97.345 ;
        RECT 300.540 97.300 300.830 97.345 ;
        RECT 304.320 97.300 304.610 97.530 ;
        RECT 286.825 97.145 287.145 97.205 ;
        RECT 279.555 97.005 287.145 97.145 ;
        RECT 286.825 96.945 287.145 97.005 ;
        RECT 292.345 96.945 292.665 97.205 ;
        RECT 293.265 96.945 293.585 97.205 ;
        RECT 296.040 97.145 296.330 97.190 ;
        RECT 304.395 97.145 304.535 97.300 ;
        RECT 296.040 97.005 304.535 97.145 ;
        RECT 296.040 96.960 296.330 97.005 ;
        RECT 279.485 96.805 279.775 96.850 ;
        RECT 281.320 96.805 281.610 96.850 ;
        RECT 284.900 96.805 285.190 96.850 ;
        RECT 279.485 96.665 285.190 96.805 ;
        RECT 279.485 96.620 279.775 96.665 ;
        RECT 281.320 96.620 281.610 96.665 ;
        RECT 284.900 96.620 285.190 96.665 ;
        RECT 266.215 96.325 278.775 96.465 ;
        RECT 279.925 96.465 280.245 96.525 ;
        RECT 282.685 96.510 283.005 96.525 ;
        RECT 285.980 96.510 286.270 96.825 ;
        RECT 288.220 96.805 288.510 96.850 ;
        RECT 286.915 96.665 288.510 96.805 ;
        RECT 280.400 96.465 280.690 96.510 ;
        RECT 279.925 96.325 280.690 96.465 ;
        RECT 247.355 95.985 249.335 96.125 ;
        RECT 249.580 96.125 249.870 96.170 ;
        RECT 251.405 96.125 251.725 96.185 ;
        RECT 249.580 95.985 251.725 96.125 ;
        RECT 249.580 95.940 249.870 95.985 ;
        RECT 251.405 95.925 251.725 95.985 ;
        RECT 252.785 95.925 253.105 96.185 ;
        RECT 253.245 96.125 253.565 96.185 ;
        RECT 254.715 96.125 254.855 96.280 ;
        RECT 265.665 96.265 265.985 96.325 ;
        RECT 275.340 96.280 275.630 96.325 ;
        RECT 279.925 96.265 280.245 96.325 ;
        RECT 280.400 96.280 280.690 96.325 ;
        RECT 282.680 96.465 283.330 96.510 ;
        RECT 285.980 96.465 286.570 96.510 ;
        RECT 282.680 96.325 286.570 96.465 ;
        RECT 282.680 96.280 283.330 96.325 ;
        RECT 286.280 96.280 286.570 96.325 ;
        RECT 282.685 96.265 283.005 96.280 ;
        RECT 257.385 96.125 257.705 96.185 ;
        RECT 253.245 95.985 257.705 96.125 ;
        RECT 253.245 95.925 253.565 95.985 ;
        RECT 257.385 95.925 257.705 95.985 ;
        RECT 278.085 96.125 278.405 96.185 ;
        RECT 284.525 96.125 284.845 96.185 ;
        RECT 278.085 95.985 284.845 96.125 ;
        RECT 278.085 95.925 278.405 95.985 ;
        RECT 284.525 95.925 284.845 95.985 ;
        RECT 284.985 96.125 285.305 96.185 ;
        RECT 286.915 96.125 287.055 96.665 ;
        RECT 288.220 96.620 288.510 96.665 ;
        RECT 294.645 96.605 294.965 96.865 ;
        RECT 306.235 96.850 306.375 97.685 ;
        RECT 307.985 97.625 308.305 97.685 ;
        RECT 307.525 96.945 307.845 97.205 ;
        RECT 295.125 96.805 295.415 96.850 ;
        RECT 296.960 96.805 297.250 96.850 ;
        RECT 300.540 96.805 300.830 96.850 ;
        RECT 295.125 96.665 300.830 96.805 ;
        RECT 295.125 96.620 295.415 96.665 ;
        RECT 296.960 96.620 297.250 96.665 ;
        RECT 300.540 96.620 300.830 96.665 ;
        RECT 290.505 96.465 290.825 96.525 ;
        RECT 301.620 96.510 301.910 96.825 ;
        RECT 306.160 96.620 306.450 96.850 ;
        RECT 298.320 96.465 298.970 96.510 ;
        RECT 301.620 96.465 302.210 96.510 ;
        RECT 290.505 96.325 302.210 96.465 ;
        RECT 290.505 96.265 290.825 96.325 ;
        RECT 284.985 95.985 287.055 96.125 ;
        RECT 284.985 95.925 285.305 95.985 ;
        RECT 287.745 95.925 288.065 96.185 ;
        RECT 291.885 95.925 292.205 96.185 ;
        RECT 297.955 96.125 298.095 96.325 ;
        RECT 298.320 96.280 298.970 96.325 ;
        RECT 301.920 96.280 302.210 96.325 ;
        RECT 306.605 96.265 306.925 96.525 ;
        RECT 299.245 96.125 299.565 96.185 ;
        RECT 297.955 95.985 299.565 96.125 ;
        RECT 299.245 95.925 299.565 95.985 ;
        RECT 162.095 95.305 311.135 95.785 ;
        RECT 166.765 95.105 167.085 95.165 ;
        RECT 176.885 95.105 177.205 95.165 ;
        RECT 166.765 94.965 177.205 95.105 ;
        RECT 166.765 94.905 167.085 94.965 ;
        RECT 169.155 94.470 169.295 94.965 ;
        RECT 176.885 94.905 177.205 94.965 ;
        RECT 177.345 95.105 177.665 95.165 ;
        RECT 177.820 95.105 178.110 95.150 ;
        RECT 183.785 95.105 184.105 95.165 ;
        RECT 177.345 94.965 184.105 95.105 ;
        RECT 177.345 94.905 177.665 94.965 ;
        RECT 177.820 94.920 178.110 94.965 ;
        RECT 183.785 94.905 184.105 94.965 ;
        RECT 185.625 95.105 185.945 95.165 ;
        RECT 188.400 95.105 188.690 95.150 ;
        RECT 185.625 94.965 188.690 95.105 ;
        RECT 185.625 94.905 185.945 94.965 ;
        RECT 188.400 94.920 188.690 94.965 ;
        RECT 190.240 95.105 190.530 95.150 ;
        RECT 193.905 95.105 194.225 95.165 ;
        RECT 190.240 94.965 194.225 95.105 ;
        RECT 190.240 94.920 190.530 94.965 ;
        RECT 193.905 94.905 194.225 94.965 ;
        RECT 208.165 94.905 208.485 95.165 ;
        RECT 208.625 95.105 208.945 95.165 ;
        RECT 225.185 95.105 225.505 95.165 ;
        RECT 232.085 95.105 232.405 95.165 ;
        RECT 208.625 94.965 224.955 95.105 ;
        RECT 208.625 94.905 208.945 94.965 ;
        RECT 172.740 94.765 173.390 94.810 ;
        RECT 176.340 94.765 176.630 94.810 ;
        RECT 172.740 94.625 176.630 94.765 ;
        RECT 172.740 94.580 173.390 94.625 ;
        RECT 176.040 94.580 176.630 94.625 ;
        RECT 186.085 94.765 186.405 94.825 ;
        RECT 190.700 94.765 190.990 94.810 ;
        RECT 192.985 94.765 193.305 94.825 ;
        RECT 186.085 94.625 193.305 94.765 ;
        RECT 164.940 94.425 165.230 94.470 ;
        RECT 164.940 94.285 168.835 94.425 ;
        RECT 164.940 94.240 165.230 94.285 ;
        RECT 164.005 93.205 164.325 93.465 ;
        RECT 168.695 93.405 168.835 94.285 ;
        RECT 169.080 94.240 169.370 94.470 ;
        RECT 169.545 94.425 169.835 94.470 ;
        RECT 171.380 94.425 171.670 94.470 ;
        RECT 174.960 94.425 175.250 94.470 ;
        RECT 169.545 94.285 175.250 94.425 ;
        RECT 169.545 94.240 169.835 94.285 ;
        RECT 171.380 94.240 171.670 94.285 ;
        RECT 174.960 94.240 175.250 94.285 ;
        RECT 176.040 94.265 176.330 94.580 ;
        RECT 186.085 94.565 186.405 94.625 ;
        RECT 190.700 94.580 190.990 94.625 ;
        RECT 192.985 94.565 193.305 94.625 ;
        RECT 200.345 94.765 200.665 94.825 ;
        RECT 208.255 94.765 208.395 94.905 ;
        RECT 224.815 94.825 224.955 94.965 ;
        RECT 225.185 94.965 225.875 95.105 ;
        RECT 225.185 94.905 225.505 94.965 ;
        RECT 210.480 94.765 210.770 94.810 ;
        RECT 200.345 94.625 207.935 94.765 ;
        RECT 208.255 94.625 210.770 94.765 ;
        RECT 200.345 94.565 200.665 94.625 ;
        RECT 183.325 94.425 183.645 94.485 ;
        RECT 185.165 94.425 185.485 94.485 ;
        RECT 183.325 94.285 184.935 94.425 ;
        RECT 170.460 94.085 170.750 94.130 ;
        RECT 175.505 94.085 175.825 94.145 ;
        RECT 170.460 93.945 175.825 94.085 ;
        RECT 170.460 93.900 170.750 93.945 ;
        RECT 175.505 93.885 175.825 93.945 ;
        RECT 169.950 93.745 170.240 93.790 ;
        RECT 171.840 93.745 172.130 93.790 ;
        RECT 174.960 93.745 175.250 93.790 ;
        RECT 169.950 93.605 175.250 93.745 ;
        RECT 169.950 93.560 170.240 93.605 ;
        RECT 171.840 93.560 172.130 93.605 ;
        RECT 174.960 93.560 175.250 93.605 ;
        RECT 173.665 93.405 173.985 93.465 ;
        RECT 168.695 93.265 173.985 93.405 ;
        RECT 173.665 93.205 173.985 93.265 ;
        RECT 174.125 93.405 174.445 93.465 ;
        RECT 176.055 93.405 176.195 94.265 ;
        RECT 183.325 94.225 183.645 94.285 ;
        RECT 184.795 94.085 184.935 94.285 ;
        RECT 185.165 94.285 193.215 94.425 ;
        RECT 185.165 94.225 185.485 94.285 ;
        RECT 191.620 94.085 191.910 94.130 ;
        RECT 192.525 94.085 192.845 94.145 ;
        RECT 184.795 93.945 187.235 94.085 ;
        RECT 187.095 93.745 187.235 93.945 ;
        RECT 191.620 93.945 192.845 94.085 ;
        RECT 193.075 94.085 193.215 94.285 ;
        RECT 193.445 94.225 193.765 94.485 ;
        RECT 194.380 94.425 194.670 94.470 ;
        RECT 205.405 94.425 205.725 94.485 ;
        RECT 207.260 94.425 207.550 94.470 ;
        RECT 194.380 94.285 205.175 94.425 ;
        RECT 194.380 94.240 194.670 94.285 ;
        RECT 194.840 94.085 195.130 94.130 ;
        RECT 196.665 94.085 196.985 94.145 ;
        RECT 193.075 93.945 196.985 94.085 ;
        RECT 205.035 94.085 205.175 94.285 ;
        RECT 205.405 94.285 207.550 94.425 ;
        RECT 205.405 94.225 205.725 94.285 ;
        RECT 207.260 94.240 207.550 94.285 ;
        RECT 207.795 94.085 207.935 94.625 ;
        RECT 210.480 94.580 210.770 94.625 ;
        RECT 224.725 94.765 225.045 94.825 ;
        RECT 225.735 94.810 225.875 94.965 ;
        RECT 227.115 94.965 232.405 95.105 ;
        RECT 224.725 94.625 225.415 94.765 ;
        RECT 224.725 94.565 225.045 94.625 ;
        RECT 208.625 94.225 208.945 94.485 ;
        RECT 209.085 94.225 209.405 94.485 ;
        RECT 210.005 94.225 210.325 94.485 ;
        RECT 210.925 94.425 211.245 94.485 ;
        RECT 225.275 94.470 225.415 94.625 ;
        RECT 225.660 94.580 225.950 94.810 ;
        RECT 210.925 94.285 224.955 94.425 ;
        RECT 210.925 94.225 211.245 94.285 ;
        RECT 224.815 94.085 224.955 94.285 ;
        RECT 225.200 94.240 225.490 94.470 ;
        RECT 226.105 94.225 226.425 94.485 ;
        RECT 227.115 94.470 227.255 94.965 ;
        RECT 232.085 94.905 232.405 94.965 ;
        RECT 241.285 94.905 241.605 95.165 ;
        RECT 244.505 95.105 244.825 95.165 ;
        RECT 244.505 94.965 246.575 95.105 ;
        RECT 244.505 94.905 244.825 94.965 ;
        RECT 246.435 94.810 246.575 94.965 ;
        RECT 248.185 94.905 248.505 95.165 ;
        RECT 268.425 95.105 268.745 95.165 ;
        RECT 248.735 94.965 268.745 95.105 ;
        RECT 228.420 94.765 228.710 94.810 ;
        RECT 245.900 94.765 246.190 94.810 ;
        RECT 228.420 94.625 246.190 94.765 ;
        RECT 228.420 94.580 228.710 94.625 ;
        RECT 245.900 94.580 246.190 94.625 ;
        RECT 246.360 94.765 246.650 94.810 ;
        RECT 248.735 94.765 248.875 94.965 ;
        RECT 268.425 94.905 268.745 94.965 ;
        RECT 277.165 94.905 277.485 95.165 ;
        RECT 279.925 94.905 280.245 95.165 ;
        RECT 282.225 94.905 282.545 95.165 ;
        RECT 283.605 95.105 283.925 95.165 ;
        RECT 288.205 95.105 288.525 95.165 ;
        RECT 283.605 94.965 288.525 95.105 ;
        RECT 283.605 94.905 283.925 94.965 ;
        RECT 288.205 94.905 288.525 94.965 ;
        RECT 296.040 94.920 296.330 95.150 ;
        RECT 246.360 94.625 248.875 94.765 ;
        RECT 249.580 94.765 249.870 94.810 ;
        RECT 255.545 94.765 255.865 94.825 ;
        RECT 259.700 94.765 259.990 94.810 ;
        RECT 262.445 94.765 262.765 94.825 ;
        RECT 263.380 94.765 263.670 94.810 ;
        RECT 249.580 94.625 255.865 94.765 ;
        RECT 246.360 94.580 246.650 94.625 ;
        RECT 249.580 94.580 249.870 94.625 ;
        RECT 227.040 94.240 227.330 94.470 ;
        RECT 227.485 94.225 227.805 94.485 ;
        RECT 228.495 94.085 228.635 94.580 ;
        RECT 255.545 94.565 255.865 94.625 ;
        RECT 256.095 94.625 259.990 94.765 ;
        RECT 228.880 94.240 229.170 94.470 ;
        RECT 229.340 94.425 229.630 94.470 ;
        RECT 230.245 94.425 230.565 94.485 ;
        RECT 229.340 94.285 230.565 94.425 ;
        RECT 229.340 94.240 229.630 94.285 ;
        RECT 205.035 93.945 207.475 94.085 ;
        RECT 207.795 93.945 224.495 94.085 ;
        RECT 224.815 93.945 228.635 94.085 ;
        RECT 191.620 93.900 191.910 93.945 ;
        RECT 192.525 93.885 192.845 93.945 ;
        RECT 194.840 93.900 195.130 93.945 ;
        RECT 196.665 93.885 196.985 93.945 ;
        RECT 191.145 93.745 191.465 93.805 ;
        RECT 204.485 93.745 204.805 93.805 ;
        RECT 207.335 93.745 207.475 93.945 ;
        RECT 209.545 93.745 209.865 93.805 ;
        RECT 210.925 93.745 211.245 93.805 ;
        RECT 187.095 93.605 207.015 93.745 ;
        RECT 207.335 93.605 211.245 93.745 ;
        RECT 224.355 93.745 224.495 93.945 ;
        RECT 225.185 93.745 225.505 93.805 ;
        RECT 227.485 93.745 227.805 93.805 ;
        RECT 224.355 93.605 227.805 93.745 ;
        RECT 191.145 93.545 191.465 93.605 ;
        RECT 204.485 93.545 204.805 93.605 ;
        RECT 187.465 93.405 187.785 93.465 ;
        RECT 174.125 93.265 187.785 93.405 ;
        RECT 174.125 93.205 174.445 93.265 ;
        RECT 187.465 93.205 187.785 93.265 ;
        RECT 206.325 93.205 206.645 93.465 ;
        RECT 206.875 93.405 207.015 93.605 ;
        RECT 209.545 93.545 209.865 93.605 ;
        RECT 210.925 93.545 211.245 93.605 ;
        RECT 225.185 93.545 225.505 93.605 ;
        RECT 227.485 93.545 227.805 93.605 ;
        RECT 228.405 93.745 228.725 93.805 ;
        RECT 228.955 93.745 229.095 94.240 ;
        RECT 230.245 94.225 230.565 94.285 ;
        RECT 239.445 94.425 239.765 94.485 ;
        RECT 241.990 94.425 242.280 94.470 ;
        RECT 239.445 94.285 242.280 94.425 ;
        RECT 239.445 94.225 239.765 94.285 ;
        RECT 241.990 94.240 242.280 94.285 ;
        RECT 242.665 94.225 242.985 94.485 ;
        RECT 243.125 94.225 243.445 94.485 ;
        RECT 244.045 94.425 244.365 94.485 ;
        RECT 243.850 94.285 244.365 94.425 ;
        RECT 244.045 94.225 244.365 94.285 ;
        RECT 244.505 94.225 244.825 94.485 ;
        RECT 244.980 94.240 245.270 94.470 ;
        RECT 245.425 94.425 245.745 94.485 ;
        RECT 246.820 94.425 247.110 94.470 ;
        RECT 247.725 94.425 248.045 94.485 ;
        RECT 249.105 94.470 249.425 94.485 ;
        RECT 249.095 94.425 249.425 94.470 ;
        RECT 245.425 94.285 248.045 94.425 ;
        RECT 248.910 94.285 249.425 94.425 ;
        RECT 242.755 94.085 242.895 94.225 ;
        RECT 245.055 94.085 245.195 94.240 ;
        RECT 245.425 94.225 245.745 94.285 ;
        RECT 246.820 94.240 247.110 94.285 ;
        RECT 247.725 94.225 248.045 94.285 ;
        RECT 249.095 94.240 249.425 94.285 ;
        RECT 249.105 94.225 249.425 94.240 ;
        RECT 250.025 94.225 250.345 94.485 ;
        RECT 250.945 94.425 251.265 94.485 ;
        RECT 250.750 94.285 251.265 94.425 ;
        RECT 250.945 94.225 251.265 94.285 ;
        RECT 251.405 94.225 251.725 94.485 ;
        RECT 254.165 94.425 254.485 94.485 ;
        RECT 256.095 94.425 256.235 94.625 ;
        RECT 259.700 94.580 259.990 94.625 ;
        RECT 260.235 94.625 262.215 94.765 ;
        RECT 260.235 94.485 260.375 94.625 ;
        RECT 254.165 94.285 256.235 94.425 ;
        RECT 256.465 94.425 256.785 94.485 ;
        RECT 259.225 94.470 259.545 94.485 ;
        RECT 258.320 94.425 258.610 94.470 ;
        RECT 256.465 94.285 258.610 94.425 ;
        RECT 254.165 94.225 254.485 94.285 ;
        RECT 256.465 94.225 256.785 94.285 ;
        RECT 258.320 94.240 258.610 94.285 ;
        RECT 259.060 94.240 259.545 94.470 ;
        RECT 259.225 94.225 259.545 94.240 ;
        RECT 260.145 94.225 260.465 94.485 ;
        RECT 260.605 94.470 260.925 94.485 ;
        RECT 262.075 94.470 262.215 94.625 ;
        RECT 262.445 94.625 263.670 94.765 ;
        RECT 262.445 94.565 262.765 94.625 ;
        RECT 263.380 94.580 263.670 94.625 ;
        RECT 264.285 94.765 264.605 94.825 ;
        RECT 281.780 94.765 282.070 94.810 ;
        RECT 287.745 94.765 288.065 94.825 ;
        RECT 264.285 94.625 288.065 94.765 ;
        RECT 264.285 94.565 264.605 94.625 ;
        RECT 281.780 94.580 282.070 94.625 ;
        RECT 287.745 94.565 288.065 94.625 ;
        RECT 288.665 94.765 288.985 94.825 ;
        RECT 294.200 94.765 294.490 94.810 ;
        RECT 288.665 94.625 294.490 94.765 ;
        RECT 296.115 94.765 296.255 94.920 ;
        RECT 298.785 94.905 299.105 95.165 ;
        RECT 299.245 95.105 299.565 95.165 ;
        RECT 307.080 95.105 307.370 95.150 ;
        RECT 308.445 95.105 308.765 95.165 ;
        RECT 299.245 94.965 304.535 95.105 ;
        RECT 299.245 94.905 299.565 94.965 ;
        RECT 297.880 94.765 298.170 94.810 ;
        RECT 296.115 94.625 298.170 94.765 ;
        RECT 298.875 94.765 299.015 94.905 ;
        RECT 300.160 94.765 300.810 94.810 ;
        RECT 303.760 94.765 304.050 94.810 ;
        RECT 298.875 94.625 304.050 94.765 ;
        RECT 304.395 94.765 304.535 94.965 ;
        RECT 307.080 94.965 308.765 95.105 ;
        RECT 307.080 94.920 307.370 94.965 ;
        RECT 308.445 94.905 308.765 94.965 ;
        RECT 308.905 94.905 309.225 95.165 ;
        RECT 304.395 94.625 308.215 94.765 ;
        RECT 288.665 94.565 288.985 94.625 ;
        RECT 294.200 94.580 294.490 94.625 ;
        RECT 297.880 94.580 298.170 94.625 ;
        RECT 300.160 94.580 300.810 94.625 ;
        RECT 303.460 94.580 304.050 94.625 ;
        RECT 260.605 94.240 260.935 94.470 ;
        RECT 262.000 94.240 262.290 94.470 ;
        RECT 260.605 94.225 260.925 94.240 ;
        RECT 262.905 94.225 263.225 94.485 ;
        RECT 263.825 94.225 264.145 94.485 ;
        RECT 278.085 94.225 278.405 94.485 ;
        RECT 278.545 94.425 278.865 94.485 ;
        RECT 279.480 94.425 279.770 94.470 ;
        RECT 283.145 94.425 283.465 94.485 ;
        RECT 284.080 94.425 284.370 94.470 ;
        RECT 278.545 94.285 284.370 94.425 ;
        RECT 278.545 94.225 278.865 94.285 ;
        RECT 279.480 94.240 279.770 94.285 ;
        RECT 283.145 94.225 283.465 94.285 ;
        RECT 284.080 94.240 284.370 94.285 ;
        RECT 284.525 94.425 284.845 94.485 ;
        RECT 285.460 94.425 285.750 94.470 ;
        RECT 284.525 94.285 285.750 94.425 ;
        RECT 284.525 94.225 284.845 94.285 ;
        RECT 285.460 94.240 285.750 94.285 ;
        RECT 286.825 94.425 287.145 94.485 ;
        RECT 293.740 94.425 294.030 94.470 ;
        RECT 286.825 94.285 294.030 94.425 ;
        RECT 286.825 94.225 287.145 94.285 ;
        RECT 293.740 94.240 294.030 94.285 ;
        RECT 242.755 93.945 245.195 94.085 ;
        RECT 247.265 94.085 247.585 94.145 ;
        RECT 264.285 94.085 264.605 94.145 ;
        RECT 247.265 93.945 264.605 94.085 ;
        RECT 247.265 93.885 247.585 93.945 ;
        RECT 264.285 93.885 264.605 93.945 ;
        RECT 276.705 94.085 277.025 94.145 ;
        RECT 279.020 94.085 279.310 94.130 ;
        RECT 276.705 93.945 279.310 94.085 ;
        RECT 276.705 93.885 277.025 93.945 ;
        RECT 279.020 93.900 279.310 93.945 ;
        RECT 278.545 93.745 278.865 93.805 ;
        RECT 228.405 93.605 278.865 93.745 ;
        RECT 279.095 93.745 279.235 93.900 ;
        RECT 282.685 93.885 283.005 94.145 ;
        RECT 286.380 94.085 286.670 94.130 ;
        RECT 293.265 94.085 293.585 94.145 ;
        RECT 286.380 93.945 293.585 94.085 ;
        RECT 286.380 93.900 286.670 93.945 ;
        RECT 293.265 93.885 293.585 93.945 ;
        RECT 280.845 93.745 281.165 93.805 ;
        RECT 282.775 93.745 282.915 93.885 ;
        RECT 279.095 93.605 281.165 93.745 ;
        RECT 228.405 93.545 228.725 93.605 ;
        RECT 278.545 93.545 278.865 93.605 ;
        RECT 280.845 93.545 281.165 93.605 ;
        RECT 282.315 93.605 282.915 93.745 ;
        RECT 210.005 93.405 210.325 93.465 ;
        RECT 206.875 93.265 210.325 93.405 ;
        RECT 210.005 93.205 210.325 93.265 ;
        RECT 211.845 93.205 212.165 93.465 ;
        RECT 224.265 93.205 224.585 93.465 ;
        RECT 230.245 93.205 230.565 93.465 ;
        RECT 243.125 93.405 243.445 93.465 ;
        RECT 244.965 93.405 245.285 93.465 ;
        RECT 243.125 93.265 245.285 93.405 ;
        RECT 243.125 93.205 243.445 93.265 ;
        RECT 244.965 93.205 245.285 93.265 ;
        RECT 247.725 93.205 248.045 93.465 ;
        RECT 261.525 93.205 261.845 93.465 ;
        RECT 264.760 93.405 265.050 93.450 ;
        RECT 275.785 93.405 276.105 93.465 ;
        RECT 264.760 93.265 276.105 93.405 ;
        RECT 264.760 93.220 265.050 93.265 ;
        RECT 275.785 93.205 276.105 93.265 ;
        RECT 277.165 93.405 277.485 93.465 ;
        RECT 282.315 93.405 282.455 93.605 ;
        RECT 277.165 93.265 282.455 93.405 ;
        RECT 284.065 93.405 284.385 93.465 ;
        RECT 284.540 93.405 284.830 93.450 ;
        RECT 284.065 93.265 284.830 93.405 ;
        RECT 294.275 93.405 294.415 94.580 ;
        RECT 296.965 94.425 297.255 94.470 ;
        RECT 298.800 94.425 299.090 94.470 ;
        RECT 302.380 94.425 302.670 94.470 ;
        RECT 296.965 94.285 302.670 94.425 ;
        RECT 296.965 94.240 297.255 94.285 ;
        RECT 298.800 94.240 299.090 94.285 ;
        RECT 302.380 94.240 302.670 94.285 ;
        RECT 303.460 94.265 303.750 94.580 ;
        RECT 306.160 94.425 306.450 94.470 ;
        RECT 307.065 94.425 307.385 94.485 ;
        RECT 308.075 94.470 308.215 94.625 ;
        RECT 306.160 94.285 307.385 94.425 ;
        RECT 306.160 94.240 306.450 94.285 ;
        RECT 307.065 94.225 307.385 94.285 ;
        RECT 308.000 94.240 308.290 94.470 ;
        RECT 295.105 94.085 295.425 94.145 ;
        RECT 296.500 94.085 296.790 94.130 ;
        RECT 305.240 94.085 305.530 94.130 ;
        RECT 295.105 93.945 296.790 94.085 ;
        RECT 295.105 93.885 295.425 93.945 ;
        RECT 296.500 93.900 296.790 93.945 ;
        RECT 297.035 93.945 305.530 94.085 ;
        RECT 297.035 93.405 297.175 93.945 ;
        RECT 305.240 93.900 305.530 93.945 ;
        RECT 297.370 93.745 297.660 93.790 ;
        RECT 299.260 93.745 299.550 93.790 ;
        RECT 302.380 93.745 302.670 93.790 ;
        RECT 297.370 93.605 302.670 93.745 ;
        RECT 297.370 93.560 297.660 93.605 ;
        RECT 299.260 93.560 299.550 93.605 ;
        RECT 302.380 93.560 302.670 93.605 ;
        RECT 294.275 93.265 297.175 93.405 ;
        RECT 298.785 93.405 299.105 93.465 ;
        RECT 300.165 93.405 300.485 93.465 ;
        RECT 301.545 93.405 301.865 93.465 ;
        RECT 298.785 93.265 301.865 93.405 ;
        RECT 277.165 93.205 277.485 93.265 ;
        RECT 284.065 93.205 284.385 93.265 ;
        RECT 284.540 93.220 284.830 93.265 ;
        RECT 298.785 93.205 299.105 93.265 ;
        RECT 300.165 93.205 300.485 93.265 ;
        RECT 301.545 93.205 301.865 93.265 ;
        RECT 302.925 93.405 303.245 93.465 ;
        RECT 303.845 93.405 304.165 93.465 ;
        RECT 302.925 93.265 304.165 93.405 ;
        RECT 302.925 93.205 303.245 93.265 ;
        RECT 303.845 93.205 304.165 93.265 ;
        RECT 162.095 92.585 311.135 93.065 ;
        RECT 203.105 92.385 203.425 92.445 ;
        RECT 173.065 92.245 203.425 92.385 ;
        RECT 173.065 92.045 173.205 92.245 ;
        RECT 203.105 92.185 203.425 92.245 ;
        RECT 203.565 92.385 203.885 92.445 ;
        RECT 212.305 92.385 212.625 92.445 ;
        RECT 203.565 92.245 212.625 92.385 ;
        RECT 203.565 92.185 203.885 92.245 ;
        RECT 212.305 92.185 212.625 92.245 ;
        RECT 226.105 92.385 226.425 92.445 ;
        RECT 228.865 92.385 229.185 92.445 ;
        RECT 233.925 92.385 234.245 92.445 ;
        RECT 244.505 92.385 244.825 92.445 ;
        RECT 246.345 92.385 246.665 92.445 ;
        RECT 258.765 92.385 259.085 92.445 ;
        RECT 260.605 92.385 260.925 92.445 ;
        RECT 226.105 92.245 234.245 92.385 ;
        RECT 226.105 92.185 226.425 92.245 ;
        RECT 228.865 92.185 229.185 92.245 ;
        RECT 233.925 92.185 234.245 92.245 ;
        RECT 234.475 92.245 244.270 92.385 ;
        RECT 227.025 92.045 227.345 92.105 ;
        RECT 171.455 91.905 173.205 92.045 ;
        RECT 206.415 91.905 227.345 92.045 ;
        RECT 165.385 91.705 165.705 91.765 ;
        RECT 171.455 91.750 171.595 91.905 ;
        RECT 171.380 91.705 171.670 91.750 ;
        RECT 165.385 91.565 171.670 91.705 ;
        RECT 165.385 91.505 165.705 91.565 ;
        RECT 171.380 91.520 171.670 91.565 ;
        RECT 178.740 91.705 179.030 91.750 ;
        RECT 183.325 91.705 183.645 91.765 ;
        RECT 206.415 91.705 206.555 91.905 ;
        RECT 227.025 91.845 227.345 91.905 ;
        RECT 229.785 92.045 230.105 92.105 ;
        RECT 233.465 92.045 233.785 92.105 ;
        RECT 229.785 91.905 233.785 92.045 ;
        RECT 229.785 91.845 230.105 91.905 ;
        RECT 233.465 91.845 233.785 91.905 ;
        RECT 178.740 91.565 183.645 91.705 ;
        RECT 178.740 91.520 179.030 91.565 ;
        RECT 183.325 91.505 183.645 91.565 ;
        RECT 196.755 91.565 206.555 91.705 ;
        RECT 206.875 91.565 211.155 91.705 ;
        RECT 182.420 91.365 182.710 91.410 ;
        RECT 193.920 91.365 194.210 91.410 ;
        RECT 194.365 91.365 194.685 91.425 ;
        RECT 173.065 91.225 194.685 91.365 ;
        RECT 165.845 91.025 166.165 91.085 ;
        RECT 173.065 91.025 173.205 91.225 ;
        RECT 182.420 91.180 182.710 91.225 ;
        RECT 193.920 91.180 194.210 91.225 ;
        RECT 194.365 91.165 194.685 91.225 ;
        RECT 195.285 91.165 195.605 91.425 ;
        RECT 196.755 91.410 196.895 91.565 ;
        RECT 196.220 91.180 196.510 91.410 ;
        RECT 196.680 91.180 196.970 91.410 ;
        RECT 197.140 91.365 197.430 91.410 ;
        RECT 198.505 91.365 198.825 91.425 ;
        RECT 197.140 91.225 198.825 91.365 ;
        RECT 197.140 91.180 197.430 91.225 ;
        RECT 177.360 91.025 177.650 91.070 ;
        RECT 179.660 91.025 179.950 91.070 ;
        RECT 165.845 90.885 173.205 91.025 ;
        RECT 173.755 90.885 177.115 91.025 ;
        RECT 165.845 90.825 166.165 90.885 ;
        RECT 173.205 90.685 173.525 90.745 ;
        RECT 173.755 90.685 173.895 90.885 ;
        RECT 173.205 90.545 173.895 90.685 ;
        RECT 174.600 90.685 174.890 90.730 ;
        RECT 175.045 90.685 175.365 90.745 ;
        RECT 174.600 90.545 175.365 90.685 ;
        RECT 173.205 90.485 173.525 90.545 ;
        RECT 174.600 90.500 174.890 90.545 ;
        RECT 175.045 90.485 175.365 90.545 ;
        RECT 175.520 90.685 175.810 90.730 ;
        RECT 176.425 90.685 176.745 90.745 ;
        RECT 175.520 90.545 176.745 90.685 ;
        RECT 176.975 90.685 177.115 90.885 ;
        RECT 177.360 90.885 179.950 91.025 ;
        RECT 177.360 90.840 177.650 90.885 ;
        RECT 179.660 90.840 179.950 90.885 ;
        RECT 192.985 90.825 193.305 91.085 ;
        RECT 194.840 91.025 195.130 91.070 ;
        RECT 196.295 91.025 196.435 91.180 ;
        RECT 198.505 91.165 198.825 91.225 ;
        RECT 203.580 91.180 203.870 91.410 ;
        RECT 206.325 91.365 206.645 91.425 ;
        RECT 206.875 91.365 207.015 91.565 ;
        RECT 206.325 91.225 207.015 91.365 ;
        RECT 207.245 91.365 207.565 91.425 ;
        RECT 208.165 91.365 208.485 91.425 ;
        RECT 207.245 91.225 208.485 91.365 ;
        RECT 203.655 91.025 203.795 91.180 ;
        RECT 206.325 91.165 206.645 91.225 ;
        RECT 207.245 91.165 207.565 91.225 ;
        RECT 208.165 91.165 208.485 91.225 ;
        RECT 208.640 91.180 208.930 91.410 ;
        RECT 194.840 90.885 196.435 91.025 ;
        RECT 196.755 90.885 203.795 91.025 ;
        RECT 208.715 91.025 208.855 91.180 ;
        RECT 210.005 91.165 210.325 91.425 ;
        RECT 211.015 91.410 211.155 91.565 ;
        RECT 211.385 91.505 211.705 91.765 ;
        RECT 211.860 91.705 212.150 91.750 ;
        RECT 212.305 91.705 212.625 91.765 ;
        RECT 229.325 91.705 229.645 91.765 ;
        RECT 234.475 91.705 234.615 92.245 ;
        RECT 243.125 91.845 243.445 92.105 ;
        RECT 244.130 92.045 244.270 92.245 ;
        RECT 244.505 92.245 248.415 92.385 ;
        RECT 244.505 92.185 244.825 92.245 ;
        RECT 246.345 92.185 246.665 92.245 ;
        RECT 244.980 92.045 245.270 92.090 ;
        RECT 244.130 91.905 245.270 92.045 ;
        RECT 244.980 91.860 245.270 91.905 ;
        RECT 211.860 91.565 212.625 91.705 ;
        RECT 211.860 91.520 212.150 91.565 ;
        RECT 212.305 91.505 212.625 91.565 ;
        RECT 228.010 91.565 229.645 91.705 ;
        RECT 210.940 91.180 211.230 91.410 ;
        RECT 212.765 91.165 213.085 91.425 ;
        RECT 213.700 91.365 213.990 91.410 ;
        RECT 216.905 91.365 217.225 91.425 ;
        RECT 228.010 91.410 228.150 91.565 ;
        RECT 229.325 91.505 229.645 91.565 ;
        RECT 230.335 91.565 234.615 91.705 ;
        RECT 243.215 91.705 243.355 91.845 ;
        RECT 244.520 91.705 244.810 91.750 ;
        RECT 247.265 91.705 247.585 91.765 ;
        RECT 243.215 91.565 243.815 91.705 ;
        RECT 213.700 91.225 217.225 91.365 ;
        RECT 213.700 91.180 213.990 91.225 ;
        RECT 216.905 91.165 217.225 91.225 ;
        RECT 227.935 91.180 228.225 91.410 ;
        RECT 228.405 91.165 228.725 91.425 ;
        RECT 229.785 91.365 230.105 91.425 ;
        RECT 230.335 91.410 230.475 91.565 ;
        RECT 229.590 91.225 230.105 91.365 ;
        RECT 229.785 91.165 230.105 91.225 ;
        RECT 230.260 91.180 230.550 91.410 ;
        RECT 231.625 91.165 231.945 91.425 ;
        RECT 232.545 91.165 232.865 91.425 ;
        RECT 233.465 91.165 233.785 91.425 ;
        RECT 242.205 91.165 242.525 91.425 ;
        RECT 242.665 91.165 242.985 91.425 ;
        RECT 243.675 91.410 243.815 91.565 ;
        RECT 244.520 91.565 247.585 91.705 ;
        RECT 244.520 91.520 244.810 91.565 ;
        RECT 246.435 91.410 246.575 91.565 ;
        RECT 247.265 91.505 247.585 91.565 ;
        RECT 248.275 91.425 248.415 92.245 ;
        RECT 258.765 92.245 260.925 92.385 ;
        RECT 258.765 92.185 259.085 92.245 ;
        RECT 260.605 92.185 260.925 92.245 ;
        RECT 261.525 92.385 261.845 92.445 ;
        RECT 267.060 92.385 267.350 92.430 ;
        RECT 261.525 92.245 267.350 92.385 ;
        RECT 261.525 92.185 261.845 92.245 ;
        RECT 267.060 92.200 267.350 92.245 ;
        RECT 267.965 92.385 268.285 92.445 ;
        RECT 269.345 92.385 269.665 92.445 ;
        RECT 281.765 92.385 282.085 92.445 ;
        RECT 267.965 92.245 282.085 92.385 ;
        RECT 267.965 92.185 268.285 92.245 ;
        RECT 269.345 92.185 269.665 92.245 ;
        RECT 281.765 92.185 282.085 92.245 ;
        RECT 301.085 92.385 301.405 92.445 ;
        RECT 308.920 92.385 309.210 92.430 ;
        RECT 301.085 92.245 309.210 92.385 ;
        RECT 301.085 92.185 301.405 92.245 ;
        RECT 308.920 92.200 309.210 92.245 ;
        RECT 256.005 92.045 256.325 92.105 ;
        RECT 262.445 92.045 262.765 92.105 ;
        RECT 256.005 91.905 262.765 92.045 ;
        RECT 256.005 91.845 256.325 91.905 ;
        RECT 243.675 91.225 244.020 91.410 ;
        RECT 243.730 91.180 244.020 91.225 ;
        RECT 245.875 91.180 246.165 91.410 ;
        RECT 246.360 91.180 246.650 91.410 ;
        RECT 247.735 91.365 248.025 91.410 ;
        RECT 247.355 91.225 248.025 91.365 ;
        RECT 224.265 91.025 224.585 91.085 ;
        RECT 208.715 90.885 224.585 91.025 ;
        RECT 194.840 90.840 195.130 90.885 ;
        RECT 177.820 90.685 178.110 90.730 ;
        RECT 178.265 90.685 178.585 90.745 ;
        RECT 176.975 90.545 178.585 90.685 ;
        RECT 175.520 90.500 175.810 90.545 ;
        RECT 176.425 90.485 176.745 90.545 ;
        RECT 177.820 90.500 178.110 90.545 ;
        RECT 178.265 90.485 178.585 90.545 ;
        RECT 185.165 90.685 185.485 90.745 ;
        RECT 196.755 90.685 196.895 90.885 ;
        RECT 224.265 90.825 224.585 90.885 ;
        RECT 225.645 91.025 225.965 91.085 ;
        RECT 225.645 90.885 228.150 91.025 ;
        RECT 225.645 90.825 225.965 90.885 ;
        RECT 185.165 90.545 196.895 90.685 ;
        RECT 185.165 90.485 185.485 90.545 ;
        RECT 198.505 90.485 198.825 90.745 ;
        RECT 204.500 90.685 204.790 90.730 ;
        RECT 205.865 90.685 206.185 90.745 ;
        RECT 204.500 90.545 206.185 90.685 ;
        RECT 204.500 90.500 204.790 90.545 ;
        RECT 205.865 90.485 206.185 90.545 ;
        RECT 206.325 90.685 206.645 90.745 ;
        RECT 207.720 90.685 208.010 90.730 ;
        RECT 206.325 90.545 208.010 90.685 ;
        RECT 206.325 90.485 206.645 90.545 ;
        RECT 207.720 90.500 208.010 90.545 ;
        RECT 209.085 90.685 209.405 90.745 ;
        RECT 209.560 90.685 209.850 90.730 ;
        RECT 209.085 90.545 209.850 90.685 ;
        RECT 209.085 90.485 209.405 90.545 ;
        RECT 209.560 90.500 209.850 90.545 ;
        RECT 215.065 90.685 215.385 90.745 ;
        RECT 227.040 90.685 227.330 90.730 ;
        RECT 215.065 90.545 227.330 90.685 ;
        RECT 228.010 90.685 228.150 90.885 ;
        RECT 228.865 90.825 229.185 91.085 ;
        RECT 231.715 91.025 231.855 91.165 ;
        RECT 229.415 90.885 231.855 91.025 ;
        RECT 229.415 90.685 229.555 90.885 ;
        RECT 232.085 90.825 232.405 91.085 ;
        RECT 243.140 91.025 243.430 91.070 ;
        RECT 245.425 91.025 245.745 91.085 ;
        RECT 243.140 90.885 245.745 91.025 ;
        RECT 243.140 90.840 243.430 90.885 ;
        RECT 245.425 90.825 245.745 90.885 ;
        RECT 228.010 90.545 229.555 90.685 ;
        RECT 215.065 90.485 215.385 90.545 ;
        RECT 227.040 90.500 227.330 90.545 ;
        RECT 230.705 90.485 231.025 90.745 ;
        RECT 231.165 90.685 231.485 90.745 ;
        RECT 241.300 90.685 241.590 90.730 ;
        RECT 231.165 90.545 241.590 90.685 ;
        RECT 231.165 90.485 231.485 90.545 ;
        RECT 241.300 90.500 241.590 90.545 ;
        RECT 241.745 90.685 242.065 90.745 ;
        RECT 245.975 90.685 246.115 91.180 ;
        RECT 247.355 91.085 247.495 91.225 ;
        RECT 247.735 91.180 248.025 91.225 ;
        RECT 248.185 91.165 248.505 91.425 ;
        RECT 260.695 91.410 260.835 91.905 ;
        RECT 262.445 91.845 262.765 91.905 ;
        RECT 263.380 92.045 263.670 92.090 ;
        RECT 282.700 92.045 282.990 92.090 ;
        RECT 263.380 91.905 266.815 92.045 ;
        RECT 263.380 91.860 263.670 91.905 ;
        RECT 262.075 91.565 265.435 91.705 ;
        RECT 262.075 91.410 262.215 91.565 ;
        RECT 265.295 91.425 265.435 91.565 ;
        RECT 260.620 91.180 260.910 91.410 ;
        RECT 262.000 91.180 262.290 91.410 ;
        RECT 262.460 91.180 262.750 91.410 ;
        RECT 246.805 90.825 247.125 91.085 ;
        RECT 247.265 90.825 247.585 91.085 ;
        RECT 259.225 91.025 259.545 91.085 ;
        RECT 261.540 91.025 261.830 91.070 ;
        RECT 259.225 90.885 261.830 91.025 ;
        RECT 259.225 90.825 259.545 90.885 ;
        RECT 261.540 90.840 261.830 90.885 ;
        RECT 249.105 90.685 249.425 90.745 ;
        RECT 241.745 90.545 249.425 90.685 ;
        RECT 241.745 90.485 242.065 90.545 ;
        RECT 249.105 90.485 249.425 90.545 ;
        RECT 250.025 90.685 250.345 90.745 ;
        RECT 262.535 90.685 262.675 91.180 ;
        RECT 263.825 91.165 264.145 91.425 ;
        RECT 265.205 91.165 265.525 91.425 ;
        RECT 265.680 91.180 265.970 91.410 ;
        RECT 266.675 91.365 266.815 91.905 ;
        RECT 270.815 91.905 282.990 92.045 ;
        RECT 267.060 91.365 267.350 91.410 ;
        RECT 266.675 91.225 267.350 91.365 ;
        RECT 267.060 91.180 267.350 91.225 ;
        RECT 264.285 91.025 264.605 91.085 ;
        RECT 264.760 91.025 265.050 91.070 ;
        RECT 264.285 90.885 265.050 91.025 ;
        RECT 265.755 91.025 265.895 91.180 ;
        RECT 267.505 91.165 267.825 91.425 ;
        RECT 268.425 91.025 268.745 91.085 ;
        RECT 270.815 91.025 270.955 91.905 ;
        RECT 282.700 91.860 282.990 91.905 ;
        RECT 284.540 91.860 284.830 92.090 ;
        RECT 278.545 91.705 278.865 91.765 ;
        RECT 278.545 91.565 281.535 91.705 ;
        RECT 278.545 91.505 278.865 91.565 ;
        RECT 278.085 91.365 278.405 91.425 ;
        RECT 279.480 91.365 279.770 91.410 ;
        RECT 278.085 91.225 279.770 91.365 ;
        RECT 281.395 91.365 281.535 91.565 ;
        RECT 281.765 91.505 282.085 91.765 ;
        RECT 282.240 91.705 282.530 91.750 ;
        RECT 283.145 91.705 283.465 91.765 ;
        RECT 282.240 91.565 283.465 91.705 ;
        RECT 284.615 91.705 284.755 91.860 ;
        RECT 290.045 91.845 290.365 92.105 ;
        RECT 295.530 92.045 295.820 92.090 ;
        RECT 297.420 92.045 297.710 92.090 ;
        RECT 300.540 92.045 300.830 92.090 ;
        RECT 295.530 91.905 300.830 92.045 ;
        RECT 295.530 91.860 295.820 91.905 ;
        RECT 297.420 91.860 297.710 91.905 ;
        RECT 300.540 91.860 300.830 91.905 ;
        RECT 302.925 92.045 303.245 92.105 ;
        RECT 303.400 92.045 303.690 92.090 ;
        RECT 302.925 91.905 303.690 92.045 ;
        RECT 302.925 91.845 303.245 91.905 ;
        RECT 303.400 91.860 303.690 91.905 ;
        RECT 287.285 91.705 287.605 91.765 ;
        RECT 293.280 91.705 293.570 91.750 ;
        RECT 307.525 91.705 307.845 91.765 ;
        RECT 284.615 91.565 307.845 91.705 ;
        RECT 282.240 91.520 282.530 91.565 ;
        RECT 283.145 91.505 283.465 91.565 ;
        RECT 287.285 91.505 287.605 91.565 ;
        RECT 293.280 91.520 293.570 91.565 ;
        RECT 307.525 91.505 307.845 91.565 ;
        RECT 283.620 91.365 283.910 91.410 ;
        RECT 284.525 91.365 284.845 91.425 ;
        RECT 291.885 91.365 292.205 91.425 ;
        RECT 281.395 91.225 283.375 91.365 ;
        RECT 278.085 91.165 278.405 91.225 ;
        RECT 279.480 91.180 279.770 91.225 ;
        RECT 265.755 90.885 270.955 91.025 ;
        RECT 277.625 91.025 277.945 91.085 ;
        RECT 280.845 91.070 281.165 91.085 ;
        RECT 279.940 91.025 280.230 91.070 ;
        RECT 277.625 90.885 280.230 91.025 ;
        RECT 264.285 90.825 264.605 90.885 ;
        RECT 264.760 90.840 265.050 90.885 ;
        RECT 268.425 90.825 268.745 90.885 ;
        RECT 277.625 90.825 277.945 90.885 ;
        RECT 279.940 90.840 280.230 90.885 ;
        RECT 280.400 90.840 280.690 91.070 ;
        RECT 280.845 90.840 281.280 91.070 ;
        RECT 283.235 91.025 283.375 91.225 ;
        RECT 283.620 91.225 284.845 91.365 ;
        RECT 283.620 91.180 283.910 91.225 ;
        RECT 284.525 91.165 284.845 91.225 ;
        RECT 290.135 91.225 292.205 91.365 ;
        RECT 290.135 91.025 290.275 91.225 ;
        RECT 291.885 91.165 292.205 91.225 ;
        RECT 292.345 91.165 292.665 91.425 ;
        RECT 294.645 91.165 294.965 91.425 ;
        RECT 295.125 91.365 295.415 91.410 ;
        RECT 296.960 91.365 297.250 91.410 ;
        RECT 300.540 91.365 300.830 91.410 ;
        RECT 295.125 91.225 300.830 91.365 ;
        RECT 295.125 91.180 295.415 91.225 ;
        RECT 296.960 91.180 297.250 91.225 ;
        RECT 300.540 91.180 300.830 91.225 ;
        RECT 301.545 91.385 301.865 91.425 ;
        RECT 301.545 91.165 301.910 91.385 ;
        RECT 303.845 91.365 304.165 91.425 ;
        RECT 306.145 91.365 306.465 91.425 ;
        RECT 308.000 91.365 308.290 91.410 ;
        RECT 303.845 91.225 308.290 91.365 ;
        RECT 303.845 91.165 304.165 91.225 ;
        RECT 306.145 91.165 306.465 91.225 ;
        RECT 308.000 91.180 308.290 91.225 ;
        RECT 283.235 90.885 290.275 91.025 ;
        RECT 290.505 91.025 290.825 91.085 ;
        RECT 301.620 91.070 301.910 91.165 ;
        RECT 296.040 91.025 296.330 91.070 ;
        RECT 290.505 90.885 296.330 91.025 ;
        RECT 265.205 90.685 265.525 90.745 ;
        RECT 250.025 90.545 265.525 90.685 ;
        RECT 250.025 90.485 250.345 90.545 ;
        RECT 265.205 90.485 265.525 90.545 ;
        RECT 266.585 90.485 266.905 90.745 ;
        RECT 268.885 90.485 269.205 90.745 ;
        RECT 276.245 90.685 276.565 90.745 ;
        RECT 278.560 90.685 278.850 90.730 ;
        RECT 276.245 90.545 278.850 90.685 ;
        RECT 280.475 90.685 280.615 90.840 ;
        RECT 280.845 90.825 281.165 90.840 ;
        RECT 290.505 90.825 290.825 90.885 ;
        RECT 296.040 90.840 296.330 90.885 ;
        RECT 298.320 91.025 298.970 91.070 ;
        RECT 301.620 91.025 302.210 91.070 ;
        RECT 298.320 90.885 302.210 91.025 ;
        RECT 298.320 90.840 298.970 90.885 ;
        RECT 301.920 90.840 302.210 90.885 ;
        RECT 302.465 91.025 302.785 91.085 ;
        RECT 304.305 91.025 304.625 91.085 ;
        RECT 302.465 90.885 304.625 91.025 ;
        RECT 302.465 90.825 302.785 90.885 ;
        RECT 304.305 90.825 304.625 90.885 ;
        RECT 282.225 90.685 282.545 90.745 ;
        RECT 280.475 90.545 282.545 90.685 ;
        RECT 276.245 90.485 276.565 90.545 ;
        RECT 278.560 90.500 278.850 90.545 ;
        RECT 282.225 90.485 282.545 90.545 ;
        RECT 291.885 90.485 292.205 90.745 ;
        RECT 292.345 90.685 292.665 90.745 ;
        RECT 302.925 90.685 303.245 90.745 ;
        RECT 292.345 90.545 303.245 90.685 ;
        RECT 292.345 90.485 292.665 90.545 ;
        RECT 302.925 90.485 303.245 90.545 ;
        RECT 162.095 89.865 311.135 90.345 ;
        RECT 165.845 89.665 166.165 89.725 ;
        RECT 169.080 89.665 169.370 89.710 ;
        RECT 165.845 89.525 169.370 89.665 ;
        RECT 165.845 89.465 166.165 89.525 ;
        RECT 169.080 89.480 169.370 89.525 ;
        RECT 175.045 89.665 175.365 89.725 ;
        RECT 180.120 89.665 180.410 89.710 ;
        RECT 175.045 89.525 180.410 89.665 ;
        RECT 175.045 89.465 175.365 89.525 ;
        RECT 180.120 89.480 180.410 89.525 ;
        RECT 186.545 89.665 186.865 89.725 ;
        RECT 204.960 89.665 205.250 89.710 ;
        RECT 206.325 89.665 206.645 89.725 ;
        RECT 186.545 89.525 206.645 89.665 ;
        RECT 186.545 89.465 186.865 89.525 ;
        RECT 204.960 89.480 205.250 89.525 ;
        RECT 206.325 89.465 206.645 89.525 ;
        RECT 207.705 89.665 208.025 89.725 ;
        RECT 229.340 89.665 229.630 89.710 ;
        RECT 207.705 89.525 229.630 89.665 ;
        RECT 207.705 89.465 208.025 89.525 ;
        RECT 229.340 89.480 229.630 89.525 ;
        RECT 243.585 89.665 243.905 89.725 ;
        RECT 246.805 89.665 247.125 89.725 ;
        RECT 243.585 89.525 247.125 89.665 ;
        RECT 243.585 89.465 243.905 89.525 ;
        RECT 246.805 89.465 247.125 89.525 ;
        RECT 249.565 89.665 249.885 89.725 ;
        RECT 258.305 89.665 258.625 89.725 ;
        RECT 249.565 89.525 258.625 89.665 ;
        RECT 249.565 89.465 249.885 89.525 ;
        RECT 258.305 89.465 258.625 89.525 ;
        RECT 263.380 89.665 263.670 89.710 ;
        RECT 267.505 89.665 267.825 89.725 ;
        RECT 263.380 89.525 267.825 89.665 ;
        RECT 263.380 89.480 263.670 89.525 ;
        RECT 267.505 89.465 267.825 89.525 ;
        RECT 277.625 89.465 277.945 89.725 ;
        RECT 286.825 89.665 287.145 89.725 ;
        RECT 288.220 89.665 288.510 89.710 ;
        RECT 286.825 89.525 288.510 89.665 ;
        RECT 286.825 89.465 287.145 89.525 ;
        RECT 288.220 89.480 288.510 89.525 ;
        RECT 290.505 89.465 290.825 89.725 ;
        RECT 303.845 89.465 304.165 89.725 ;
        RECT 174.125 89.370 174.445 89.385 ;
        RECT 170.560 89.325 170.850 89.370 ;
        RECT 173.800 89.325 174.450 89.370 ;
        RECT 170.560 89.185 174.450 89.325 ;
        RECT 170.560 89.140 171.150 89.185 ;
        RECT 173.800 89.140 174.450 89.185 ;
        RECT 170.860 88.825 171.150 89.140 ;
        RECT 174.125 89.125 174.445 89.140 ;
        RECT 176.425 89.125 176.745 89.385 ;
        RECT 176.885 89.325 177.205 89.385 ;
        RECT 180.580 89.325 180.870 89.370 ;
        RECT 187.925 89.325 188.245 89.385 ;
        RECT 176.885 89.185 178.035 89.325 ;
        RECT 176.885 89.125 177.205 89.185 ;
        RECT 177.895 89.030 178.035 89.185 ;
        RECT 180.580 89.185 188.245 89.325 ;
        RECT 180.580 89.140 180.870 89.185 ;
        RECT 187.925 89.125 188.245 89.185 ;
        RECT 188.860 89.325 189.150 89.370 ;
        RECT 195.745 89.325 196.065 89.385 ;
        RECT 188.860 89.185 196.065 89.325 ;
        RECT 188.860 89.140 189.150 89.185 ;
        RECT 171.940 88.985 172.230 89.030 ;
        RECT 175.520 88.985 175.810 89.030 ;
        RECT 177.355 88.985 177.645 89.030 ;
        RECT 171.940 88.845 177.645 88.985 ;
        RECT 171.940 88.800 172.230 88.845 ;
        RECT 175.520 88.800 175.810 88.845 ;
        RECT 177.355 88.800 177.645 88.845 ;
        RECT 177.820 88.800 178.110 89.030 ;
        RECT 178.265 88.985 178.585 89.045 ;
        RECT 188.935 88.985 189.075 89.140 ;
        RECT 195.745 89.125 196.065 89.185 ;
        RECT 203.105 89.125 203.425 89.385 ;
        RECT 204.040 89.325 204.330 89.370 ;
        RECT 215.065 89.325 215.385 89.385 ;
        RECT 250.945 89.325 251.265 89.385 ;
        RECT 204.040 89.185 208.395 89.325 ;
        RECT 204.040 89.140 204.330 89.185 ;
        RECT 178.265 88.845 189.075 88.985 ;
        RECT 178.265 88.785 178.585 88.845 ;
        RECT 189.765 88.785 190.085 89.045 ;
        RECT 192.985 88.985 193.305 89.045 ;
        RECT 194.825 88.985 195.145 89.045 ;
        RECT 202.200 88.985 202.490 89.030 ;
        RECT 203.565 88.985 203.885 89.045 ;
        RECT 192.985 88.845 203.885 88.985 ;
        RECT 192.985 88.785 193.305 88.845 ;
        RECT 194.825 88.785 195.145 88.845 ;
        RECT 202.200 88.800 202.490 88.845 ;
        RECT 203.565 88.785 203.885 88.845 ;
        RECT 204.485 88.785 204.805 89.045 ;
        RECT 205.865 88.785 206.185 89.045 ;
        RECT 208.255 89.030 208.395 89.185 ;
        RECT 208.715 89.185 215.385 89.325 ;
        RECT 208.715 89.030 208.855 89.185 ;
        RECT 215.065 89.125 215.385 89.185 ;
        RECT 216.995 89.185 251.265 89.325 ;
        RECT 207.380 88.985 207.670 89.030 ;
        RECT 207.380 88.800 207.705 88.985 ;
        RECT 208.180 88.800 208.470 89.030 ;
        RECT 208.640 88.800 208.930 89.030 ;
        RECT 181.500 88.645 181.790 88.690 ;
        RECT 183.325 88.645 183.645 88.705 ;
        RECT 181.500 88.505 183.645 88.645 ;
        RECT 181.500 88.460 181.790 88.505 ;
        RECT 183.325 88.445 183.645 88.505 ;
        RECT 190.685 88.445 191.005 88.705 ;
        RECT 171.940 88.305 172.230 88.350 ;
        RECT 175.060 88.305 175.350 88.350 ;
        RECT 176.950 88.305 177.240 88.350 ;
        RECT 171.940 88.165 177.240 88.305 ;
        RECT 205.955 88.305 206.095 88.785 ;
        RECT 206.325 88.645 206.645 88.705 ;
        RECT 207.565 88.645 207.705 88.800 ;
        RECT 209.085 88.785 209.405 89.045 ;
        RECT 211.845 88.985 212.165 89.045 ;
        RECT 216.995 89.030 217.135 89.185 ;
        RECT 250.945 89.125 251.265 89.185 ;
        RECT 259.685 89.325 260.005 89.385 ;
        RECT 262.000 89.325 262.290 89.370 ;
        RECT 270.280 89.325 270.570 89.370 ;
        RECT 298.780 89.325 299.430 89.370 ;
        RECT 300.165 89.325 300.485 89.385 ;
        RECT 302.380 89.325 302.670 89.370 ;
        RECT 259.685 89.185 263.135 89.325 ;
        RECT 259.685 89.125 260.005 89.185 ;
        RECT 262.000 89.140 262.290 89.185 ;
        RECT 215.540 88.985 215.830 89.030 ;
        RECT 211.845 88.845 215.830 88.985 ;
        RECT 211.845 88.785 212.165 88.845 ;
        RECT 215.540 88.800 215.830 88.845 ;
        RECT 216.000 88.800 216.290 89.030 ;
        RECT 216.920 88.800 217.210 89.030 ;
        RECT 217.380 88.985 217.670 89.030 ;
        RECT 225.645 88.985 225.965 89.045 ;
        RECT 217.380 88.845 225.965 88.985 ;
        RECT 217.380 88.800 217.670 88.845 ;
        RECT 210.005 88.645 210.325 88.705 ;
        RECT 206.325 88.505 210.325 88.645 ;
        RECT 206.325 88.445 206.645 88.505 ;
        RECT 210.005 88.445 210.325 88.505 ;
        RECT 216.075 88.645 216.215 88.800 ;
        RECT 225.645 88.785 225.965 88.845 ;
        RECT 230.705 88.785 231.025 89.045 ;
        RECT 231.165 88.785 231.485 89.045 ;
        RECT 242.665 88.785 242.985 89.045 ;
        RECT 243.600 88.800 243.890 89.030 ;
        RECT 238.985 88.645 239.305 88.705 ;
        RECT 243.125 88.645 243.445 88.705 ;
        RECT 216.075 88.505 243.445 88.645 ;
        RECT 243.675 88.645 243.815 88.800 ;
        RECT 244.045 88.785 244.365 89.045 ;
        RECT 244.505 88.985 244.825 89.045 ;
        RECT 244.980 88.985 245.270 89.030 ;
        RECT 244.505 88.845 245.270 88.985 ;
        RECT 244.505 88.785 244.825 88.845 ;
        RECT 244.980 88.800 245.270 88.845 ;
        RECT 245.440 88.985 245.730 89.030 ;
        RECT 247.725 88.985 248.045 89.045 ;
        RECT 245.440 88.845 248.045 88.985 ;
        RECT 245.440 88.800 245.730 88.845 ;
        RECT 247.725 88.785 248.045 88.845 ;
        RECT 250.485 88.985 250.805 89.045 ;
        RECT 260.160 88.985 260.450 89.030 ;
        RECT 250.485 88.845 260.450 88.985 ;
        RECT 250.485 88.785 250.805 88.845 ;
        RECT 260.160 88.800 260.450 88.845 ;
        RECT 260.900 88.985 261.190 89.030 ;
        RECT 260.900 88.800 261.295 88.985 ;
        RECT 243.675 88.505 260.375 88.645 ;
        RECT 216.075 88.305 216.215 88.505 ;
        RECT 238.985 88.445 239.305 88.505 ;
        RECT 243.125 88.445 243.445 88.505 ;
        RECT 260.235 88.365 260.375 88.505 ;
        RECT 205.955 88.165 216.215 88.305 ;
        RECT 234.385 88.305 234.705 88.365 ;
        RECT 252.785 88.305 253.105 88.365 ;
        RECT 234.385 88.165 253.105 88.305 ;
        RECT 171.940 88.120 172.230 88.165 ;
        RECT 175.060 88.120 175.350 88.165 ;
        RECT 176.950 88.120 177.240 88.165 ;
        RECT 234.385 88.105 234.705 88.165 ;
        RECT 252.785 88.105 253.105 88.165 ;
        RECT 260.145 88.105 260.465 88.365 ;
        RECT 261.155 88.305 261.295 88.800 ;
        RECT 261.525 88.785 261.845 89.045 ;
        RECT 262.445 89.030 262.765 89.045 ;
        RECT 262.445 88.985 262.775 89.030 ;
        RECT 262.275 88.845 262.775 88.985 ;
        RECT 262.995 88.985 263.135 89.185 ;
        RECT 270.280 89.185 282.915 89.325 ;
        RECT 270.280 89.140 270.570 89.185 ;
        RECT 263.825 88.985 264.145 89.045 ;
        RECT 262.995 88.845 264.145 88.985 ;
        RECT 262.445 88.800 262.775 88.845 ;
        RECT 262.445 88.785 262.765 88.800 ;
        RECT 263.825 88.785 264.145 88.845 ;
        RECT 275.340 88.800 275.630 89.030 ;
        RECT 266.125 88.445 266.445 88.705 ;
        RECT 266.585 88.645 266.905 88.705 ;
        RECT 275.415 88.645 275.555 88.800 ;
        RECT 276.705 88.785 277.025 89.045 ;
        RECT 279.005 88.785 279.325 89.045 ;
        RECT 282.775 89.030 282.915 89.185 ;
        RECT 298.780 89.185 302.670 89.325 ;
        RECT 298.780 89.140 299.430 89.185 ;
        RECT 300.165 89.125 300.485 89.185 ;
        RECT 302.080 89.140 302.670 89.185 ;
        RECT 282.700 88.985 282.990 89.030 ;
        RECT 285.445 88.985 285.765 89.045 ;
        RECT 282.700 88.845 285.765 88.985 ;
        RECT 282.700 88.800 282.990 88.845 ;
        RECT 285.445 88.785 285.765 88.845 ;
        RECT 288.665 88.985 288.985 89.045 ;
        RECT 292.345 88.985 292.665 89.045 ;
        RECT 288.665 88.845 292.665 88.985 ;
        RECT 288.665 88.785 288.985 88.845 ;
        RECT 292.345 88.785 292.665 88.845 ;
        RECT 295.585 88.985 295.875 89.030 ;
        RECT 297.420 88.985 297.710 89.030 ;
        RECT 301.000 88.985 301.290 89.030 ;
        RECT 295.585 88.845 301.290 88.985 ;
        RECT 295.585 88.800 295.875 88.845 ;
        RECT 297.420 88.800 297.710 88.845 ;
        RECT 301.000 88.800 301.290 88.845 ;
        RECT 302.080 88.825 302.370 89.140 ;
        RECT 302.925 88.985 303.245 89.045 ;
        RECT 305.240 88.985 305.530 89.030 ;
        RECT 302.925 88.845 305.530 88.985 ;
        RECT 302.925 88.785 303.245 88.845 ;
        RECT 305.240 88.800 305.530 88.845 ;
        RECT 266.585 88.505 275.555 88.645 ;
        RECT 266.585 88.445 266.905 88.505 ;
        RECT 275.785 88.445 276.105 88.705 ;
        RECT 287.285 88.445 287.605 88.705 ;
        RECT 295.105 88.445 295.425 88.705 ;
        RECT 296.500 88.645 296.790 88.690 ;
        RECT 304.305 88.645 304.625 88.705 ;
        RECT 296.500 88.505 304.625 88.645 ;
        RECT 296.500 88.460 296.790 88.505 ;
        RECT 304.305 88.445 304.625 88.505 ;
        RECT 267.965 88.305 268.285 88.365 ;
        RECT 291.885 88.305 292.205 88.365 ;
        RECT 261.155 88.165 268.285 88.305 ;
        RECT 267.965 88.105 268.285 88.165 ;
        RECT 275.875 88.165 292.205 88.305 ;
        RECT 173.205 87.965 173.525 88.025 ;
        RECT 178.280 87.965 178.570 88.010 ;
        RECT 173.205 87.825 178.570 87.965 ;
        RECT 173.205 87.765 173.525 87.825 ;
        RECT 178.280 87.780 178.570 87.825 ;
        RECT 195.285 87.965 195.605 88.025 ;
        RECT 199.425 87.965 199.745 88.025 ;
        RECT 206.325 87.965 206.645 88.025 ;
        RECT 195.285 87.825 206.645 87.965 ;
        RECT 195.285 87.765 195.605 87.825 ;
        RECT 199.425 87.765 199.745 87.825 ;
        RECT 206.325 87.765 206.645 87.825 ;
        RECT 206.800 87.965 207.090 88.010 ;
        RECT 207.245 87.965 207.565 88.025 ;
        RECT 206.800 87.825 207.565 87.965 ;
        RECT 206.800 87.780 207.090 87.825 ;
        RECT 207.245 87.765 207.565 87.825 ;
        RECT 210.480 87.965 210.770 88.010 ;
        RECT 210.925 87.965 211.245 88.025 ;
        RECT 210.480 87.825 211.245 87.965 ;
        RECT 210.480 87.780 210.770 87.825 ;
        RECT 210.925 87.765 211.245 87.825 ;
        RECT 211.385 87.965 211.705 88.025 ;
        RECT 218.300 87.965 218.590 88.010 ;
        RECT 211.385 87.825 218.590 87.965 ;
        RECT 211.385 87.765 211.705 87.825 ;
        RECT 218.300 87.780 218.590 87.825 ;
        RECT 230.245 87.765 230.565 88.025 ;
        RECT 232.085 87.965 232.405 88.025 ;
        RECT 275.875 87.965 276.015 88.165 ;
        RECT 291.885 88.105 292.205 88.165 ;
        RECT 295.990 88.305 296.280 88.350 ;
        RECT 297.880 88.305 298.170 88.350 ;
        RECT 301.000 88.305 301.290 88.350 ;
        RECT 295.990 88.165 301.290 88.305 ;
        RECT 295.990 88.120 296.280 88.165 ;
        RECT 297.880 88.120 298.170 88.165 ;
        RECT 301.000 88.120 301.290 88.165 ;
        RECT 232.085 87.825 276.015 87.965 ;
        RECT 232.085 87.765 232.405 87.825 ;
        RECT 276.245 87.765 276.565 88.025 ;
        RECT 300.165 87.965 300.485 88.025 ;
        RECT 305.700 87.965 305.990 88.010 ;
        RECT 300.165 87.825 305.990 87.965 ;
        RECT 300.165 87.765 300.485 87.825 ;
        RECT 305.700 87.780 305.990 87.825 ;
        RECT 162.095 87.145 311.135 87.625 ;
        RECT 165.385 86.945 165.705 87.005 ;
        RECT 165.860 86.945 166.150 86.990 ;
        RECT 165.385 86.805 166.150 86.945 ;
        RECT 165.385 86.745 165.705 86.805 ;
        RECT 165.860 86.760 166.150 86.805 ;
        RECT 168.145 86.945 168.465 87.005 ;
        RECT 168.145 86.805 177.575 86.945 ;
        RECT 168.145 86.745 168.465 86.805 ;
        RECT 168.720 86.605 169.010 86.650 ;
        RECT 171.840 86.605 172.130 86.650 ;
        RECT 173.730 86.605 174.020 86.650 ;
        RECT 168.720 86.465 174.020 86.605 ;
        RECT 168.720 86.420 169.010 86.465 ;
        RECT 171.840 86.420 172.130 86.465 ;
        RECT 173.730 86.420 174.020 86.465 ;
        RECT 173.205 86.065 173.525 86.325 ;
        RECT 174.585 86.065 174.905 86.325 ;
        RECT 177.435 85.970 177.575 86.805 ;
        RECT 186.085 86.745 186.405 87.005 ;
        RECT 212.765 86.945 213.085 87.005 ;
        RECT 186.635 86.805 213.085 86.945 ;
        RECT 178.740 86.265 179.030 86.310 ;
        RECT 182.880 86.265 183.170 86.310 ;
        RECT 183.325 86.265 183.645 86.325 ;
        RECT 178.740 86.125 183.645 86.265 ;
        RECT 178.740 86.080 179.030 86.125 ;
        RECT 182.880 86.080 183.170 86.125 ;
        RECT 183.325 86.065 183.645 86.125 ;
        RECT 167.640 85.630 167.930 85.945 ;
        RECT 168.720 85.925 169.010 85.970 ;
        RECT 172.300 85.925 172.590 85.970 ;
        RECT 174.135 85.925 174.425 85.970 ;
        RECT 168.720 85.785 174.425 85.925 ;
        RECT 168.720 85.740 169.010 85.785 ;
        RECT 172.300 85.740 172.590 85.785 ;
        RECT 174.135 85.740 174.425 85.785 ;
        RECT 177.360 85.925 177.650 85.970 ;
        RECT 186.635 85.925 186.775 86.805 ;
        RECT 212.765 86.745 213.085 86.805 ;
        RECT 245.885 86.945 246.205 87.005 ;
        RECT 245.885 86.805 250.255 86.945 ;
        RECT 245.885 86.745 246.205 86.805 ;
        RECT 187.925 86.605 188.245 86.665 ;
        RECT 188.860 86.605 189.150 86.650 ;
        RECT 242.665 86.605 242.985 86.665 ;
        RECT 187.925 86.465 189.150 86.605 ;
        RECT 187.925 86.405 188.245 86.465 ;
        RECT 188.860 86.420 189.150 86.465 ;
        RECT 197.215 86.465 242.985 86.605 ;
        RECT 193.460 86.265 193.750 86.310 ;
        RECT 193.460 86.125 196.895 86.265 ;
        RECT 193.460 86.080 193.750 86.125 ;
        RECT 177.360 85.785 186.775 85.925 ;
        RECT 177.360 85.740 177.650 85.785 ;
        RECT 187.020 85.740 187.310 85.970 ;
        RECT 167.340 85.585 167.930 85.630 ;
        RECT 170.580 85.585 171.230 85.630 ;
        RECT 171.825 85.585 172.145 85.645 ;
        RECT 167.340 85.445 172.145 85.585 ;
        RECT 167.340 85.400 167.630 85.445 ;
        RECT 170.580 85.400 171.230 85.445 ;
        RECT 171.825 85.385 172.145 85.445 ;
        RECT 175.965 85.585 176.285 85.645 ;
        RECT 177.820 85.585 178.110 85.630 ;
        RECT 175.965 85.445 178.110 85.585 ;
        RECT 175.965 85.385 176.285 85.445 ;
        RECT 177.820 85.400 178.110 85.445 ;
        RECT 181.500 85.585 181.790 85.630 ;
        RECT 183.785 85.585 184.105 85.645 ;
        RECT 181.500 85.445 184.105 85.585 ;
        RECT 187.095 85.585 187.235 85.740 ;
        RECT 187.925 85.725 188.245 85.985 ;
        RECT 189.765 85.725 190.085 85.985 ;
        RECT 190.225 85.725 190.545 85.985 ;
        RECT 194.365 85.725 194.685 85.985 ;
        RECT 195.745 85.725 196.065 85.985 ;
        RECT 196.755 85.970 196.895 86.125 ;
        RECT 197.215 85.970 197.355 86.465 ;
        RECT 242.665 86.405 242.985 86.465 ;
        RECT 244.045 86.605 244.365 86.665 ;
        RECT 250.115 86.605 250.255 86.805 ;
        RECT 250.485 86.745 250.805 87.005 ;
        RECT 270.725 86.945 271.045 87.005 ;
        RECT 255.865 86.805 271.045 86.945 ;
        RECT 255.865 86.605 256.005 86.805 ;
        RECT 270.725 86.745 271.045 86.805 ;
        RECT 276.705 86.945 277.025 87.005 ;
        RECT 281.780 86.945 282.070 86.990 ;
        RECT 276.705 86.805 282.070 86.945 ;
        RECT 276.705 86.745 277.025 86.805 ;
        RECT 281.780 86.760 282.070 86.805 ;
        RECT 291.885 86.945 292.205 87.005 ;
        RECT 296.485 86.945 296.805 87.005 ;
        RECT 297.420 86.945 297.710 86.990 ;
        RECT 291.885 86.805 297.710 86.945 ;
        RECT 291.885 86.745 292.205 86.805 ;
        RECT 296.485 86.745 296.805 86.805 ;
        RECT 297.420 86.760 297.710 86.805 ;
        RECT 304.305 86.745 304.625 87.005 ;
        RECT 244.045 86.465 249.795 86.605 ;
        RECT 250.115 86.465 256.005 86.605 ;
        RECT 260.145 86.605 260.465 86.665 ;
        RECT 276.245 86.605 276.565 86.665 ;
        RECT 260.145 86.465 276.565 86.605 ;
        RECT 244.045 86.405 244.365 86.465 ;
        RECT 198.045 86.265 198.365 86.325 ;
        RECT 204.040 86.265 204.330 86.310 ;
        RECT 249.120 86.265 249.410 86.310 ;
        RECT 198.045 86.125 203.795 86.265 ;
        RECT 198.045 86.065 198.365 86.125 ;
        RECT 196.680 85.740 196.970 85.970 ;
        RECT 197.140 85.740 197.430 85.970 ;
        RECT 197.600 85.925 197.890 85.970 ;
        RECT 200.805 85.925 201.125 85.985 ;
        RECT 197.600 85.785 201.125 85.925 ;
        RECT 197.600 85.740 197.890 85.785 ;
        RECT 200.805 85.725 201.125 85.785 ;
        RECT 203.105 85.725 203.425 85.985 ;
        RECT 203.655 85.925 203.795 86.125 ;
        RECT 204.040 86.125 206.555 86.265 ;
        RECT 204.040 86.080 204.330 86.125 ;
        RECT 205.405 85.925 205.725 85.985 ;
        RECT 206.415 85.970 206.555 86.125 ;
        RECT 242.755 86.125 249.410 86.265 ;
        RECT 242.755 85.985 242.895 86.125 ;
        RECT 249.120 86.080 249.410 86.125 ;
        RECT 249.655 86.265 249.795 86.465 ;
        RECT 260.145 86.405 260.465 86.465 ;
        RECT 276.245 86.405 276.565 86.465 ;
        RECT 289.550 86.605 289.840 86.650 ;
        RECT 291.440 86.605 291.730 86.650 ;
        RECT 294.560 86.605 294.850 86.650 ;
        RECT 289.550 86.465 294.850 86.605 ;
        RECT 289.550 86.420 289.840 86.465 ;
        RECT 291.440 86.420 291.730 86.465 ;
        RECT 294.560 86.420 294.850 86.465 ;
        RECT 250.025 86.265 250.345 86.325 ;
        RECT 249.655 86.125 250.345 86.265 ;
        RECT 203.655 85.785 205.725 85.925 ;
        RECT 205.405 85.725 205.725 85.785 ;
        RECT 206.340 85.740 206.630 85.970 ;
        RECT 206.785 85.725 207.105 85.985 ;
        RECT 207.245 85.725 207.565 85.985 ;
        RECT 211.400 85.925 211.690 85.970 ;
        RECT 212.765 85.925 213.085 85.985 ;
        RECT 211.400 85.785 213.085 85.925 ;
        RECT 211.400 85.740 211.690 85.785 ;
        RECT 212.765 85.725 213.085 85.785 ;
        RECT 223.345 85.925 223.665 85.985 ;
        RECT 242.665 85.925 242.985 85.985 ;
        RECT 223.345 85.785 242.985 85.925 ;
        RECT 223.345 85.725 223.665 85.785 ;
        RECT 242.665 85.725 242.985 85.785 ;
        RECT 243.125 85.925 243.445 85.985 ;
        RECT 243.600 85.925 243.890 85.970 ;
        RECT 243.125 85.785 243.890 85.925 ;
        RECT 243.125 85.725 243.445 85.785 ;
        RECT 243.600 85.740 243.890 85.785 ;
        RECT 244.045 85.925 244.365 85.985 ;
        RECT 244.520 85.925 244.810 85.970 ;
        RECT 244.045 85.785 244.810 85.925 ;
        RECT 189.855 85.585 189.995 85.725 ;
        RECT 187.095 85.445 189.995 85.585 ;
        RECT 195.300 85.585 195.590 85.630 ;
        RECT 202.185 85.585 202.505 85.645 ;
        RECT 195.300 85.445 202.505 85.585 ;
        RECT 205.495 85.585 205.635 85.725 ;
        RECT 210.005 85.585 210.325 85.645 ;
        RECT 210.480 85.585 210.770 85.630 ;
        RECT 217.365 85.585 217.685 85.645 ;
        RECT 205.495 85.445 209.775 85.585 ;
        RECT 181.500 85.400 181.790 85.445 ;
        RECT 183.785 85.385 184.105 85.445 ;
        RECT 195.300 85.400 195.590 85.445 ;
        RECT 202.185 85.385 202.505 85.445 ;
        RECT 175.505 85.045 175.825 85.305 ;
        RECT 179.645 85.045 179.965 85.305 ;
        RECT 181.960 85.245 182.250 85.290 ;
        RECT 186.085 85.245 186.405 85.305 ;
        RECT 181.960 85.105 186.405 85.245 ;
        RECT 181.960 85.060 182.250 85.105 ;
        RECT 186.085 85.045 186.405 85.105 ;
        RECT 195.745 85.245 196.065 85.305 ;
        RECT 198.045 85.245 198.365 85.305 ;
        RECT 195.745 85.105 198.365 85.245 ;
        RECT 195.745 85.045 196.065 85.105 ;
        RECT 198.045 85.045 198.365 85.105 ;
        RECT 198.965 85.045 199.285 85.305 ;
        RECT 208.640 85.245 208.930 85.290 ;
        RECT 209.085 85.245 209.405 85.305 ;
        RECT 208.640 85.105 209.405 85.245 ;
        RECT 209.635 85.245 209.775 85.445 ;
        RECT 210.005 85.445 210.770 85.585 ;
        RECT 210.005 85.385 210.325 85.445 ;
        RECT 210.480 85.400 210.770 85.445 ;
        RECT 211.935 85.445 217.685 85.585 ;
        RECT 211.935 85.245 212.075 85.445 ;
        RECT 217.365 85.385 217.685 85.445 ;
        RECT 224.725 85.585 225.045 85.645 ;
        RECT 229.325 85.585 229.645 85.645 ;
        RECT 224.725 85.445 229.645 85.585 ;
        RECT 243.675 85.585 243.815 85.740 ;
        RECT 244.045 85.725 244.365 85.785 ;
        RECT 244.520 85.740 244.810 85.785 ;
        RECT 245.440 85.925 245.730 85.970 ;
        RECT 247.280 85.925 247.570 85.970 ;
        RECT 245.440 85.785 247.570 85.925 ;
        RECT 245.440 85.740 245.730 85.785 ;
        RECT 247.280 85.740 247.570 85.785 ;
        RECT 248.660 85.925 248.950 85.970 ;
        RECT 249.655 85.925 249.795 86.125 ;
        RECT 250.025 86.065 250.345 86.125 ;
        RECT 256.005 86.265 256.325 86.325 ;
        RECT 262.445 86.265 262.765 86.325 ;
        RECT 281.765 86.265 282.085 86.325 ;
        RECT 295.105 86.265 295.425 86.325 ;
        RECT 256.005 86.125 262.765 86.265 ;
        RECT 256.005 86.065 256.325 86.125 ;
        RECT 262.445 86.065 262.765 86.125 ;
        RECT 264.835 86.125 282.085 86.265 ;
        RECT 264.835 85.985 264.975 86.125 ;
        RECT 281.765 86.065 282.085 86.125 ;
        RECT 288.755 86.125 295.425 86.265 ;
        RECT 248.660 85.785 249.795 85.925 ;
        RECT 256.925 85.925 257.245 85.985 ;
        RECT 264.745 85.925 265.065 85.985 ;
        RECT 256.925 85.785 265.065 85.925 ;
        RECT 248.660 85.740 248.950 85.785 ;
        RECT 245.515 85.585 245.655 85.740 ;
        RECT 243.675 85.445 245.655 85.585 ;
        RECT 224.725 85.385 225.045 85.445 ;
        RECT 229.325 85.385 229.645 85.445 ;
        RECT 209.635 85.105 212.075 85.245 ;
        RECT 208.640 85.060 208.930 85.105 ;
        RECT 209.085 85.045 209.405 85.105 ;
        RECT 212.305 85.045 212.625 85.305 ;
        RECT 228.865 85.245 229.185 85.305 ;
        RECT 229.785 85.245 230.105 85.305 ;
        RECT 228.865 85.105 230.105 85.245 ;
        RECT 228.865 85.045 229.185 85.105 ;
        RECT 229.785 85.045 230.105 85.105 ;
        RECT 240.825 85.245 241.145 85.305 ;
        RECT 242.680 85.245 242.970 85.290 ;
        RECT 240.825 85.105 242.970 85.245 ;
        RECT 240.825 85.045 241.145 85.105 ;
        RECT 242.680 85.060 242.970 85.105 ;
        RECT 244.045 85.245 244.365 85.305 ;
        RECT 244.520 85.245 244.810 85.290 ;
        RECT 246.805 85.245 247.125 85.305 ;
        RECT 244.045 85.105 247.125 85.245 ;
        RECT 247.355 85.245 247.495 85.740 ;
        RECT 256.925 85.725 257.245 85.785 ;
        RECT 264.745 85.725 265.065 85.785 ;
        RECT 266.125 85.725 266.445 85.985 ;
        RECT 278.560 85.925 278.850 85.970 ;
        RECT 279.005 85.925 279.325 85.985 ;
        RECT 278.560 85.785 279.325 85.925 ;
        RECT 278.560 85.740 278.850 85.785 ;
        RECT 279.005 85.725 279.325 85.785 ;
        RECT 282.700 85.740 282.990 85.970 ;
        RECT 284.065 85.925 284.385 85.985 ;
        RECT 283.870 85.785 284.385 85.925 ;
        RECT 249.705 85.585 249.995 85.630 ;
        RECT 270.265 85.585 270.585 85.645 ;
        RECT 282.775 85.585 282.915 85.740 ;
        RECT 284.065 85.725 284.385 85.785 ;
        RECT 286.365 85.925 286.685 85.985 ;
        RECT 288.755 85.970 288.895 86.125 ;
        RECT 295.105 86.065 295.425 86.125 ;
        RECT 296.025 86.265 296.345 86.325 ;
        RECT 300.640 86.265 300.930 86.310 ;
        RECT 296.025 86.125 300.930 86.265 ;
        RECT 296.025 86.065 296.345 86.125 ;
        RECT 300.640 86.080 300.930 86.125 ;
        RECT 304.765 86.265 305.085 86.325 ;
        RECT 306.620 86.265 306.910 86.310 ;
        RECT 304.765 86.125 306.910 86.265 ;
        RECT 304.765 86.065 305.085 86.125 ;
        RECT 306.620 86.080 306.910 86.125 ;
        RECT 307.525 86.065 307.845 86.325 ;
        RECT 288.680 85.925 288.970 85.970 ;
        RECT 286.365 85.785 288.970 85.925 ;
        RECT 286.365 85.725 286.685 85.785 ;
        RECT 288.680 85.740 288.970 85.785 ;
        RECT 289.145 85.925 289.435 85.970 ;
        RECT 290.980 85.925 291.270 85.970 ;
        RECT 294.560 85.925 294.850 85.970 ;
        RECT 289.145 85.785 294.850 85.925 ;
        RECT 289.145 85.740 289.435 85.785 ;
        RECT 290.980 85.740 291.270 85.785 ;
        RECT 294.560 85.740 294.850 85.785 ;
        RECT 295.640 85.925 295.930 85.945 ;
        RECT 300.165 85.925 300.485 85.985 ;
        RECT 295.640 85.785 300.485 85.925 ;
        RECT 249.705 85.445 269.805 85.585 ;
        RECT 249.705 85.400 249.995 85.445 ;
        RECT 248.645 85.245 248.965 85.305 ;
        RECT 247.355 85.105 248.965 85.245 ;
        RECT 244.045 85.045 244.365 85.105 ;
        RECT 244.520 85.060 244.810 85.105 ;
        RECT 246.805 85.045 247.125 85.105 ;
        RECT 248.645 85.045 248.965 85.105 ;
        RECT 249.105 85.245 249.425 85.305 ;
        RECT 261.525 85.245 261.845 85.305 ;
        RECT 266.585 85.245 266.905 85.305 ;
        RECT 249.105 85.105 266.905 85.245 ;
        RECT 269.665 85.245 269.805 85.445 ;
        RECT 270.265 85.445 282.915 85.585 ;
        RECT 270.265 85.385 270.585 85.445 ;
        RECT 290.045 85.385 290.365 85.645 ;
        RECT 295.640 85.630 295.930 85.785 ;
        RECT 300.165 85.725 300.485 85.785 ;
        RECT 306.145 85.725 306.465 85.985 ;
        RECT 309.365 85.725 309.685 85.985 ;
        RECT 292.340 85.585 292.990 85.630 ;
        RECT 295.640 85.585 296.230 85.630 ;
        RECT 292.340 85.445 296.230 85.585 ;
        RECT 292.340 85.400 292.990 85.445 ;
        RECT 295.940 85.400 296.230 85.445 ;
        RECT 296.945 85.585 297.265 85.645 ;
        RECT 299.720 85.585 300.010 85.630 ;
        RECT 296.945 85.445 300.010 85.585 ;
        RECT 296.945 85.385 297.265 85.445 ;
        RECT 299.720 85.400 300.010 85.445 ;
        RECT 283.620 85.245 283.910 85.290 ;
        RECT 288.205 85.245 288.525 85.305 ;
        RECT 269.665 85.105 288.525 85.245 ;
        RECT 249.105 85.045 249.425 85.105 ;
        RECT 261.525 85.045 261.845 85.105 ;
        RECT 266.585 85.045 266.905 85.105 ;
        RECT 283.620 85.060 283.910 85.105 ;
        RECT 288.205 85.045 288.525 85.105 ;
        RECT 297.865 85.045 298.185 85.305 ;
        RECT 300.165 85.045 300.485 85.305 ;
        RECT 307.525 85.245 307.845 85.305 ;
        RECT 308.460 85.245 308.750 85.290 ;
        RECT 307.525 85.105 308.750 85.245 ;
        RECT 307.525 85.045 307.845 85.105 ;
        RECT 308.460 85.060 308.750 85.105 ;
        RECT 162.095 84.425 311.135 84.905 ;
        RECT 168.605 84.225 168.925 84.285 ;
        RECT 170.920 84.225 171.210 84.270 ;
        RECT 168.605 84.085 171.210 84.225 ;
        RECT 168.605 84.025 168.925 84.085 ;
        RECT 170.920 84.040 171.210 84.085 ;
        RECT 171.825 84.225 172.145 84.285 ;
        RECT 174.125 84.225 174.445 84.285 ;
        RECT 171.825 84.085 174.445 84.225 ;
        RECT 171.825 84.025 172.145 84.085 ;
        RECT 174.125 84.025 174.445 84.085 ;
        RECT 174.585 84.225 174.905 84.285 ;
        RECT 174.585 84.085 179.875 84.225 ;
        RECT 174.585 84.025 174.905 84.085 ;
        RECT 171.915 83.885 172.055 84.025 ;
        RECT 172.400 83.885 172.690 83.930 ;
        RECT 175.640 83.885 176.290 83.930 ;
        RECT 171.915 83.745 176.290 83.885 ;
        RECT 172.400 83.700 172.990 83.745 ;
        RECT 175.640 83.700 176.290 83.745 ;
        RECT 172.700 83.385 172.990 83.700 ;
        RECT 179.735 83.590 179.875 84.085 ;
        RECT 183.325 84.025 183.645 84.285 ;
        RECT 183.785 84.225 184.105 84.285 ;
        RECT 231.625 84.225 231.945 84.285 ;
        RECT 234.845 84.225 235.165 84.285 ;
        RECT 183.785 84.085 215.755 84.225 ;
        RECT 183.785 84.025 184.105 84.085 ;
        RECT 192.985 83.885 193.305 83.945 ;
        RECT 185.715 83.745 193.305 83.885 ;
        RECT 185.715 83.605 185.855 83.745 ;
        RECT 192.985 83.685 193.305 83.745 ;
        RECT 206.800 83.885 207.090 83.930 ;
        RECT 210.465 83.885 210.785 83.945 ;
        RECT 212.305 83.885 212.625 83.945 ;
        RECT 206.800 83.745 210.785 83.885 ;
        RECT 206.800 83.700 207.090 83.745 ;
        RECT 210.465 83.685 210.785 83.745 ;
        RECT 211.015 83.745 212.625 83.885 ;
        RECT 173.780 83.545 174.070 83.590 ;
        RECT 177.360 83.545 177.650 83.590 ;
        RECT 179.195 83.545 179.485 83.590 ;
        RECT 173.780 83.405 179.485 83.545 ;
        RECT 173.780 83.360 174.070 83.405 ;
        RECT 177.360 83.360 177.650 83.405 ;
        RECT 179.195 83.360 179.485 83.405 ;
        RECT 179.660 83.360 179.950 83.590 ;
        RECT 184.260 83.360 184.550 83.590 ;
        RECT 175.505 83.205 175.825 83.265 ;
        RECT 178.280 83.205 178.570 83.250 ;
        RECT 175.505 83.065 178.570 83.205 ;
        RECT 184.335 83.205 184.475 83.360 ;
        RECT 185.165 83.345 185.485 83.605 ;
        RECT 185.625 83.345 185.945 83.605 ;
        RECT 189.765 83.345 190.085 83.605 ;
        RECT 205.405 83.545 205.725 83.605 ;
        RECT 211.015 83.590 211.155 83.745 ;
        RECT 212.305 83.685 212.625 83.745 ;
        RECT 215.615 83.885 215.755 84.085 ;
        RECT 227.115 84.085 235.165 84.225 ;
        RECT 220.125 83.885 220.445 83.945 ;
        RECT 215.615 83.745 220.445 83.885 ;
        RECT 210.020 83.545 210.310 83.590 ;
        RECT 205.405 83.405 210.310 83.545 ;
        RECT 205.405 83.345 205.725 83.405 ;
        RECT 210.020 83.360 210.310 83.405 ;
        RECT 210.940 83.360 211.230 83.590 ;
        RECT 211.385 83.345 211.705 83.605 ;
        RECT 211.845 83.345 212.165 83.605 ;
        RECT 215.615 83.590 215.755 83.745 ;
        RECT 220.125 83.685 220.445 83.745 ;
        RECT 215.540 83.360 215.830 83.590 ;
        RECT 216.000 83.360 216.290 83.590 ;
        RECT 216.460 83.360 216.750 83.590 ;
        RECT 187.005 83.205 187.325 83.265 ;
        RECT 184.335 83.065 187.325 83.205 ;
        RECT 175.505 83.005 175.825 83.065 ;
        RECT 178.280 83.020 178.570 83.065 ;
        RECT 187.005 83.005 187.325 83.065 ;
        RECT 187.465 83.205 187.785 83.265 ;
        RECT 190.700 83.205 190.990 83.250 ;
        RECT 187.465 83.065 190.990 83.205 ;
        RECT 187.465 83.005 187.785 83.065 ;
        RECT 190.700 83.020 190.990 83.065 ;
        RECT 202.185 83.205 202.505 83.265 ;
        RECT 216.075 83.205 216.215 83.360 ;
        RECT 202.185 83.065 216.215 83.205 ;
        RECT 216.535 83.205 216.675 83.360 ;
        RECT 217.365 83.345 217.685 83.605 ;
        RECT 226.565 83.545 226.885 83.605 ;
        RECT 227.115 83.590 227.255 84.085 ;
        RECT 231.625 84.025 231.945 84.085 ;
        RECT 234.845 84.025 235.165 84.085 ;
        RECT 241.745 84.025 242.065 84.285 ;
        RECT 245.885 84.225 246.205 84.285 ;
        RECT 245.510 84.085 246.205 84.225 ;
        RECT 227.485 83.885 227.805 83.945 ;
        RECT 240.825 83.885 241.145 83.945 ;
        RECT 227.485 83.745 241.145 83.885 ;
        RECT 241.835 83.885 241.975 84.025 ;
        RECT 244.060 83.885 244.350 83.930 ;
        RECT 244.965 83.885 245.285 83.945 ;
        RECT 241.835 83.745 243.355 83.885 ;
        RECT 227.485 83.685 227.805 83.745 ;
        RECT 240.825 83.685 241.145 83.745 ;
        RECT 221.365 83.405 226.885 83.545 ;
        RECT 221.365 83.205 221.505 83.405 ;
        RECT 226.565 83.345 226.885 83.405 ;
        RECT 227.040 83.360 227.330 83.590 ;
        RECT 227.945 83.545 228.265 83.605 ;
        RECT 227.575 83.405 228.265 83.545 ;
        RECT 216.535 83.065 221.505 83.205 ;
        RECT 202.185 83.005 202.505 83.065 ;
        RECT 173.780 82.865 174.070 82.910 ;
        RECT 176.900 82.865 177.190 82.910 ;
        RECT 178.790 82.865 179.080 82.910 ;
        RECT 173.780 82.725 179.080 82.865 ;
        RECT 187.095 82.865 187.235 83.005 ;
        RECT 188.385 82.865 188.705 82.925 ;
        RECT 187.095 82.725 188.705 82.865 ;
        RECT 173.780 82.680 174.070 82.725 ;
        RECT 176.900 82.680 177.190 82.725 ;
        RECT 178.790 82.680 179.080 82.725 ;
        RECT 188.385 82.665 188.705 82.725 ;
        RECT 190.225 82.865 190.545 82.925 ;
        RECT 204.485 82.865 204.805 82.925 ;
        RECT 190.225 82.725 204.805 82.865 ;
        RECT 190.225 82.665 190.545 82.725 ;
        RECT 204.485 82.665 204.805 82.725 ;
        RECT 213.240 82.865 213.530 82.910 ;
        RECT 215.525 82.865 215.845 82.925 ;
        RECT 213.240 82.725 215.845 82.865 ;
        RECT 213.240 82.680 213.530 82.725 ;
        RECT 215.525 82.665 215.845 82.725 ;
        RECT 175.965 82.525 176.285 82.585 ;
        RECT 188.860 82.525 189.150 82.570 ;
        RECT 175.965 82.385 189.150 82.525 ;
        RECT 175.965 82.325 176.285 82.385 ;
        RECT 188.860 82.340 189.150 82.385 ;
        RECT 190.685 82.525 191.005 82.585 ;
        RECT 203.105 82.525 203.425 82.585 ;
        RECT 190.685 82.385 203.425 82.525 ;
        RECT 190.685 82.325 191.005 82.385 ;
        RECT 203.105 82.325 203.425 82.385 ;
        RECT 207.705 82.525 208.025 82.585 ;
        RECT 209.545 82.525 209.865 82.585 ;
        RECT 207.705 82.385 209.865 82.525 ;
        RECT 207.705 82.325 208.025 82.385 ;
        RECT 209.545 82.325 209.865 82.385 ;
        RECT 214.160 82.525 214.450 82.570 ;
        RECT 214.605 82.525 214.925 82.585 ;
        RECT 214.160 82.385 214.925 82.525 ;
        RECT 214.160 82.340 214.450 82.385 ;
        RECT 214.605 82.325 214.925 82.385 ;
        RECT 215.985 82.525 216.305 82.585 ;
        RECT 227.575 82.525 227.715 83.405 ;
        RECT 227.945 83.345 228.265 83.405 ;
        RECT 228.405 83.345 228.725 83.605 ;
        RECT 228.880 83.545 229.170 83.590 ;
        RECT 229.325 83.545 229.645 83.605 ;
        RECT 239.445 83.545 239.765 83.605 ;
        RECT 228.880 83.405 239.765 83.545 ;
        RECT 228.880 83.360 229.170 83.405 ;
        RECT 229.325 83.345 229.645 83.405 ;
        RECT 239.445 83.345 239.765 83.405 ;
        RECT 241.760 83.360 242.050 83.590 ;
        RECT 242.220 83.545 242.510 83.590 ;
        RECT 242.665 83.545 242.985 83.605 ;
        RECT 242.220 83.405 242.985 83.545 ;
        RECT 243.215 83.545 243.355 83.745 ;
        RECT 244.060 83.745 245.285 83.885 ;
        RECT 244.060 83.700 244.350 83.745 ;
        RECT 244.965 83.685 245.285 83.745 ;
        RECT 245.510 83.590 245.650 84.085 ;
        RECT 245.885 84.025 246.205 84.085 ;
        RECT 246.345 84.225 246.665 84.285 ;
        RECT 248.185 84.225 248.505 84.285 ;
        RECT 252.340 84.225 252.630 84.270 ;
        RECT 246.345 84.085 252.630 84.225 ;
        RECT 246.345 84.025 246.665 84.085 ;
        RECT 248.185 84.025 248.505 84.085 ;
        RECT 252.340 84.040 252.630 84.085 ;
        RECT 254.625 84.225 254.945 84.285 ;
        RECT 264.300 84.225 264.590 84.270 ;
        RECT 254.625 84.085 264.590 84.225 ;
        RECT 254.625 84.025 254.945 84.085 ;
        RECT 264.300 84.040 264.590 84.085 ;
        RECT 297.865 84.025 298.185 84.285 ;
        RECT 247.695 83.885 247.985 83.930 ;
        RECT 248.645 83.885 248.965 83.945 ;
        RECT 256.465 83.885 256.785 83.945 ;
        RECT 247.695 83.745 248.965 83.885 ;
        RECT 247.695 83.700 247.985 83.745 ;
        RECT 248.645 83.685 248.965 83.745 ;
        RECT 255.865 83.745 256.785 83.885 ;
        RECT 243.575 83.545 243.865 83.590 ;
        RECT 243.215 83.405 243.865 83.545 ;
        RECT 242.220 83.360 242.510 83.405 ;
        RECT 241.835 83.205 241.975 83.360 ;
        RECT 242.665 83.345 242.985 83.405 ;
        RECT 243.575 83.360 243.865 83.405 ;
        RECT 244.520 83.360 244.810 83.590 ;
        RECT 245.435 83.360 245.725 83.590 ;
        RECT 244.045 83.205 244.365 83.265 ;
        RECT 244.595 83.205 244.735 83.360 ;
        RECT 228.495 83.065 243.790 83.205 ;
        RECT 228.495 82.925 228.635 83.065 ;
        RECT 228.405 82.665 228.725 82.925 ;
        RECT 231.165 82.865 231.485 82.925 ;
        RECT 229.415 82.725 231.485 82.865 ;
        RECT 215.985 82.385 227.715 82.525 ;
        RECT 227.945 82.525 228.265 82.585 ;
        RECT 229.415 82.525 229.555 82.725 ;
        RECT 231.165 82.665 231.485 82.725 ;
        RECT 241.745 82.865 242.065 82.925 ;
        RECT 242.220 82.865 242.510 82.910 ;
        RECT 241.745 82.725 242.510 82.865 ;
        RECT 243.650 82.865 243.790 83.065 ;
        RECT 244.045 83.065 244.735 83.205 ;
        RECT 244.965 83.205 245.285 83.265 ;
        RECT 245.510 83.205 245.650 83.360 ;
        RECT 245.885 83.345 246.205 83.605 ;
        RECT 246.805 83.545 247.125 83.605 ;
        RECT 249.580 83.545 249.870 83.590 ;
        RECT 246.805 83.405 249.870 83.545 ;
        RECT 246.805 83.345 247.125 83.405 ;
        RECT 249.580 83.360 249.870 83.405 ;
        RECT 244.965 83.065 245.650 83.205 ;
        RECT 244.045 83.005 244.365 83.065 ;
        RECT 244.965 83.005 245.285 83.065 ;
        RECT 246.345 82.865 246.665 82.925 ;
        RECT 243.650 82.725 246.665 82.865 ;
        RECT 241.745 82.665 242.065 82.725 ;
        RECT 242.220 82.680 242.510 82.725 ;
        RECT 246.345 82.665 246.665 82.725 ;
        RECT 246.820 82.865 247.110 82.910 ;
        RECT 249.105 82.865 249.425 82.925 ;
        RECT 246.820 82.725 249.425 82.865 ;
        RECT 249.655 82.865 249.795 83.360 ;
        RECT 250.025 83.345 250.345 83.605 ;
        RECT 252.785 83.545 253.105 83.605 ;
        RECT 255.865 83.545 256.005 83.745 ;
        RECT 256.465 83.685 256.785 83.745 ;
        RECT 259.685 83.685 260.005 83.945 ;
        RECT 260.160 83.885 260.450 83.930 ;
        RECT 271.645 83.885 271.965 83.945 ;
        RECT 283.605 83.885 283.925 83.945 ;
        RECT 260.160 83.745 283.925 83.885 ;
        RECT 260.160 83.700 260.450 83.745 ;
        RECT 271.645 83.685 271.965 83.745 ;
        RECT 283.605 83.685 283.925 83.745 ;
        RECT 296.040 83.885 296.330 83.930 ;
        RECT 297.955 83.885 298.095 84.025 ;
        RECT 296.040 83.745 298.095 83.885 ;
        RECT 298.320 83.885 298.970 83.930 ;
        RECT 301.920 83.885 302.210 83.930 ;
        RECT 302.925 83.885 303.245 83.945 ;
        RECT 298.320 83.745 303.245 83.885 ;
        RECT 296.040 83.700 296.330 83.745 ;
        RECT 298.320 83.700 298.970 83.745 ;
        RECT 301.620 83.700 302.210 83.745 ;
        RECT 252.785 83.405 256.005 83.545 ;
        RECT 258.780 83.545 259.070 83.590 ;
        RECT 259.225 83.545 259.545 83.605 ;
        RECT 258.780 83.405 259.545 83.545 ;
        RECT 252.785 83.345 253.105 83.405 ;
        RECT 258.780 83.360 259.070 83.405 ;
        RECT 259.225 83.345 259.545 83.405 ;
        RECT 255.085 83.205 255.405 83.265 ;
        RECT 259.775 83.205 259.915 83.685 ;
        RECT 260.620 83.360 260.910 83.590 ;
        RECT 261.065 83.545 261.385 83.605 ;
        RECT 262.000 83.545 262.290 83.590 ;
        RECT 261.065 83.405 262.290 83.545 ;
        RECT 255.085 83.065 259.915 83.205 ;
        RECT 260.695 83.205 260.835 83.360 ;
        RECT 261.065 83.345 261.385 83.405 ;
        RECT 262.000 83.360 262.290 83.405 ;
        RECT 263.380 83.545 263.670 83.590 ;
        RECT 265.680 83.545 265.970 83.590 ;
        RECT 263.380 83.405 265.970 83.545 ;
        RECT 263.380 83.360 263.670 83.405 ;
        RECT 265.680 83.360 265.970 83.405 ;
        RECT 266.585 83.345 266.905 83.605 ;
        RECT 286.365 83.545 286.685 83.605 ;
        RECT 287.760 83.545 288.050 83.590 ;
        RECT 286.365 83.405 288.050 83.545 ;
        RECT 286.365 83.345 286.685 83.405 ;
        RECT 287.760 83.360 288.050 83.405 ;
        RECT 295.125 83.545 295.415 83.590 ;
        RECT 296.960 83.545 297.250 83.590 ;
        RECT 300.540 83.545 300.830 83.590 ;
        RECT 295.125 83.405 300.830 83.545 ;
        RECT 295.125 83.360 295.415 83.405 ;
        RECT 296.960 83.360 297.250 83.405 ;
        RECT 300.540 83.360 300.830 83.405 ;
        RECT 301.620 83.385 301.910 83.700 ;
        RECT 302.925 83.685 303.245 83.745 ;
        RECT 304.765 83.885 305.085 83.945 ;
        RECT 305.700 83.885 305.990 83.930 ;
        RECT 306.605 83.885 306.925 83.945 ;
        RECT 304.765 83.745 306.925 83.885 ;
        RECT 304.765 83.685 305.085 83.745 ;
        RECT 305.700 83.700 305.990 83.745 ;
        RECT 306.605 83.685 306.925 83.745 ;
        RECT 260.695 83.065 261.755 83.205 ;
        RECT 255.085 83.005 255.405 83.065 ;
        RECT 250.960 82.865 251.250 82.910 ;
        RECT 249.655 82.725 251.250 82.865 ;
        RECT 246.820 82.680 247.110 82.725 ;
        RECT 249.105 82.665 249.425 82.725 ;
        RECT 250.960 82.680 251.250 82.725 ;
        RECT 253.245 82.865 253.565 82.925 ;
        RECT 260.695 82.865 260.835 83.065 ;
        RECT 253.245 82.725 260.835 82.865 ;
        RECT 261.615 82.865 261.755 83.065 ;
        RECT 262.905 83.005 263.225 83.265 ;
        RECT 267.505 83.005 267.825 83.265 ;
        RECT 294.185 83.205 294.505 83.265 ;
        RECT 294.660 83.205 294.950 83.250 ;
        RECT 294.185 83.065 294.950 83.205 ;
        RECT 294.185 83.005 294.505 83.065 ;
        RECT 294.660 83.020 294.950 83.065 ;
        RECT 296.025 83.205 296.345 83.265 ;
        RECT 296.025 83.065 305.915 83.205 ;
        RECT 296.025 83.005 296.345 83.065 ;
        RECT 295.530 82.865 295.820 82.910 ;
        RECT 297.420 82.865 297.710 82.910 ;
        RECT 300.540 82.865 300.830 82.910 ;
        RECT 261.615 82.725 262.675 82.865 ;
        RECT 253.245 82.665 253.565 82.725 ;
        RECT 227.945 82.385 229.555 82.525 ;
        RECT 229.800 82.525 230.090 82.570 ;
        RECT 233.005 82.525 233.325 82.585 ;
        RECT 229.800 82.385 233.325 82.525 ;
        RECT 215.985 82.325 216.305 82.385 ;
        RECT 227.945 82.325 228.265 82.385 ;
        RECT 229.800 82.340 230.090 82.385 ;
        RECT 233.005 82.325 233.325 82.385 ;
        RECT 233.465 82.525 233.785 82.585 ;
        RECT 242.680 82.525 242.970 82.570 ;
        RECT 233.465 82.385 242.970 82.525 ;
        RECT 233.465 82.325 233.785 82.385 ;
        RECT 242.680 82.340 242.970 82.385 ;
        RECT 247.265 82.525 247.585 82.585 ;
        RECT 247.740 82.525 248.030 82.570 ;
        RECT 247.265 82.385 248.030 82.525 ;
        RECT 247.265 82.325 247.585 82.385 ;
        RECT 247.740 82.340 248.030 82.385 ;
        RECT 261.540 82.525 261.830 82.570 ;
        RECT 262.000 82.525 262.290 82.570 ;
        RECT 261.540 82.385 262.290 82.525 ;
        RECT 262.535 82.525 262.675 82.725 ;
        RECT 295.530 82.725 300.830 82.865 ;
        RECT 295.530 82.680 295.820 82.725 ;
        RECT 297.420 82.680 297.710 82.725 ;
        RECT 300.540 82.680 300.830 82.725 ;
        RECT 302.925 82.865 303.245 82.925 ;
        RECT 303.860 82.865 304.150 82.910 ;
        RECT 302.925 82.725 304.150 82.865 ;
        RECT 305.775 82.865 305.915 83.065 ;
        RECT 306.145 83.005 306.465 83.265 ;
        RECT 306.620 83.020 306.910 83.250 ;
        RECT 306.695 82.865 306.835 83.020 ;
        RECT 305.775 82.725 306.835 82.865 ;
        RECT 302.925 82.665 303.245 82.725 ;
        RECT 303.860 82.680 304.150 82.725 ;
        RECT 264.745 82.525 265.065 82.585 ;
        RECT 262.535 82.385 265.065 82.525 ;
        RECT 261.540 82.340 261.830 82.385 ;
        RECT 262.000 82.340 262.290 82.385 ;
        RECT 264.745 82.325 265.065 82.385 ;
        RECT 296.945 82.525 297.265 82.585 ;
        RECT 303.400 82.525 303.690 82.570 ;
        RECT 296.945 82.385 303.690 82.525 ;
        RECT 296.945 82.325 297.265 82.385 ;
        RECT 303.400 82.340 303.690 82.385 ;
        RECT 162.095 81.705 311.135 82.185 ;
        RECT 164.925 81.505 165.245 81.565 ;
        RECT 165.860 81.505 166.150 81.550 ;
        RECT 183.785 81.505 184.105 81.565 ;
        RECT 164.925 81.365 184.105 81.505 ;
        RECT 164.925 81.305 165.245 81.365 ;
        RECT 165.860 81.320 166.150 81.365 ;
        RECT 183.785 81.305 184.105 81.365 ;
        RECT 186.085 81.505 186.405 81.565 ;
        RECT 190.225 81.505 190.545 81.565 ;
        RECT 192.540 81.505 192.830 81.550 ;
        RECT 186.085 81.365 192.830 81.505 ;
        RECT 186.085 81.305 186.405 81.365 ;
        RECT 190.225 81.305 190.545 81.365 ;
        RECT 192.540 81.320 192.830 81.365 ;
        RECT 194.380 81.505 194.670 81.550 ;
        RECT 194.825 81.505 195.145 81.565 ;
        RECT 195.760 81.505 196.050 81.550 ;
        RECT 199.885 81.505 200.205 81.565 ;
        RECT 194.380 81.365 200.205 81.505 ;
        RECT 194.380 81.320 194.670 81.365 ;
        RECT 194.825 81.305 195.145 81.365 ;
        RECT 195.760 81.320 196.050 81.365 ;
        RECT 199.885 81.305 200.205 81.365 ;
        RECT 205.865 81.505 206.185 81.565 ;
        RECT 215.985 81.505 216.305 81.565 ;
        RECT 205.865 81.365 216.305 81.505 ;
        RECT 205.865 81.305 206.185 81.365 ;
        RECT 215.985 81.305 216.305 81.365 ;
        RECT 224.265 81.505 224.585 81.565 ;
        RECT 224.740 81.505 225.030 81.550 ;
        RECT 243.585 81.505 243.905 81.565 ;
        RECT 255.085 81.505 255.405 81.565 ;
        RECT 258.765 81.505 259.085 81.565 ;
        RECT 224.265 81.365 243.905 81.505 ;
        RECT 224.265 81.305 224.585 81.365 ;
        RECT 224.740 81.320 225.030 81.365 ;
        RECT 243.585 81.305 243.905 81.365 ;
        RECT 244.130 81.365 259.085 81.505 ;
        RECT 168.720 81.165 169.010 81.210 ;
        RECT 171.840 81.165 172.130 81.210 ;
        RECT 173.730 81.165 174.020 81.210 ;
        RECT 179.645 81.165 179.965 81.225 ;
        RECT 168.720 81.025 174.020 81.165 ;
        RECT 168.720 80.980 169.010 81.025 ;
        RECT 171.840 80.980 172.130 81.025 ;
        RECT 173.730 80.980 174.020 81.025 ;
        RECT 174.215 81.025 179.965 81.165 ;
        RECT 173.220 80.825 173.510 80.870 ;
        RECT 174.215 80.825 174.355 81.025 ;
        RECT 179.645 80.965 179.965 81.025 ;
        RECT 182.865 81.165 183.185 81.225 ;
        RECT 202.660 81.165 202.950 81.210 ;
        RECT 207.705 81.165 208.025 81.225 ;
        RECT 182.865 81.025 195.515 81.165 ;
        RECT 182.865 80.965 183.185 81.025 ;
        RECT 173.220 80.685 174.355 80.825 ;
        RECT 174.600 80.825 174.890 80.870 ;
        RECT 176.885 80.825 177.205 80.885 ;
        RECT 174.600 80.685 177.205 80.825 ;
        RECT 173.220 80.640 173.510 80.685 ;
        RECT 174.600 80.640 174.890 80.685 ;
        RECT 176.885 80.625 177.205 80.685 ;
        RECT 183.325 80.625 183.645 80.885 ;
        RECT 184.705 80.825 185.025 80.885 ;
        RECT 187.925 80.825 188.245 80.885 ;
        RECT 191.605 80.825 191.925 80.885 ;
        RECT 195.375 80.870 195.515 81.025 ;
        RECT 202.660 81.025 208.025 81.165 ;
        RECT 202.660 80.980 202.950 81.025 ;
        RECT 207.705 80.965 208.025 81.025 ;
        RECT 208.165 81.165 208.485 81.225 ;
        RECT 210.480 81.165 210.770 81.210 ;
        RECT 225.185 81.165 225.505 81.225 ;
        RECT 208.165 81.025 225.505 81.165 ;
        RECT 208.165 80.965 208.485 81.025 ;
        RECT 210.480 80.980 210.770 81.025 ;
        RECT 225.185 80.965 225.505 81.025 ;
        RECT 225.660 81.165 225.950 81.210 ;
        RECT 226.105 81.165 226.425 81.225 ;
        RECT 225.660 81.025 226.425 81.165 ;
        RECT 225.660 80.980 225.950 81.025 ;
        RECT 226.105 80.965 226.425 81.025 ;
        RECT 229.325 80.965 229.645 81.225 ;
        RECT 229.785 81.165 230.105 81.225 ;
        RECT 239.905 81.165 240.225 81.225 ;
        RECT 244.130 81.165 244.270 81.365 ;
        RECT 255.085 81.305 255.405 81.365 ;
        RECT 258.765 81.305 259.085 81.365 ;
        RECT 262.905 81.505 263.225 81.565 ;
        RECT 263.380 81.505 263.670 81.550 ;
        RECT 262.905 81.365 263.670 81.505 ;
        RECT 262.905 81.305 263.225 81.365 ;
        RECT 263.380 81.320 263.670 81.365 ;
        RECT 264.375 81.365 266.355 81.505 ;
        RECT 229.785 81.025 240.225 81.165 ;
        RECT 229.785 80.965 230.105 81.025 ;
        RECT 239.905 80.965 240.225 81.025 ;
        RECT 243.190 81.025 244.270 81.165 ;
        RECT 256.465 81.165 256.785 81.225 ;
        RECT 259.700 81.165 259.990 81.210 ;
        RECT 264.375 81.165 264.515 81.365 ;
        RECT 256.465 81.025 258.540 81.165 ;
        RECT 193.000 80.825 193.290 80.870 ;
        RECT 184.705 80.685 185.395 80.825 ;
        RECT 184.705 80.625 185.025 80.685 ;
        RECT 167.640 80.190 167.930 80.505 ;
        RECT 168.720 80.485 169.010 80.530 ;
        RECT 172.300 80.485 172.590 80.530 ;
        RECT 174.135 80.485 174.425 80.530 ;
        RECT 168.720 80.345 174.425 80.485 ;
        RECT 168.720 80.300 169.010 80.345 ;
        RECT 172.300 80.300 172.590 80.345 ;
        RECT 174.135 80.300 174.425 80.345 ;
        RECT 167.340 80.145 167.930 80.190 ;
        RECT 170.580 80.145 171.230 80.190 ;
        RECT 172.745 80.145 173.065 80.205 ;
        RECT 167.340 80.005 173.065 80.145 ;
        RECT 167.340 79.960 167.630 80.005 ;
        RECT 170.580 79.960 171.230 80.005 ;
        RECT 172.745 79.945 173.065 80.005 ;
        RECT 182.420 80.145 182.710 80.190 ;
        RECT 184.705 80.145 185.025 80.205 ;
        RECT 182.420 80.005 185.025 80.145 ;
        RECT 182.420 79.960 182.710 80.005 ;
        RECT 184.705 79.945 185.025 80.005 ;
        RECT 180.565 79.605 180.885 79.865 ;
        RECT 182.880 79.805 183.170 79.850 ;
        RECT 185.255 79.805 185.395 80.685 ;
        RECT 187.925 80.685 193.290 80.825 ;
        RECT 187.925 80.625 188.245 80.685 ;
        RECT 191.605 80.625 191.925 80.685 ;
        RECT 193.000 80.640 193.290 80.685 ;
        RECT 195.300 80.640 195.590 80.870 ;
        RECT 197.600 80.825 197.890 80.870 ;
        RECT 206.325 80.825 206.645 80.885 ;
        RECT 212.765 80.825 213.085 80.885 ;
        RECT 229.415 80.825 229.555 80.965 ;
        RECT 233.465 80.825 233.785 80.885 ;
        RECT 197.600 80.685 206.645 80.825 ;
        RECT 197.600 80.640 197.890 80.685 ;
        RECT 190.685 80.485 191.005 80.545 ;
        RECT 192.540 80.485 192.830 80.530 ;
        RECT 190.685 80.345 192.830 80.485 ;
        RECT 193.075 80.485 193.215 80.640 ;
        RECT 206.325 80.625 206.645 80.685 ;
        RECT 206.875 80.685 213.085 80.825 ;
        RECT 196.680 80.485 196.970 80.530 ;
        RECT 199.425 80.485 199.745 80.545 ;
        RECT 193.075 80.345 196.435 80.485 ;
        RECT 190.685 80.285 191.005 80.345 ;
        RECT 192.540 80.300 192.830 80.345 ;
        RECT 196.295 80.145 196.435 80.345 ;
        RECT 196.680 80.345 199.745 80.485 ;
        RECT 196.680 80.300 196.970 80.345 ;
        RECT 199.425 80.285 199.745 80.345 ;
        RECT 201.740 80.485 202.030 80.530 ;
        RECT 202.185 80.485 202.505 80.545 ;
        RECT 204.025 80.485 204.345 80.545 ;
        RECT 201.740 80.345 202.505 80.485 ;
        RECT 201.740 80.300 202.030 80.345 ;
        RECT 202.185 80.285 202.505 80.345 ;
        RECT 202.735 80.345 204.345 80.485 ;
        RECT 202.735 80.145 202.875 80.345 ;
        RECT 204.025 80.285 204.345 80.345 ;
        RECT 204.485 80.485 204.805 80.545 ;
        RECT 204.960 80.485 205.250 80.530 ;
        RECT 206.875 80.485 207.015 80.685 ;
        RECT 212.765 80.625 213.085 80.685 ;
        RECT 213.775 80.685 229.555 80.825 ;
        RECT 231.715 80.685 233.785 80.825 ;
        RECT 213.775 80.530 213.915 80.685 ;
        RECT 204.485 80.345 207.015 80.485 ;
        RECT 207.260 80.485 207.550 80.530 ;
        RECT 213.700 80.485 213.990 80.530 ;
        RECT 215.080 80.485 215.370 80.530 ;
        RECT 207.260 80.345 213.990 80.485 ;
        RECT 204.485 80.285 204.805 80.345 ;
        RECT 204.960 80.300 205.250 80.345 ;
        RECT 207.260 80.300 207.550 80.345 ;
        RECT 213.700 80.300 213.990 80.345 ;
        RECT 214.235 80.345 217.135 80.485 ;
        RECT 196.295 80.005 202.875 80.145 ;
        RECT 203.105 80.145 203.425 80.205 ;
        RECT 207.335 80.145 207.475 80.300 ;
        RECT 203.105 80.005 207.475 80.145 ;
        RECT 208.625 80.145 208.945 80.205 ;
        RECT 210.940 80.145 211.230 80.190 ;
        RECT 214.235 80.145 214.375 80.345 ;
        RECT 215.080 80.300 215.370 80.345 ;
        RECT 208.625 80.005 211.230 80.145 ;
        RECT 203.105 79.945 203.425 80.005 ;
        RECT 208.625 79.945 208.945 80.005 ;
        RECT 210.940 79.960 211.230 80.005 ;
        RECT 213.775 80.005 214.375 80.145 ;
        RECT 216.995 80.145 217.135 80.345 ;
        RECT 217.365 80.285 217.685 80.545 ;
        RECT 225.185 80.485 225.505 80.545 ;
        RECT 227.025 80.485 227.345 80.545 ;
        RECT 231.715 80.530 231.855 80.685 ;
        RECT 233.465 80.625 233.785 80.685 ;
        RECT 239.445 80.825 239.765 80.885 ;
        RECT 243.190 80.825 243.330 81.025 ;
        RECT 256.465 80.965 256.785 81.025 ;
        RECT 254.165 80.825 254.485 80.885 ;
        RECT 258.400 80.825 258.540 81.025 ;
        RECT 259.700 81.025 264.515 81.165 ;
        RECT 259.700 80.980 259.990 81.025 ;
        RECT 264.745 80.965 265.065 81.225 ;
        RECT 239.445 80.685 243.330 80.825 ;
        RECT 239.445 80.625 239.765 80.685 ;
        RECT 229.110 80.485 229.400 80.530 ;
        RECT 217.915 80.345 220.815 80.485 ;
        RECT 217.915 80.145 218.055 80.345 ;
        RECT 216.995 80.005 218.055 80.145 ;
        RECT 220.675 80.145 220.815 80.345 ;
        RECT 225.185 80.345 229.400 80.485 ;
        RECT 225.185 80.285 225.505 80.345 ;
        RECT 227.025 80.285 227.345 80.345 ;
        RECT 229.110 80.300 229.400 80.345 ;
        RECT 231.175 80.300 231.465 80.530 ;
        RECT 231.640 80.300 231.930 80.530 ;
        RECT 223.820 80.145 224.110 80.190 ;
        RECT 227.485 80.145 227.805 80.205 ;
        RECT 220.675 80.005 227.805 80.145 ;
        RECT 185.625 79.805 185.945 79.865 ;
        RECT 182.880 79.665 185.945 79.805 ;
        RECT 182.880 79.620 183.170 79.665 ;
        RECT 185.625 79.605 185.945 79.665 ;
        RECT 204.025 79.805 204.345 79.865 ;
        RECT 213.775 79.805 213.915 80.005 ;
        RECT 223.820 79.960 224.110 80.005 ;
        RECT 227.485 79.945 227.805 80.005 ;
        RECT 229.785 79.945 230.105 80.205 ;
        RECT 230.260 80.145 230.550 80.190 ;
        RECT 230.705 80.145 231.025 80.205 ;
        RECT 230.260 80.005 231.025 80.145 ;
        RECT 231.255 80.145 231.395 80.300 ;
        RECT 233.005 80.285 233.325 80.545 ;
        RECT 233.925 80.285 234.245 80.545 ;
        RECT 234.385 80.475 234.705 80.545 ;
        RECT 238.525 80.485 238.845 80.545 ;
        RECT 239.000 80.485 239.290 80.530 ;
        RECT 234.385 80.335 235.075 80.475 ;
        RECT 234.385 80.285 234.705 80.335 ;
        RECT 233.465 80.145 233.785 80.205 ;
        RECT 231.255 80.005 233.785 80.145 ;
        RECT 234.935 80.145 235.075 80.335 ;
        RECT 238.525 80.345 239.290 80.485 ;
        RECT 238.525 80.285 238.845 80.345 ;
        RECT 239.000 80.300 239.290 80.345 ;
        RECT 239.905 80.285 240.225 80.545 ;
        RECT 240.365 80.285 240.685 80.545 ;
        RECT 240.840 80.485 241.130 80.530 ;
        RECT 241.745 80.485 242.065 80.545 ;
        RECT 243.190 80.530 243.330 80.685 ;
        RECT 244.130 80.685 256.005 80.825 ;
        RECT 258.400 80.685 260.375 80.825 ;
        RECT 244.130 80.545 244.270 80.685 ;
        RECT 254.165 80.625 254.485 80.685 ;
        RECT 240.840 80.345 242.065 80.485 ;
        RECT 240.840 80.300 241.130 80.345 ;
        RECT 240.915 80.145 241.055 80.300 ;
        RECT 241.745 80.285 242.065 80.345 ;
        RECT 243.115 80.300 243.405 80.530 ;
        RECT 244.045 80.285 244.365 80.545 ;
        RECT 244.505 80.530 244.825 80.545 ;
        RECT 244.505 80.300 244.990 80.530 ;
        RECT 245.440 80.485 245.730 80.530 ;
        RECT 245.885 80.485 246.205 80.545 ;
        RECT 245.440 80.345 246.205 80.485 ;
        RECT 245.440 80.300 245.730 80.345 ;
        RECT 244.505 80.285 244.825 80.300 ;
        RECT 245.885 80.285 246.205 80.345 ;
        RECT 246.805 80.285 247.125 80.545 ;
        RECT 248.645 80.285 248.965 80.545 ;
        RECT 249.105 80.485 249.425 80.545 ;
        RECT 250.040 80.485 250.330 80.530 ;
        RECT 249.105 80.345 250.330 80.485 ;
        RECT 249.105 80.285 249.425 80.345 ;
        RECT 250.040 80.300 250.330 80.345 ;
        RECT 250.945 80.285 251.265 80.545 ;
        RECT 255.865 80.485 256.005 80.685 ;
        RECT 255.865 80.345 256.235 80.485 ;
        RECT 243.600 80.145 243.890 80.190 ;
        RECT 234.935 80.005 241.055 80.145 ;
        RECT 241.375 80.005 243.890 80.145 ;
        RECT 230.260 79.960 230.550 80.005 ;
        RECT 230.705 79.945 231.025 80.005 ;
        RECT 233.465 79.945 233.785 80.005 ;
        RECT 241.375 79.865 241.515 80.005 ;
        RECT 243.600 79.960 243.890 80.005 ;
        RECT 247.265 79.945 247.585 80.205 ;
        RECT 247.740 80.145 248.030 80.190 ;
        RECT 253.245 80.145 253.565 80.205 ;
        RECT 247.740 80.005 253.565 80.145 ;
        RECT 256.095 80.145 256.235 80.345 ;
        RECT 256.465 80.285 256.785 80.545 ;
        RECT 256.925 80.485 257.245 80.545 ;
        RECT 256.925 80.345 257.440 80.485 ;
        RECT 256.925 80.285 257.245 80.345 ;
        RECT 257.860 80.300 258.150 80.530 ;
        RECT 257.935 80.145 258.075 80.300 ;
        RECT 258.305 80.285 258.625 80.545 ;
        RECT 258.765 80.530 259.085 80.545 ;
        RECT 260.235 80.530 260.375 80.685 ;
        RECT 258.765 80.485 259.095 80.530 ;
        RECT 258.765 80.345 259.280 80.485 ;
        RECT 258.765 80.300 259.095 80.345 ;
        RECT 260.160 80.300 260.450 80.530 ;
        RECT 258.765 80.285 259.085 80.300 ;
        RECT 260.605 80.285 260.925 80.545 ;
        RECT 262.485 80.485 262.775 80.530 ;
        RECT 261.155 80.345 262.775 80.485 ;
        RECT 261.155 80.145 261.295 80.345 ;
        RECT 262.485 80.300 262.775 80.345 ;
        RECT 263.840 80.485 264.130 80.530 ;
        RECT 264.285 80.485 264.605 80.545 ;
        RECT 264.835 80.530 264.975 80.965 ;
        RECT 263.840 80.345 264.605 80.485 ;
        RECT 263.840 80.300 264.130 80.345 ;
        RECT 264.285 80.285 264.605 80.345 ;
        RECT 264.760 80.300 265.050 80.530 ;
        RECT 265.220 80.300 265.510 80.530 ;
        RECT 256.095 80.005 261.295 80.145 ;
        RECT 247.740 79.960 248.030 80.005 ;
        RECT 248.275 79.865 248.415 80.005 ;
        RECT 253.245 79.945 253.565 80.005 ;
        RECT 261.525 79.945 261.845 80.205 ;
        RECT 261.985 79.945 262.305 80.205 ;
        RECT 265.295 80.145 265.435 80.300 ;
        RECT 265.665 80.285 265.985 80.545 ;
        RECT 266.215 80.485 266.355 81.365 ;
        RECT 267.045 81.305 267.365 81.565 ;
        RECT 269.345 81.305 269.665 81.565 ;
        RECT 276.245 81.505 276.565 81.565 ;
        RECT 277.180 81.505 277.470 81.550 ;
        RECT 276.245 81.365 277.470 81.505 ;
        RECT 276.245 81.305 276.565 81.365 ;
        RECT 277.180 81.320 277.470 81.365 ;
        RECT 280.385 81.505 280.705 81.565 ;
        RECT 302.940 81.505 303.230 81.550 ;
        RECT 280.385 81.365 303.230 81.505 ;
        RECT 280.385 81.305 280.705 81.365 ;
        RECT 302.940 81.320 303.230 81.365 ;
        RECT 266.600 81.165 266.890 81.210 ;
        RECT 278.545 81.165 278.865 81.225 ;
        RECT 284.065 81.165 284.385 81.225 ;
        RECT 266.600 81.025 267.735 81.165 ;
        RECT 266.600 80.980 266.890 81.025 ;
        RECT 267.595 80.870 267.735 81.025 ;
        RECT 278.545 81.025 284.385 81.165 ;
        RECT 278.545 80.965 278.865 81.025 ;
        RECT 284.065 80.965 284.385 81.025 ;
        RECT 295.070 81.165 295.360 81.210 ;
        RECT 296.960 81.165 297.250 81.210 ;
        RECT 300.080 81.165 300.370 81.210 ;
        RECT 295.070 81.025 300.370 81.165 ;
        RECT 295.070 80.980 295.360 81.025 ;
        RECT 296.960 80.980 297.250 81.025 ;
        RECT 300.080 80.980 300.370 81.025 ;
        RECT 267.520 80.640 267.810 80.870 ;
        RECT 276.705 80.825 277.025 80.885 ;
        RECT 280.385 80.825 280.705 80.885 ;
        RECT 276.705 80.685 280.705 80.825 ;
        RECT 276.705 80.625 277.025 80.685 ;
        RECT 280.385 80.625 280.705 80.685 ;
        RECT 281.765 80.825 282.085 80.885 ;
        RECT 282.685 80.825 283.005 80.885 ;
        RECT 281.765 80.685 283.005 80.825 ;
        RECT 281.765 80.625 282.085 80.685 ;
        RECT 282.685 80.625 283.005 80.685 ;
        RECT 283.145 80.625 283.465 80.885 ;
        RECT 286.365 80.825 286.685 80.885 ;
        RECT 291.440 80.825 291.730 80.870 ;
        RECT 286.365 80.685 291.730 80.825 ;
        RECT 286.365 80.625 286.685 80.685 ;
        RECT 291.440 80.640 291.730 80.685 ;
        RECT 267.060 80.485 267.350 80.530 ;
        RECT 266.215 80.345 267.350 80.485 ;
        RECT 267.060 80.300 267.350 80.345 ;
        RECT 268.425 80.285 268.745 80.545 ;
        RECT 269.805 80.485 270.125 80.545 ;
        RECT 275.340 80.485 275.630 80.530 ;
        RECT 269.805 80.345 275.630 80.485 ;
        RECT 269.805 80.285 270.125 80.345 ;
        RECT 275.340 80.300 275.630 80.345 ;
        RECT 275.785 80.485 276.105 80.545 ;
        RECT 276.260 80.485 276.550 80.530 ;
        RECT 278.085 80.485 278.405 80.545 ;
        RECT 275.785 80.345 278.405 80.485 ;
        RECT 275.785 80.285 276.105 80.345 ;
        RECT 276.260 80.300 276.550 80.345 ;
        RECT 278.085 80.285 278.405 80.345 ;
        RECT 290.505 80.485 290.825 80.545 ;
        RECT 294.185 80.485 294.505 80.545 ;
        RECT 290.505 80.345 294.505 80.485 ;
        RECT 290.505 80.285 290.825 80.345 ;
        RECT 294.185 80.285 294.505 80.345 ;
        RECT 294.665 80.485 294.955 80.530 ;
        RECT 296.500 80.485 296.790 80.530 ;
        RECT 300.080 80.485 300.370 80.530 ;
        RECT 294.665 80.345 300.370 80.485 ;
        RECT 294.665 80.300 294.955 80.345 ;
        RECT 296.500 80.300 296.790 80.345 ;
        RECT 300.080 80.300 300.370 80.345 ;
        RECT 281.305 80.145 281.625 80.205 ;
        RECT 282.240 80.145 282.530 80.190 ;
        RECT 284.065 80.145 284.385 80.205 ;
        RECT 264.835 80.005 281.995 80.145 ;
        RECT 264.835 79.865 264.975 80.005 ;
        RECT 281.305 79.945 281.625 80.005 ;
        RECT 204.025 79.665 213.915 79.805 ;
        RECT 223.345 79.805 223.665 79.865 ;
        RECT 224.740 79.805 225.030 79.850 ;
        RECT 223.345 79.665 225.030 79.805 ;
        RECT 204.025 79.605 204.345 79.665 ;
        RECT 223.345 79.605 223.665 79.665 ;
        RECT 224.740 79.620 225.030 79.665 ;
        RECT 228.420 79.805 228.710 79.850 ;
        RECT 228.865 79.805 229.185 79.865 ;
        RECT 228.420 79.665 229.185 79.805 ;
        RECT 228.420 79.620 228.710 79.665 ;
        RECT 228.865 79.605 229.185 79.665 ;
        RECT 232.085 79.605 232.405 79.865 ;
        RECT 241.285 79.605 241.605 79.865 ;
        RECT 241.745 79.605 242.065 79.865 ;
        RECT 242.205 79.605 242.525 79.865 ;
        RECT 244.505 79.805 244.825 79.865 ;
        RECT 245.900 79.805 246.190 79.850 ;
        RECT 244.505 79.665 246.190 79.805 ;
        RECT 244.505 79.605 244.825 79.665 ;
        RECT 245.900 79.620 246.190 79.665 ;
        RECT 248.185 79.605 248.505 79.865 ;
        RECT 249.105 79.605 249.425 79.865 ;
        RECT 249.565 79.805 249.885 79.865 ;
        RECT 255.545 79.805 255.865 79.865 ;
        RECT 258.765 79.805 259.085 79.865 ;
        RECT 249.565 79.665 259.085 79.805 ;
        RECT 249.565 79.605 249.885 79.665 ;
        RECT 255.545 79.605 255.865 79.665 ;
        RECT 258.765 79.605 259.085 79.665 ;
        RECT 264.745 79.605 265.065 79.865 ;
        RECT 280.385 79.605 280.705 79.865 ;
        RECT 281.855 79.805 281.995 80.005 ;
        RECT 282.240 80.005 284.385 80.145 ;
        RECT 282.240 79.960 282.530 80.005 ;
        RECT 284.065 79.945 284.385 80.005 ;
        RECT 285.905 80.145 286.225 80.205 ;
        RECT 287.760 80.145 288.050 80.190 ;
        RECT 285.905 80.005 288.050 80.145 ;
        RECT 285.905 79.945 286.225 80.005 ;
        RECT 287.760 79.960 288.050 80.005 ;
        RECT 295.565 79.945 295.885 80.205 ;
        RECT 301.160 80.190 301.450 80.505 ;
        RECT 297.860 80.145 298.510 80.190 ;
        RECT 301.160 80.145 301.750 80.190 ;
        RECT 302.465 80.145 302.785 80.205 ;
        RECT 303.845 80.145 304.165 80.205 ;
        RECT 297.860 80.005 304.165 80.145 ;
        RECT 297.860 79.960 298.510 80.005 ;
        RECT 301.460 79.960 301.750 80.005 ;
        RECT 302.465 79.945 302.785 80.005 ;
        RECT 303.845 79.945 304.165 80.005 ;
        RECT 304.765 80.145 305.085 80.205 ;
        RECT 305.685 80.145 306.005 80.205 ;
        RECT 304.765 80.005 306.005 80.145 ;
        RECT 304.765 79.945 305.085 80.005 ;
        RECT 305.685 79.945 306.005 80.005 ;
        RECT 296.945 79.805 297.265 79.865 ;
        RECT 281.855 79.665 297.265 79.805 ;
        RECT 296.945 79.605 297.265 79.665 ;
        RECT 162.095 78.985 311.135 79.465 ;
        RECT 176.885 78.785 177.205 78.845 ;
        RECT 204.025 78.785 204.345 78.845 ;
        RECT 205.005 78.785 205.295 78.830 ;
        RECT 176.885 78.645 189.075 78.785 ;
        RECT 176.885 78.585 177.205 78.645 ;
        RECT 173.665 78.445 173.985 78.505 ;
        RECT 175.060 78.445 175.350 78.490 ;
        RECT 179.645 78.445 179.965 78.505 ;
        RECT 173.665 78.305 179.965 78.445 ;
        RECT 173.665 78.245 173.985 78.305 ;
        RECT 175.060 78.260 175.350 78.305 ;
        RECT 179.645 78.245 179.965 78.305 ;
        RECT 180.560 78.445 181.210 78.490 ;
        RECT 184.160 78.445 184.450 78.490 ;
        RECT 180.560 78.305 184.450 78.445 ;
        RECT 180.560 78.260 181.210 78.305 ;
        RECT 183.860 78.260 184.450 78.305 ;
        RECT 174.125 78.105 174.445 78.165 ;
        RECT 174.600 78.105 174.890 78.150 ;
        RECT 174.125 77.965 174.890 78.105 ;
        RECT 174.125 77.905 174.445 77.965 ;
        RECT 174.600 77.920 174.890 77.965 ;
        RECT 176.885 77.905 177.205 78.165 ;
        RECT 177.365 78.105 177.655 78.150 ;
        RECT 179.200 78.105 179.490 78.150 ;
        RECT 182.780 78.105 183.070 78.150 ;
        RECT 177.365 77.965 183.070 78.105 ;
        RECT 177.365 77.920 177.655 77.965 ;
        RECT 179.200 77.920 179.490 77.965 ;
        RECT 182.780 77.920 183.070 77.965 ;
        RECT 183.860 77.945 184.150 78.260 ;
        RECT 175.980 77.765 176.270 77.810 ;
        RECT 178.280 77.765 178.570 77.810 ;
        RECT 180.565 77.765 180.885 77.825 ;
        RECT 175.980 77.625 177.575 77.765 ;
        RECT 175.980 77.580 176.270 77.625 ;
        RECT 172.760 77.085 173.050 77.130 ;
        RECT 175.965 77.085 176.285 77.145 ;
        RECT 172.760 76.945 176.285 77.085 ;
        RECT 177.435 77.085 177.575 77.625 ;
        RECT 178.280 77.625 180.885 77.765 ;
        RECT 178.280 77.580 178.570 77.625 ;
        RECT 180.565 77.565 180.885 77.625 ;
        RECT 181.945 77.765 182.265 77.825 ;
        RECT 183.875 77.765 184.015 77.945 ;
        RECT 188.385 77.905 188.705 78.165 ;
        RECT 188.935 78.105 189.075 78.645 ;
        RECT 204.025 78.645 205.295 78.785 ;
        RECT 204.025 78.585 204.345 78.645 ;
        RECT 205.005 78.600 205.295 78.645 ;
        RECT 206.325 78.785 206.645 78.845 ;
        RECT 213.685 78.785 214.005 78.845 ;
        RECT 206.325 78.645 214.005 78.785 ;
        RECT 206.325 78.585 206.645 78.645 ;
        RECT 213.685 78.585 214.005 78.645 ;
        RECT 215.985 78.585 216.305 78.845 ;
        RECT 216.445 78.785 216.765 78.845 ;
        RECT 217.380 78.785 217.670 78.830 ;
        RECT 219.205 78.785 219.525 78.845 ;
        RECT 216.445 78.645 219.525 78.785 ;
        RECT 216.445 78.585 216.765 78.645 ;
        RECT 217.380 78.600 217.670 78.645 ;
        RECT 219.205 78.585 219.525 78.645 ;
        RECT 228.465 78.785 228.755 78.830 ;
        RECT 229.325 78.785 229.645 78.845 ;
        RECT 228.465 78.645 229.645 78.785 ;
        RECT 228.465 78.600 228.755 78.645 ;
        RECT 229.325 78.585 229.645 78.645 ;
        RECT 239.905 78.785 240.225 78.845 ;
        RECT 258.305 78.785 258.625 78.845 ;
        RECT 239.905 78.645 258.625 78.785 ;
        RECT 239.905 78.585 240.225 78.645 ;
        RECT 258.305 78.585 258.625 78.645 ;
        RECT 258.765 78.585 259.085 78.845 ;
        RECT 259.685 78.785 260.005 78.845 ;
        RECT 260.160 78.785 260.450 78.830 ;
        RECT 261.065 78.785 261.385 78.845 ;
        RECT 259.685 78.645 260.450 78.785 ;
        RECT 259.685 78.585 260.005 78.645 ;
        RECT 260.160 78.600 260.450 78.645 ;
        RECT 260.720 78.645 261.385 78.785 ;
        RECT 190.225 78.445 190.545 78.505 ;
        RECT 198.060 78.445 198.350 78.490 ;
        RECT 216.075 78.445 216.215 78.585 ;
        RECT 216.920 78.445 217.210 78.490 ;
        RECT 190.225 78.305 203.795 78.445 ;
        RECT 216.075 78.305 217.210 78.445 ;
        RECT 190.225 78.245 190.545 78.305 ;
        RECT 198.060 78.260 198.350 78.305 ;
        RECT 191.620 78.105 191.910 78.150 ;
        RECT 193.920 78.105 194.210 78.150 ;
        RECT 188.935 77.965 194.210 78.105 ;
        RECT 191.620 77.920 191.910 77.965 ;
        RECT 193.920 77.920 194.210 77.965 ;
        RECT 197.585 78.105 197.905 78.165 ;
        RECT 198.520 78.105 198.810 78.150 ;
        RECT 197.585 77.965 198.810 78.105 ;
        RECT 197.585 77.905 197.905 77.965 ;
        RECT 198.520 77.920 198.810 77.965 ;
        RECT 199.425 77.905 199.745 78.165 ;
        RECT 199.885 77.905 200.205 78.165 ;
        RECT 200.360 77.920 200.650 78.150 ;
        RECT 186.545 77.765 186.865 77.825 ;
        RECT 188.845 77.765 189.165 77.825 ;
        RECT 192.525 77.765 192.845 77.825 ;
        RECT 181.945 77.625 192.845 77.765 ;
        RECT 181.945 77.565 182.265 77.625 ;
        RECT 186.545 77.565 186.865 77.625 ;
        RECT 188.845 77.565 189.165 77.625 ;
        RECT 192.525 77.565 192.845 77.625 ;
        RECT 198.045 77.765 198.365 77.825 ;
        RECT 200.435 77.765 200.575 77.920 ;
        RECT 203.105 77.905 203.425 78.165 ;
        RECT 203.655 78.105 203.795 78.305 ;
        RECT 216.920 78.260 217.210 78.305 ;
        RECT 217.825 78.445 218.145 78.505 ;
        RECT 226.580 78.445 226.870 78.490 ;
        RECT 227.485 78.445 227.805 78.505 ;
        RECT 217.825 78.305 221.505 78.445 ;
        RECT 217.825 78.245 218.145 78.305 ;
        RECT 206.800 78.105 207.090 78.150 ;
        RECT 212.305 78.105 212.625 78.165 ;
        RECT 203.655 77.965 207.090 78.105 ;
        RECT 206.800 77.920 207.090 77.965 ;
        RECT 207.335 77.965 212.625 78.105 ;
        RECT 207.335 77.765 207.475 77.965 ;
        RECT 212.305 77.905 212.625 77.965 ;
        RECT 213.685 78.105 214.005 78.165 ;
        RECT 219.220 78.105 219.510 78.150 ;
        RECT 213.685 77.965 219.510 78.105 ;
        RECT 213.685 77.905 214.005 77.965 ;
        RECT 219.220 77.920 219.510 77.965 ;
        RECT 220.125 77.905 220.445 78.165 ;
        RECT 221.365 78.105 221.505 78.305 ;
        RECT 226.580 78.305 227.805 78.445 ;
        RECT 226.580 78.260 226.870 78.305 ;
        RECT 227.485 78.245 227.805 78.305 ;
        RECT 231.165 78.445 231.485 78.505 ;
        RECT 241.745 78.445 242.065 78.505 ;
        RECT 243.140 78.445 243.430 78.490 ;
        RECT 231.165 78.305 237.375 78.445 ;
        RECT 231.165 78.245 231.485 78.305 ;
        RECT 224.740 78.105 225.030 78.150 ;
        RECT 221.365 77.965 225.030 78.105 ;
        RECT 237.235 78.105 237.375 78.305 ;
        RECT 241.745 78.305 243.430 78.445 ;
        RECT 241.745 78.245 242.065 78.305 ;
        RECT 243.140 78.260 243.430 78.305 ;
        RECT 256.005 78.445 256.325 78.505 ;
        RECT 257.845 78.445 258.165 78.505 ;
        RECT 256.005 78.305 258.165 78.445 ;
        RECT 258.855 78.445 258.995 78.585 ;
        RECT 260.720 78.445 260.860 78.645 ;
        RECT 261.065 78.585 261.385 78.645 ;
        RECT 263.380 78.785 263.670 78.830 ;
        RECT 267.045 78.785 267.365 78.845 ;
        RECT 263.380 78.645 267.365 78.785 ;
        RECT 263.380 78.600 263.670 78.645 ;
        RECT 267.045 78.585 267.365 78.645 ;
        RECT 267.520 78.785 267.810 78.830 ;
        RECT 268.425 78.785 268.745 78.845 ;
        RECT 267.520 78.645 268.745 78.785 ;
        RECT 267.520 78.600 267.810 78.645 ;
        RECT 268.425 78.585 268.745 78.645 ;
        RECT 279.005 78.585 279.325 78.845 ;
        RECT 279.095 78.445 279.235 78.585 ;
        RECT 258.855 78.305 260.860 78.445 ;
        RECT 276.795 78.305 279.235 78.445 ;
        RECT 280.380 78.445 281.030 78.490 ;
        RECT 283.980 78.445 284.270 78.490 ;
        RECT 280.380 78.305 284.270 78.445 ;
        RECT 256.005 78.245 256.325 78.305 ;
        RECT 257.845 78.245 258.165 78.305 ;
        RECT 244.520 78.105 244.810 78.150 ;
        RECT 249.105 78.105 249.425 78.165 ;
        RECT 237.235 77.965 244.270 78.105 ;
        RECT 224.740 77.920 225.030 77.965 ;
        RECT 198.045 77.625 200.575 77.765 ;
        RECT 201.355 77.625 207.475 77.765 ;
        RECT 198.045 77.565 198.365 77.625 ;
        RECT 177.770 77.425 178.060 77.470 ;
        RECT 179.660 77.425 179.950 77.470 ;
        RECT 182.780 77.425 183.070 77.470 ;
        RECT 177.770 77.285 183.070 77.425 ;
        RECT 177.770 77.240 178.060 77.285 ;
        RECT 179.660 77.240 179.950 77.285 ;
        RECT 182.780 77.240 183.070 77.285 ;
        RECT 185.625 77.225 185.945 77.485 ;
        RECT 180.105 77.085 180.425 77.145 ;
        RECT 183.325 77.085 183.645 77.145 ;
        RECT 177.435 76.945 183.645 77.085 ;
        RECT 172.760 76.900 173.050 76.945 ;
        RECT 175.965 76.885 176.285 76.945 ;
        RECT 180.105 76.885 180.425 76.945 ;
        RECT 183.325 76.885 183.645 76.945 ;
        RECT 187.005 77.085 187.325 77.145 ;
        RECT 192.065 77.085 192.385 77.145 ;
        RECT 201.355 77.085 201.495 77.625 ;
        RECT 210.465 77.565 210.785 77.825 ;
        RECT 211.845 77.765 212.165 77.825 ;
        RECT 211.845 77.625 217.135 77.765 ;
        RECT 211.845 77.565 212.165 77.625 ;
        RECT 204.025 77.425 204.345 77.485 ;
        RECT 204.025 77.285 205.635 77.425 ;
        RECT 204.025 77.225 204.345 77.285 ;
        RECT 187.005 76.945 201.495 77.085 ;
        RECT 187.005 76.885 187.325 76.945 ;
        RECT 192.065 76.885 192.385 76.945 ;
        RECT 201.725 76.885 202.045 77.145 ;
        RECT 204.485 77.085 204.805 77.145 ;
        RECT 204.960 77.085 205.250 77.130 ;
        RECT 204.485 76.945 205.250 77.085 ;
        RECT 205.495 77.085 205.635 77.285 ;
        RECT 205.865 77.225 206.185 77.485 ;
        RECT 211.385 77.425 211.705 77.485 ;
        RECT 216.995 77.425 217.135 77.625 ;
        RECT 217.840 77.580 218.130 77.810 ;
        RECT 226.120 77.765 226.410 77.810 ;
        RECT 232.085 77.765 232.405 77.825 ;
        RECT 226.120 77.625 232.405 77.765 ;
        RECT 226.120 77.580 226.410 77.625 ;
        RECT 217.915 77.425 218.055 77.580 ;
        RECT 232.085 77.565 232.405 77.625 ;
        RECT 242.205 77.765 242.525 77.825 ;
        RECT 243.600 77.765 243.890 77.810 ;
        RECT 242.205 77.625 243.890 77.765 ;
        RECT 244.130 77.765 244.270 77.965 ;
        RECT 244.520 77.965 249.425 78.105 ;
        RECT 244.520 77.920 244.810 77.965 ;
        RECT 249.105 77.905 249.425 77.965 ;
        RECT 252.325 78.105 252.645 78.165 ;
        RECT 255.085 78.105 255.405 78.165 ;
        RECT 257.400 78.105 257.690 78.150 ;
        RECT 252.325 77.965 257.690 78.105 ;
        RECT 252.325 77.905 252.645 77.965 ;
        RECT 255.085 77.905 255.405 77.965 ;
        RECT 257.400 77.920 257.690 77.965 ;
        RECT 258.305 77.905 258.625 78.165 ;
        RECT 258.765 77.905 259.085 78.165 ;
        RECT 259.315 78.150 259.455 78.305 ;
        RECT 259.240 77.920 259.530 78.150 ;
        RECT 260.605 77.905 260.925 78.165 ;
        RECT 261.525 77.905 261.845 78.165 ;
        RECT 261.985 77.905 262.305 78.165 ;
        RECT 262.460 77.920 262.750 78.150 ;
        RECT 256.465 77.765 256.785 77.825 ;
        RECT 257.845 77.765 258.165 77.825 ;
        RECT 261.065 77.765 261.385 77.825 ;
        RECT 262.535 77.765 262.675 77.920 ;
        RECT 266.585 77.905 266.905 78.165 ;
        RECT 276.795 78.150 276.935 78.305 ;
        RECT 280.380 78.260 281.030 78.305 ;
        RECT 283.680 78.260 284.270 78.305 ;
        RECT 283.680 78.165 283.970 78.260 ;
        RECT 285.905 78.245 286.225 78.505 ;
        RECT 276.720 77.920 277.010 78.150 ;
        RECT 277.185 78.105 277.475 78.150 ;
        RECT 279.020 78.105 279.310 78.150 ;
        RECT 282.600 78.105 282.890 78.150 ;
        RECT 277.185 77.965 282.890 78.105 ;
        RECT 277.185 77.920 277.475 77.965 ;
        RECT 279.020 77.920 279.310 77.965 ;
        RECT 282.600 77.920 282.890 77.965 ;
        RECT 283.605 78.105 283.970 78.165 ;
        RECT 286.825 78.105 287.145 78.165 ;
        RECT 283.605 77.965 287.145 78.105 ;
        RECT 283.605 77.945 283.970 77.965 ;
        RECT 283.605 77.905 283.925 77.945 ;
        RECT 286.825 77.905 287.145 77.965 ;
        RECT 291.440 77.920 291.730 78.150 ;
        RECT 244.130 77.625 246.115 77.765 ;
        RECT 242.205 77.565 242.525 77.625 ;
        RECT 243.600 77.580 243.890 77.625 ;
        RECT 211.385 77.285 216.675 77.425 ;
        RECT 216.995 77.285 218.055 77.425 ;
        RECT 218.285 77.425 218.605 77.485 ;
        RECT 225.660 77.425 225.950 77.470 ;
        RECT 228.865 77.425 229.185 77.485 ;
        RECT 218.285 77.285 225.415 77.425 ;
        RECT 211.385 77.225 211.705 77.285 ;
        RECT 214.145 77.085 214.465 77.145 ;
        RECT 205.495 76.945 214.465 77.085 ;
        RECT 204.485 76.885 204.805 76.945 ;
        RECT 204.960 76.900 205.250 76.945 ;
        RECT 214.145 76.885 214.465 76.945 ;
        RECT 215.080 77.085 215.370 77.130 ;
        RECT 215.985 77.085 216.305 77.145 ;
        RECT 215.080 76.945 216.305 77.085 ;
        RECT 216.535 77.085 216.675 77.285 ;
        RECT 218.285 77.225 218.605 77.285 ;
        RECT 221.060 77.085 221.350 77.130 ;
        RECT 216.535 76.945 221.350 77.085 ;
        RECT 215.080 76.900 215.370 76.945 ;
        RECT 215.985 76.885 216.305 76.945 ;
        RECT 221.060 76.900 221.350 76.945 ;
        RECT 223.805 76.885 224.125 77.145 ;
        RECT 225.275 77.085 225.415 77.285 ;
        RECT 225.660 77.285 229.185 77.425 ;
        RECT 225.660 77.240 225.950 77.285 ;
        RECT 228.865 77.225 229.185 77.285 ;
        RECT 233.005 77.425 233.325 77.485 ;
        RECT 245.440 77.425 245.730 77.470 ;
        RECT 233.005 77.285 245.730 77.425 ;
        RECT 233.005 77.225 233.325 77.285 ;
        RECT 245.440 77.240 245.730 77.285 ;
        RECT 228.405 77.085 228.725 77.145 ;
        RECT 225.275 76.945 228.725 77.085 ;
        RECT 228.405 76.885 228.725 76.945 ;
        RECT 229.340 77.085 229.630 77.130 ;
        RECT 230.705 77.085 231.025 77.145 ;
        RECT 229.340 76.945 231.025 77.085 ;
        RECT 229.340 76.900 229.630 76.945 ;
        RECT 230.705 76.885 231.025 76.945 ;
        RECT 233.465 77.085 233.785 77.145 ;
        RECT 243.585 77.085 243.905 77.145 ;
        RECT 233.465 76.945 243.905 77.085 ;
        RECT 233.465 76.885 233.785 76.945 ;
        RECT 243.585 76.885 243.905 76.945 ;
        RECT 244.505 76.885 244.825 77.145 ;
        RECT 245.975 77.085 246.115 77.625 ;
        RECT 256.465 77.625 258.165 77.765 ;
        RECT 256.465 77.565 256.785 77.625 ;
        RECT 257.845 77.565 258.165 77.625 ;
        RECT 258.400 77.625 260.860 77.765 ;
        RECT 258.400 77.085 258.540 77.625 ;
        RECT 260.720 77.425 260.860 77.625 ;
        RECT 261.065 77.625 262.675 77.765 ;
        RECT 265.205 77.765 265.525 77.825 ;
        RECT 265.680 77.765 265.970 77.810 ;
        RECT 265.205 77.625 265.970 77.765 ;
        RECT 261.065 77.565 261.385 77.625 ;
        RECT 265.205 77.565 265.525 77.625 ;
        RECT 265.680 77.580 265.970 77.625 ;
        RECT 278.085 77.565 278.405 77.825 ;
        RECT 290.060 77.765 290.350 77.810 ;
        RECT 290.505 77.765 290.825 77.825 ;
        RECT 291.515 77.765 291.655 77.920 ;
        RECT 290.060 77.625 291.655 77.765 ;
        RECT 290.060 77.580 290.350 77.625 ;
        RECT 290.505 77.565 290.825 77.625 ;
        RECT 268.425 77.425 268.745 77.485 ;
        RECT 276.705 77.425 277.025 77.485 ;
        RECT 260.720 77.285 268.745 77.425 ;
        RECT 268.425 77.225 268.745 77.285 ;
        RECT 269.665 77.285 277.025 77.425 ;
        RECT 245.975 76.945 258.540 77.085 ;
        RECT 259.225 77.085 259.545 77.145 ;
        RECT 261.985 77.085 262.305 77.145 ;
        RECT 259.225 76.945 262.305 77.085 ;
        RECT 259.225 76.885 259.545 76.945 ;
        RECT 261.985 76.885 262.305 76.945 ;
        RECT 262.905 77.085 263.225 77.145 ;
        RECT 267.505 77.085 267.825 77.145 ;
        RECT 269.665 77.085 269.805 77.285 ;
        RECT 276.705 77.225 277.025 77.285 ;
        RECT 277.590 77.425 277.880 77.470 ;
        RECT 279.480 77.425 279.770 77.470 ;
        RECT 282.600 77.425 282.890 77.470 ;
        RECT 277.590 77.285 282.890 77.425 ;
        RECT 277.590 77.240 277.880 77.285 ;
        RECT 279.480 77.240 279.770 77.285 ;
        RECT 282.600 77.240 282.890 77.285 ;
        RECT 262.905 76.945 269.805 77.085 ;
        RECT 275.325 77.085 275.645 77.145 ;
        RECT 285.460 77.085 285.750 77.130 ;
        RECT 275.325 76.945 285.750 77.085 ;
        RECT 262.905 76.885 263.225 76.945 ;
        RECT 267.505 76.885 267.825 76.945 ;
        RECT 275.325 76.885 275.645 76.945 ;
        RECT 285.460 76.900 285.750 76.945 ;
        RECT 296.485 77.085 296.805 77.145 ;
        RECT 306.145 77.085 306.465 77.145 ;
        RECT 296.485 76.945 306.465 77.085 ;
        RECT 296.485 76.885 296.805 76.945 ;
        RECT 306.145 76.885 306.465 76.945 ;
        RECT 162.095 76.265 311.135 76.745 ;
        RECT 174.600 76.065 174.890 76.110 ;
        RECT 175.505 76.065 175.825 76.125 ;
        RECT 184.245 76.065 184.565 76.125 ;
        RECT 174.600 75.925 184.565 76.065 ;
        RECT 174.600 75.880 174.890 75.925 ;
        RECT 175.505 75.865 175.825 75.925 ;
        RECT 184.245 75.865 184.565 75.925 ;
        RECT 187.005 76.065 187.325 76.125 ;
        RECT 187.940 76.065 188.230 76.110 ;
        RECT 212.305 76.065 212.625 76.125 ;
        RECT 187.005 75.925 188.230 76.065 ;
        RECT 187.005 75.865 187.325 75.925 ;
        RECT 187.940 75.880 188.230 75.925 ;
        RECT 189.395 75.925 212.625 76.065 ;
        RECT 166.730 75.725 167.020 75.770 ;
        RECT 168.620 75.725 168.910 75.770 ;
        RECT 171.740 75.725 172.030 75.770 ;
        RECT 166.730 75.585 172.030 75.725 ;
        RECT 166.730 75.540 167.020 75.585 ;
        RECT 168.620 75.540 168.910 75.585 ;
        RECT 171.740 75.540 172.030 75.585 ;
        RECT 180.070 75.725 180.360 75.770 ;
        RECT 181.960 75.725 182.250 75.770 ;
        RECT 185.080 75.725 185.370 75.770 ;
        RECT 180.070 75.585 185.370 75.725 ;
        RECT 180.070 75.540 180.360 75.585 ;
        RECT 181.960 75.540 182.250 75.585 ;
        RECT 185.080 75.540 185.370 75.585 ;
        RECT 185.625 75.725 185.945 75.785 ;
        RECT 188.860 75.725 189.150 75.770 ;
        RECT 185.625 75.585 189.150 75.725 ;
        RECT 185.625 75.525 185.945 75.585 ;
        RECT 188.860 75.540 189.150 75.585 ;
        RECT 165.860 75.385 166.150 75.430 ;
        RECT 174.585 75.385 174.905 75.445 ;
        RECT 179.200 75.385 179.490 75.430 ;
        RECT 188.385 75.385 188.705 75.445 ;
        RECT 165.860 75.245 188.705 75.385 ;
        RECT 165.860 75.200 166.150 75.245 ;
        RECT 174.585 75.185 174.905 75.245 ;
        RECT 179.200 75.200 179.490 75.245 ;
        RECT 188.385 75.185 188.705 75.245 ;
        RECT 166.325 75.045 166.615 75.090 ;
        RECT 168.160 75.045 168.450 75.090 ;
        RECT 171.740 75.045 172.030 75.090 ;
        RECT 166.325 74.905 172.030 75.045 ;
        RECT 166.325 74.860 166.615 74.905 ;
        RECT 168.160 74.860 168.450 74.905 ;
        RECT 171.740 74.860 172.030 74.905 ;
        RECT 172.820 74.750 173.110 75.065 ;
        RECT 179.665 75.045 179.955 75.090 ;
        RECT 181.500 75.045 181.790 75.090 ;
        RECT 185.080 75.045 185.370 75.090 ;
        RECT 179.665 74.905 185.370 75.045 ;
        RECT 179.665 74.860 179.955 74.905 ;
        RECT 181.500 74.860 181.790 74.905 ;
        RECT 185.080 74.860 185.370 74.905 ;
        RECT 186.085 75.065 186.405 75.105 ;
        RECT 186.085 74.845 186.450 75.065 ;
        RECT 189.395 75.045 189.535 75.925 ;
        RECT 212.305 75.865 212.625 75.925 ;
        RECT 219.665 76.065 219.985 76.125 ;
        RECT 236.685 76.065 237.005 76.125 ;
        RECT 219.665 75.925 221.275 76.065 ;
        RECT 219.665 75.865 219.985 75.925 ;
        RECT 194.480 75.725 194.770 75.770 ;
        RECT 197.600 75.725 197.890 75.770 ;
        RECT 199.490 75.725 199.780 75.770 ;
        RECT 194.480 75.585 199.780 75.725 ;
        RECT 194.480 75.540 194.770 75.585 ;
        RECT 197.600 75.540 197.890 75.585 ;
        RECT 199.490 75.540 199.780 75.585 ;
        RECT 200.345 75.725 200.665 75.785 ;
        RECT 213.685 75.725 214.005 75.785 ;
        RECT 200.345 75.585 214.005 75.725 ;
        RECT 200.345 75.525 200.665 75.585 ;
        RECT 213.685 75.525 214.005 75.585 ;
        RECT 215.490 75.725 215.780 75.770 ;
        RECT 217.380 75.725 217.670 75.770 ;
        RECT 220.500 75.725 220.790 75.770 ;
        RECT 215.490 75.585 220.790 75.725 ;
        RECT 221.135 75.725 221.275 75.925 ;
        RECT 223.435 75.925 237.005 76.065 ;
        RECT 223.435 75.770 223.575 75.925 ;
        RECT 236.685 75.865 237.005 75.925 ;
        RECT 238.080 76.065 238.370 76.110 ;
        RECT 241.285 76.065 241.605 76.125 ;
        RECT 238.080 75.925 241.605 76.065 ;
        RECT 238.080 75.880 238.370 75.925 ;
        RECT 241.285 75.865 241.605 75.925 ;
        RECT 255.085 76.065 255.405 76.125 ;
        RECT 258.305 76.065 258.625 76.125 ;
        RECT 255.085 75.925 258.625 76.065 ;
        RECT 255.085 75.865 255.405 75.925 ;
        RECT 258.305 75.865 258.625 75.925 ;
        RECT 258.765 76.065 259.085 76.125 ;
        RECT 262.445 76.065 262.765 76.125 ;
        RECT 258.765 75.925 262.765 76.065 ;
        RECT 258.765 75.865 259.085 75.925 ;
        RECT 262.445 75.865 262.765 75.925 ;
        RECT 277.640 76.065 277.930 76.110 ;
        RECT 278.085 76.065 278.405 76.125 ;
        RECT 277.640 75.925 278.405 76.065 ;
        RECT 277.640 75.880 277.930 75.925 ;
        RECT 278.085 75.865 278.405 75.925 ;
        RECT 282.685 76.065 283.005 76.125 ;
        RECT 287.760 76.065 288.050 76.110 ;
        RECT 282.685 75.925 288.050 76.065 ;
        RECT 282.685 75.865 283.005 75.925 ;
        RECT 287.760 75.880 288.050 75.925 ;
        RECT 294.200 76.065 294.490 76.110 ;
        RECT 295.565 76.065 295.885 76.125 ;
        RECT 304.765 76.065 305.085 76.125 ;
        RECT 294.200 75.925 295.885 76.065 ;
        RECT 294.200 75.880 294.490 75.925 ;
        RECT 295.565 75.865 295.885 75.925 ;
        RECT 296.115 75.925 305.085 76.065 ;
        RECT 223.360 75.725 223.650 75.770 ;
        RECT 221.135 75.585 223.650 75.725 ;
        RECT 215.490 75.540 215.780 75.585 ;
        RECT 217.380 75.540 217.670 75.585 ;
        RECT 220.500 75.540 220.790 75.585 ;
        RECT 223.360 75.540 223.650 75.585 ;
        RECT 224.280 75.540 224.570 75.770 ;
        RECT 229.325 75.725 229.645 75.785 ;
        RECT 254.625 75.725 254.945 75.785 ;
        RECT 259.685 75.725 260.005 75.785 ;
        RECT 270.265 75.725 270.585 75.785 ;
        RECT 229.325 75.585 254.945 75.725 ;
        RECT 190.685 75.185 191.005 75.445 ;
        RECT 191.620 75.385 191.910 75.430 ;
        RECT 203.580 75.385 203.870 75.430 ;
        RECT 204.025 75.385 204.345 75.445 ;
        RECT 191.620 75.245 204.345 75.385 ;
        RECT 191.620 75.200 191.910 75.245 ;
        RECT 203.580 75.200 203.870 75.245 ;
        RECT 204.025 75.185 204.345 75.245 ;
        RECT 204.500 75.385 204.790 75.430 ;
        RECT 206.785 75.385 207.105 75.445 ;
        RECT 211.400 75.385 211.690 75.430 ;
        RECT 211.845 75.385 212.165 75.445 ;
        RECT 204.500 75.245 212.165 75.385 ;
        RECT 204.500 75.200 204.790 75.245 ;
        RECT 206.785 75.185 207.105 75.245 ;
        RECT 211.400 75.200 211.690 75.245 ;
        RECT 211.845 75.185 212.165 75.245 ;
        RECT 215.985 75.185 216.305 75.445 ;
        RECT 218.285 75.385 218.605 75.445 ;
        RECT 224.355 75.385 224.495 75.540 ;
        RECT 229.325 75.525 229.645 75.585 ;
        RECT 254.625 75.525 254.945 75.585 ;
        RECT 257.475 75.585 258.540 75.725 ;
        RECT 257.475 75.445 257.615 75.585 ;
        RECT 218.285 75.245 224.495 75.385 ;
        RECT 237.145 75.385 237.465 75.445 ;
        RECT 255.085 75.385 255.405 75.445 ;
        RECT 237.145 75.245 255.405 75.385 ;
        RECT 218.285 75.185 218.605 75.245 ;
        RECT 167.240 74.520 167.530 74.750 ;
        RECT 169.520 74.705 170.170 74.750 ;
        RECT 172.820 74.705 173.410 74.750 ;
        RECT 169.520 74.565 174.815 74.705 ;
        RECT 169.520 74.520 170.170 74.565 ;
        RECT 173.120 74.520 173.410 74.565 ;
        RECT 167.315 74.365 167.455 74.520 ;
        RECT 174.125 74.365 174.445 74.425 ;
        RECT 167.315 74.225 174.445 74.365 ;
        RECT 174.675 74.365 174.815 74.565 ;
        RECT 180.565 74.505 180.885 74.765 ;
        RECT 186.160 74.750 186.450 74.845 ;
        RECT 187.095 74.905 189.535 75.045 ;
        RECT 190.240 75.045 190.530 75.090 ;
        RECT 191.145 75.045 191.465 75.105 ;
        RECT 190.240 74.905 191.465 75.045 ;
        RECT 182.860 74.705 183.510 74.750 ;
        RECT 186.160 74.705 186.750 74.750 ;
        RECT 182.860 74.565 186.750 74.705 ;
        RECT 182.860 74.520 183.510 74.565 ;
        RECT 186.460 74.520 186.750 74.565 ;
        RECT 175.045 74.365 175.365 74.425 ;
        RECT 181.945 74.365 182.265 74.425 ;
        RECT 174.675 74.225 182.265 74.365 ;
        RECT 174.125 74.165 174.445 74.225 ;
        RECT 175.045 74.165 175.365 74.225 ;
        RECT 181.945 74.165 182.265 74.225 ;
        RECT 182.405 74.365 182.725 74.425 ;
        RECT 184.705 74.365 185.025 74.425 ;
        RECT 187.095 74.365 187.235 74.905 ;
        RECT 190.240 74.860 190.530 74.905 ;
        RECT 188.400 74.520 188.690 74.750 ;
        RECT 189.305 74.705 189.625 74.765 ;
        RECT 190.315 74.705 190.455 74.860 ;
        RECT 191.145 74.845 191.465 74.905 ;
        RECT 189.305 74.565 190.455 74.705 ;
        RECT 192.525 74.705 192.845 74.765 ;
        RECT 193.400 74.750 193.690 75.065 ;
        RECT 194.480 75.045 194.770 75.090 ;
        RECT 198.060 75.045 198.350 75.090 ;
        RECT 199.895 75.045 200.185 75.090 ;
        RECT 194.480 74.905 200.185 75.045 ;
        RECT 194.480 74.860 194.770 74.905 ;
        RECT 198.060 74.860 198.350 74.905 ;
        RECT 199.895 74.860 200.185 74.905 ;
        RECT 200.360 75.045 200.650 75.090 ;
        RECT 210.465 75.045 210.785 75.105 ;
        RECT 214.145 75.045 214.465 75.105 ;
        RECT 214.620 75.045 214.910 75.090 ;
        RECT 200.360 74.905 214.910 75.045 ;
        RECT 200.360 74.860 200.650 74.905 ;
        RECT 210.465 74.845 210.785 74.905 ;
        RECT 214.145 74.845 214.465 74.905 ;
        RECT 214.620 74.860 214.910 74.905 ;
        RECT 215.085 75.045 215.375 75.090 ;
        RECT 216.920 75.045 217.210 75.090 ;
        RECT 220.500 75.045 220.790 75.090 ;
        RECT 215.085 74.905 220.790 75.045 ;
        RECT 215.085 74.860 215.375 74.905 ;
        RECT 216.920 74.860 217.210 74.905 ;
        RECT 220.500 74.860 220.790 74.905 ;
        RECT 193.100 74.705 193.690 74.750 ;
        RECT 196.340 74.705 196.990 74.750 ;
        RECT 192.525 74.565 196.990 74.705 ;
        RECT 182.405 74.225 187.235 74.365 ;
        RECT 188.475 74.365 188.615 74.520 ;
        RECT 189.305 74.505 189.625 74.565 ;
        RECT 192.525 74.505 192.845 74.565 ;
        RECT 193.100 74.520 193.390 74.565 ;
        RECT 196.340 74.520 196.990 74.565 ;
        RECT 198.980 74.520 199.270 74.750 ;
        RECT 200.805 74.705 201.125 74.765 ;
        RECT 205.420 74.705 205.710 74.750 ;
        RECT 200.805 74.565 205.710 74.705 ;
        RECT 191.145 74.365 191.465 74.425 ;
        RECT 188.475 74.225 191.465 74.365 ;
        RECT 199.055 74.365 199.195 74.520 ;
        RECT 200.805 74.505 201.125 74.565 ;
        RECT 205.420 74.520 205.710 74.565 ;
        RECT 207.260 74.520 207.550 74.750 ;
        RECT 201.280 74.365 201.570 74.410 ;
        RECT 199.055 74.225 201.570 74.365 ;
        RECT 182.405 74.165 182.725 74.225 ;
        RECT 184.705 74.165 185.025 74.225 ;
        RECT 191.145 74.165 191.465 74.225 ;
        RECT 201.280 74.180 201.570 74.225 ;
        RECT 203.105 74.165 203.425 74.425 ;
        RECT 207.335 74.365 207.475 74.520 ;
        RECT 211.845 74.505 212.165 74.765 ;
        RECT 212.305 74.505 212.625 74.765 ;
        RECT 218.285 74.750 218.605 74.765 ;
        RECT 221.580 74.750 221.870 75.065 ;
        RECT 222.055 74.750 222.195 75.245 ;
        RECT 237.145 75.185 237.465 75.245 ;
        RECT 255.085 75.185 255.405 75.245 ;
        RECT 257.385 75.185 257.705 75.445 ;
        RECT 258.400 75.385 258.540 75.585 ;
        RECT 259.685 75.585 270.585 75.725 ;
        RECT 259.685 75.525 260.005 75.585 ;
        RECT 270.265 75.525 270.585 75.585 ;
        RECT 279.890 75.725 280.180 75.770 ;
        RECT 281.780 75.725 282.070 75.770 ;
        RECT 284.900 75.725 285.190 75.770 ;
        RECT 279.890 75.585 285.190 75.725 ;
        RECT 279.890 75.540 280.180 75.585 ;
        RECT 281.780 75.540 282.070 75.585 ;
        RECT 284.900 75.540 285.190 75.585 ;
        RECT 285.445 75.725 285.765 75.785 ;
        RECT 294.660 75.725 294.950 75.770 ;
        RECT 296.115 75.725 296.255 75.925 ;
        RECT 304.765 75.865 305.085 75.925 ;
        RECT 285.445 75.585 296.255 75.725 ;
        RECT 297.520 75.725 297.810 75.770 ;
        RECT 300.640 75.725 300.930 75.770 ;
        RECT 302.530 75.725 302.820 75.770 ;
        RECT 297.520 75.585 302.820 75.725 ;
        RECT 285.445 75.525 285.765 75.585 ;
        RECT 294.660 75.540 294.950 75.585 ;
        RECT 297.520 75.540 297.810 75.585 ;
        RECT 300.640 75.540 300.930 75.585 ;
        RECT 302.530 75.540 302.820 75.585 ;
        RECT 264.285 75.385 264.605 75.445 ;
        RECT 258.400 75.245 259.915 75.385 ;
        RECT 225.185 74.845 225.505 75.105 ;
        RECT 237.605 74.845 237.925 75.105 ;
        RECT 238.080 74.860 238.370 75.090 ;
        RECT 218.280 74.705 218.930 74.750 ;
        RECT 221.580 74.705 222.195 74.750 ;
        RECT 222.885 74.705 223.205 74.765 ;
        RECT 213.775 74.565 223.205 74.705 ;
        RECT 213.775 74.365 213.915 74.565 ;
        RECT 218.280 74.520 218.930 74.565 ;
        RECT 221.880 74.520 222.170 74.565 ;
        RECT 218.285 74.505 218.605 74.520 ;
        RECT 222.885 74.505 223.205 74.565 ;
        RECT 232.545 74.705 232.865 74.765 ;
        RECT 238.155 74.705 238.295 74.860 ;
        RECT 257.845 74.845 258.165 75.105 ;
        RECT 259.775 75.090 259.915 75.245 ;
        RECT 261.155 75.245 264.605 75.385 ;
        RECT 258.325 74.860 258.615 75.090 ;
        RECT 259.240 74.860 259.530 75.090 ;
        RECT 259.700 74.860 259.990 75.090 ;
        RECT 260.390 75.045 260.680 75.090 ;
        RECT 261.155 75.045 261.295 75.245 ;
        RECT 264.285 75.185 264.605 75.245 ;
        RECT 274.880 75.385 275.170 75.430 ;
        RECT 276.705 75.385 277.025 75.445 ;
        RECT 274.880 75.245 277.025 75.385 ;
        RECT 274.880 75.200 275.170 75.245 ;
        RECT 276.705 75.185 277.025 75.245 ;
        RECT 280.385 75.185 280.705 75.445 ;
        RECT 280.845 75.385 281.165 75.445 ;
        RECT 290.965 75.385 291.285 75.445 ;
        RECT 296.025 75.385 296.345 75.445 ;
        RECT 280.845 75.245 286.595 75.385 ;
        RECT 280.845 75.185 281.165 75.245 ;
        RECT 260.390 74.905 261.295 75.045 ;
        RECT 260.390 74.860 260.680 74.905 ;
        RECT 232.545 74.565 238.295 74.705 ;
        RECT 257.385 74.705 257.705 74.765 ;
        RECT 258.400 74.705 258.540 74.860 ;
        RECT 257.385 74.565 258.540 74.705 ;
        RECT 259.315 74.705 259.455 74.860 ;
        RECT 261.525 74.845 261.845 75.105 ;
        RECT 261.985 74.845 262.305 75.105 ;
        RECT 262.445 74.845 262.765 75.105 ;
        RECT 262.905 74.845 263.225 75.105 ;
        RECT 263.380 75.045 263.670 75.090 ;
        RECT 265.665 75.045 265.985 75.105 ;
        RECT 263.380 74.905 265.985 75.045 ;
        RECT 263.380 74.860 263.670 74.905 ;
        RECT 265.665 74.845 265.985 74.905 ;
        RECT 268.425 75.045 268.745 75.105 ;
        RECT 275.800 75.045 276.090 75.090 ;
        RECT 268.425 74.905 276.090 75.045 ;
        RECT 268.425 74.845 268.745 74.905 ;
        RECT 275.800 74.860 276.090 74.905 ;
        RECT 278.545 75.045 278.865 75.105 ;
        RECT 279.020 75.045 279.310 75.090 ;
        RECT 278.545 74.905 279.310 75.045 ;
        RECT 262.075 74.705 262.215 74.845 ;
        RECT 259.315 74.565 262.215 74.705 ;
        RECT 270.725 74.705 271.045 74.765 ;
        RECT 275.325 74.705 275.645 74.765 ;
        RECT 270.725 74.565 275.645 74.705 ;
        RECT 275.875 74.705 276.015 74.860 ;
        RECT 278.545 74.845 278.865 74.905 ;
        RECT 279.020 74.860 279.310 74.905 ;
        RECT 279.485 75.045 279.775 75.090 ;
        RECT 281.320 75.045 281.610 75.090 ;
        RECT 284.900 75.045 285.190 75.090 ;
        RECT 279.485 74.905 285.190 75.045 ;
        RECT 279.485 74.860 279.775 74.905 ;
        RECT 281.320 74.860 281.610 74.905 ;
        RECT 284.900 74.860 285.190 74.905 ;
        RECT 280.845 74.705 281.165 74.765 ;
        RECT 285.980 74.750 286.270 75.065 ;
        RECT 286.455 75.045 286.595 75.245 ;
        RECT 290.965 75.245 296.345 75.385 ;
        RECT 290.965 75.185 291.285 75.245 ;
        RECT 296.025 75.185 296.345 75.245 ;
        RECT 296.945 75.385 297.265 75.445 ;
        RECT 303.400 75.385 303.690 75.430 ;
        RECT 296.945 75.245 303.690 75.385 ;
        RECT 296.945 75.185 297.265 75.245 ;
        RECT 303.400 75.200 303.690 75.245 ;
        RECT 292.360 75.045 292.650 75.090 ;
        RECT 286.455 74.905 292.650 75.045 ;
        RECT 292.360 74.860 292.650 74.905 ;
        RECT 275.875 74.565 281.165 74.705 ;
        RECT 232.545 74.505 232.865 74.565 ;
        RECT 257.385 74.505 257.705 74.565 ;
        RECT 207.335 74.225 213.915 74.365 ;
        RECT 214.160 74.365 214.450 74.410 ;
        RECT 215.525 74.365 215.845 74.425 ;
        RECT 214.160 74.225 215.845 74.365 ;
        RECT 214.160 74.180 214.450 74.225 ;
        RECT 215.525 74.165 215.845 74.225 ;
        RECT 220.125 74.365 220.445 74.425 ;
        RECT 231.165 74.365 231.485 74.425 ;
        RECT 220.125 74.225 231.485 74.365 ;
        RECT 220.125 74.165 220.445 74.225 ;
        RECT 231.165 74.165 231.485 74.225 ;
        RECT 236.225 74.165 236.545 74.425 ;
        RECT 238.985 74.365 239.305 74.425 ;
        RECT 245.885 74.365 246.205 74.425 ;
        RECT 238.985 74.225 246.205 74.365 ;
        RECT 238.985 74.165 239.305 74.225 ;
        RECT 245.885 74.165 246.205 74.225 ;
        RECT 256.925 74.365 257.245 74.425 ;
        RECT 259.315 74.365 259.455 74.565 ;
        RECT 270.725 74.505 271.045 74.565 ;
        RECT 275.325 74.505 275.645 74.565 ;
        RECT 280.845 74.505 281.165 74.565 ;
        RECT 282.680 74.705 283.330 74.750 ;
        RECT 285.980 74.705 286.570 74.750 ;
        RECT 286.825 74.705 287.145 74.765 ;
        RECT 296.440 74.750 296.730 75.065 ;
        RECT 297.520 75.045 297.810 75.090 ;
        RECT 301.100 75.045 301.390 75.090 ;
        RECT 302.935 75.045 303.225 75.090 ;
        RECT 297.520 74.905 303.225 75.045 ;
        RECT 297.520 74.860 297.810 74.905 ;
        RECT 301.100 74.860 301.390 74.905 ;
        RECT 302.935 74.860 303.225 74.905 ;
        RECT 296.140 74.705 296.730 74.750 ;
        RECT 299.380 74.705 300.030 74.750 ;
        RECT 302.020 74.705 302.310 74.750 ;
        RECT 304.305 74.705 304.625 74.765 ;
        RECT 282.680 74.565 295.335 74.705 ;
        RECT 282.680 74.520 283.330 74.565 ;
        RECT 286.280 74.520 286.570 74.565 ;
        RECT 286.825 74.505 287.145 74.565 ;
        RECT 256.925 74.225 259.455 74.365 ;
        RECT 261.080 74.365 261.370 74.410 ;
        RECT 263.365 74.365 263.685 74.425 ;
        RECT 261.080 74.225 263.685 74.365 ;
        RECT 256.925 74.165 257.245 74.225 ;
        RECT 261.080 74.180 261.370 74.225 ;
        RECT 263.365 74.165 263.685 74.225 ;
        RECT 264.300 74.365 264.590 74.410 ;
        RECT 265.205 74.365 265.525 74.425 ;
        RECT 264.300 74.225 265.525 74.365 ;
        RECT 264.300 74.180 264.590 74.225 ;
        RECT 265.205 74.165 265.525 74.225 ;
        RECT 270.265 74.365 270.585 74.425 ;
        RECT 271.645 74.365 271.965 74.425 ;
        RECT 270.265 74.225 271.965 74.365 ;
        RECT 270.265 74.165 270.585 74.225 ;
        RECT 271.645 74.165 271.965 74.225 ;
        RECT 272.105 74.365 272.425 74.425 ;
        RECT 285.445 74.365 285.765 74.425 ;
        RECT 272.105 74.225 285.765 74.365 ;
        RECT 272.105 74.165 272.425 74.225 ;
        RECT 285.445 74.165 285.765 74.225 ;
        RECT 291.885 74.165 292.205 74.425 ;
        RECT 295.195 74.365 295.335 74.565 ;
        RECT 296.140 74.565 300.395 74.705 ;
        RECT 296.140 74.520 296.430 74.565 ;
        RECT 299.380 74.520 300.030 74.565 ;
        RECT 300.255 74.365 300.395 74.565 ;
        RECT 302.020 74.565 304.625 74.705 ;
        RECT 302.020 74.520 302.310 74.565 ;
        RECT 304.305 74.505 304.625 74.565 ;
        RECT 303.845 74.365 304.165 74.425 ;
        RECT 295.195 74.225 304.165 74.365 ;
        RECT 303.845 74.165 304.165 74.225 ;
        RECT 162.095 73.545 311.135 74.025 ;
        RECT 174.125 73.345 174.445 73.405 ;
        RECT 177.820 73.345 178.110 73.390 ;
        RECT 174.125 73.205 178.110 73.345 ;
        RECT 174.125 73.145 174.445 73.205 ;
        RECT 177.820 73.160 178.110 73.205 ;
        RECT 180.565 73.345 180.885 73.405 ;
        RECT 182.880 73.345 183.170 73.390 ;
        RECT 180.565 73.205 183.170 73.345 ;
        RECT 180.565 73.145 180.885 73.205 ;
        RECT 182.880 73.160 183.170 73.205 ;
        RECT 185.180 73.345 185.470 73.390 ;
        RECT 186.545 73.345 186.865 73.405 ;
        RECT 185.180 73.205 186.865 73.345 ;
        RECT 185.180 73.160 185.470 73.205 ;
        RECT 186.545 73.145 186.865 73.205 ;
        RECT 202.185 73.345 202.505 73.405 ;
        RECT 202.185 73.205 232.315 73.345 ;
        RECT 202.185 73.145 202.505 73.205 ;
        RECT 170.100 73.005 170.390 73.050 ;
        RECT 172.745 73.005 173.065 73.065 ;
        RECT 173.340 73.005 173.990 73.050 ;
        RECT 170.100 72.865 173.990 73.005 ;
        RECT 170.100 72.820 170.690 72.865 ;
        RECT 170.400 72.505 170.690 72.820 ;
        RECT 172.745 72.805 173.065 72.865 ;
        RECT 173.340 72.820 173.990 72.865 ;
        RECT 175.965 72.805 176.285 73.065 ;
        RECT 192.525 73.005 192.845 73.065 ;
        RECT 200.805 73.050 201.125 73.065 ;
        RECT 200.800 73.005 201.450 73.050 ;
        RECT 204.400 73.005 204.690 73.050 ;
        RECT 177.435 72.865 192.295 73.005 ;
        RECT 177.435 72.725 177.575 72.865 ;
        RECT 171.480 72.665 171.770 72.710 ;
        RECT 175.060 72.665 175.350 72.710 ;
        RECT 176.895 72.665 177.185 72.710 ;
        RECT 171.480 72.525 177.185 72.665 ;
        RECT 171.480 72.480 171.770 72.525 ;
        RECT 175.060 72.480 175.350 72.525 ;
        RECT 176.895 72.480 177.185 72.525 ;
        RECT 177.345 72.465 177.665 72.725 ;
        RECT 179.185 72.665 179.505 72.725 ;
        RECT 179.660 72.665 179.950 72.710 ;
        RECT 179.185 72.525 179.950 72.665 ;
        RECT 179.185 72.465 179.505 72.525 ;
        RECT 179.660 72.480 179.950 72.525 ;
        RECT 184.705 72.465 185.025 72.725 ;
        RECT 188.400 72.665 188.690 72.710 ;
        RECT 190.225 72.665 190.545 72.725 ;
        RECT 192.155 72.710 192.295 72.865 ;
        RECT 192.525 72.865 204.690 73.005 ;
        RECT 192.525 72.805 192.845 72.865 ;
        RECT 200.800 72.820 201.450 72.865 ;
        RECT 204.100 72.820 204.690 72.865 ;
        RECT 200.805 72.805 201.125 72.820 ;
        RECT 188.400 72.525 190.545 72.665 ;
        RECT 188.400 72.480 188.690 72.525 ;
        RECT 190.225 72.465 190.545 72.525 ;
        RECT 192.080 72.665 192.370 72.710 ;
        RECT 193.460 72.665 193.750 72.710 ;
        RECT 192.080 72.525 193.750 72.665 ;
        RECT 192.080 72.480 192.370 72.525 ;
        RECT 193.460 72.480 193.750 72.525 ;
        RECT 197.605 72.665 197.895 72.710 ;
        RECT 199.440 72.665 199.730 72.710 ;
        RECT 203.020 72.665 203.310 72.710 ;
        RECT 197.605 72.525 203.310 72.665 ;
        RECT 197.605 72.480 197.895 72.525 ;
        RECT 199.440 72.480 199.730 72.525 ;
        RECT 203.020 72.480 203.310 72.525 ;
        RECT 204.100 72.505 204.390 72.820 ;
        RECT 206.785 72.805 207.105 73.065 ;
        RECT 215.525 72.805 215.845 73.065 ;
        RECT 217.820 73.005 218.470 73.050 ;
        RECT 221.420 73.005 221.710 73.050 ;
        RECT 222.885 73.005 223.205 73.065 ;
        RECT 217.820 72.865 223.205 73.005 ;
        RECT 217.820 72.820 218.470 72.865 ;
        RECT 221.120 72.820 221.710 72.865 ;
        RECT 206.340 72.665 206.630 72.710 ;
        RECT 207.705 72.665 208.025 72.725 ;
        RECT 208.180 72.665 208.470 72.710 ;
        RECT 206.340 72.525 207.015 72.665 ;
        RECT 206.340 72.480 206.630 72.525 ;
        RECT 168.620 72.325 168.910 72.370 ;
        RECT 173.665 72.325 173.985 72.385 ;
        RECT 168.620 72.185 173.985 72.325 ;
        RECT 168.620 72.140 168.910 72.185 ;
        RECT 173.665 72.125 173.985 72.185 ;
        RECT 175.505 72.325 175.825 72.385 ;
        RECT 180.120 72.325 180.410 72.370 ;
        RECT 175.505 72.185 180.410 72.325 ;
        RECT 175.505 72.125 175.825 72.185 ;
        RECT 179.735 72.045 179.875 72.185 ;
        RECT 180.120 72.140 180.410 72.185 ;
        RECT 180.565 72.325 180.885 72.385 ;
        RECT 181.040 72.325 181.330 72.370 ;
        RECT 185.625 72.325 185.945 72.385 ;
        RECT 180.565 72.185 185.945 72.325 ;
        RECT 180.565 72.125 180.885 72.185 ;
        RECT 181.040 72.140 181.330 72.185 ;
        RECT 185.625 72.125 185.945 72.185 ;
        RECT 192.525 72.325 192.845 72.385 ;
        RECT 197.140 72.325 197.430 72.370 ;
        RECT 192.525 72.185 197.430 72.325 ;
        RECT 192.525 72.125 192.845 72.185 ;
        RECT 197.140 72.140 197.430 72.185 ;
        RECT 198.520 72.325 198.810 72.370 ;
        RECT 201.265 72.325 201.585 72.385 ;
        RECT 198.520 72.185 201.585 72.325 ;
        RECT 198.520 72.140 198.810 72.185 ;
        RECT 201.265 72.125 201.585 72.185 ;
        RECT 171.480 71.985 171.770 72.030 ;
        RECT 174.600 71.985 174.890 72.030 ;
        RECT 176.490 71.985 176.780 72.030 ;
        RECT 171.480 71.845 176.780 71.985 ;
        RECT 171.480 71.800 171.770 71.845 ;
        RECT 174.600 71.800 174.890 71.845 ;
        RECT 176.490 71.800 176.780 71.845 ;
        RECT 179.645 71.785 179.965 72.045 ;
        RECT 198.010 71.985 198.300 72.030 ;
        RECT 199.900 71.985 200.190 72.030 ;
        RECT 203.020 71.985 203.310 72.030 ;
        RECT 206.875 71.985 207.015 72.525 ;
        RECT 207.705 72.525 208.470 72.665 ;
        RECT 207.705 72.465 208.025 72.525 ;
        RECT 208.180 72.480 208.470 72.525 ;
        RECT 214.145 72.465 214.465 72.725 ;
        RECT 214.625 72.665 214.915 72.710 ;
        RECT 216.460 72.665 216.750 72.710 ;
        RECT 220.040 72.665 220.330 72.710 ;
        RECT 214.625 72.525 220.330 72.665 ;
        RECT 214.625 72.480 214.915 72.525 ;
        RECT 216.460 72.480 216.750 72.525 ;
        RECT 220.040 72.480 220.330 72.525 ;
        RECT 221.120 72.505 221.410 72.820 ;
        RECT 222.885 72.805 223.205 72.865 ;
        RECT 228.865 73.005 229.185 73.065 ;
        RECT 231.180 73.005 231.470 73.050 ;
        RECT 228.865 72.865 231.470 73.005 ;
        RECT 232.175 73.005 232.315 73.205 ;
        RECT 232.545 73.145 232.865 73.405 ;
        RECT 237.605 73.345 237.925 73.405 ;
        RECT 239.000 73.345 239.290 73.390 ;
        RECT 237.605 73.205 239.290 73.345 ;
        RECT 237.605 73.145 237.925 73.205 ;
        RECT 239.000 73.160 239.290 73.205 ;
        RECT 241.285 73.145 241.605 73.405 ;
        RECT 244.965 73.345 245.285 73.405 ;
        RECT 242.755 73.205 245.285 73.345 ;
        RECT 237.145 73.005 237.465 73.065 ;
        RECT 242.755 73.050 242.895 73.205 ;
        RECT 244.965 73.145 245.285 73.205 ;
        RECT 245.885 73.345 246.205 73.405 ;
        RECT 257.845 73.345 258.165 73.405 ;
        RECT 261.525 73.345 261.845 73.405 ;
        RECT 265.665 73.345 265.985 73.405 ;
        RECT 245.885 73.205 258.165 73.345 ;
        RECT 245.885 73.145 246.205 73.205 ;
        RECT 257.845 73.145 258.165 73.205 ;
        RECT 258.400 73.205 260.375 73.345 ;
        RECT 232.175 72.865 237.465 73.005 ;
        RECT 228.865 72.805 229.185 72.865 ;
        RECT 231.180 72.820 231.470 72.865 ;
        RECT 237.145 72.805 237.465 72.865 ;
        RECT 242.680 72.820 242.970 73.050 ;
        RECT 251.865 73.005 252.185 73.065 ;
        RECT 258.400 73.005 258.540 73.205 ;
        RECT 243.650 72.865 258.540 73.005 ;
        RECT 258.765 73.005 259.085 73.065 ;
        RECT 259.240 73.005 259.530 73.050 ;
        RECT 258.765 72.865 259.530 73.005 ;
        RECT 229.785 72.465 230.105 72.725 ;
        RECT 230.705 72.465 231.025 72.725 ;
        RECT 231.640 72.665 231.930 72.710 ;
        RECT 232.085 72.665 232.405 72.725 ;
        RECT 231.640 72.525 232.405 72.665 ;
        RECT 231.640 72.480 231.930 72.525 ;
        RECT 232.085 72.465 232.405 72.525 ;
        RECT 233.465 72.665 233.785 72.725 ;
        RECT 236.685 72.710 237.005 72.725 ;
        RECT 235.780 72.665 236.070 72.710 ;
        RECT 233.465 72.525 236.070 72.665 ;
        RECT 233.465 72.465 233.785 72.525 ;
        RECT 235.780 72.480 236.070 72.525 ;
        RECT 236.520 72.480 237.005 72.710 ;
        RECT 236.685 72.465 237.005 72.480 ;
        RECT 237.605 72.465 237.925 72.725 ;
        RECT 238.310 72.665 238.600 72.710 ;
        RECT 241.285 72.665 241.605 72.725 ;
        RECT 242.205 72.710 242.525 72.725 ;
        RECT 242.195 72.665 242.525 72.710 ;
        RECT 238.310 72.525 241.605 72.665 ;
        RECT 242.010 72.525 242.525 72.665 ;
        RECT 238.310 72.480 238.600 72.525 ;
        RECT 241.285 72.465 241.605 72.525 ;
        RECT 242.195 72.480 242.525 72.525 ;
        RECT 243.140 72.665 243.430 72.710 ;
        RECT 243.650 72.665 243.790 72.865 ;
        RECT 251.865 72.805 252.185 72.865 ;
        RECT 258.765 72.805 259.085 72.865 ;
        RECT 259.240 72.820 259.530 72.865 ;
        RECT 243.140 72.525 243.790 72.665 ;
        RECT 243.140 72.480 243.430 72.525 ;
        RECT 242.205 72.465 242.525 72.480 ;
        RECT 244.040 72.465 244.360 72.725 ;
        RECT 244.575 72.665 244.865 72.710 ;
        RECT 245.885 72.665 246.205 72.725 ;
        RECT 256.005 72.665 256.325 72.725 ;
        RECT 258.320 72.665 258.610 72.710 ;
        RECT 244.575 72.525 246.205 72.665 ;
        RECT 244.575 72.480 244.865 72.525 ;
        RECT 245.885 72.465 246.205 72.525 ;
        RECT 255.865 72.525 258.610 72.665 ;
        RECT 255.865 72.465 256.325 72.525 ;
        RECT 258.320 72.480 258.610 72.525 ;
        RECT 209.100 72.325 209.390 72.370 ;
        RECT 211.385 72.325 211.705 72.385 ;
        RECT 209.100 72.185 211.705 72.325 ;
        RECT 209.100 72.140 209.390 72.185 ;
        RECT 211.385 72.125 211.705 72.185 ;
        RECT 212.305 72.325 212.625 72.385 ;
        RECT 215.525 72.325 215.845 72.385 ;
        RECT 222.900 72.325 223.190 72.370 ;
        RECT 255.865 72.325 256.005 72.465 ;
        RECT 212.305 72.185 256.005 72.325 ;
        RECT 212.305 72.125 212.625 72.185 ;
        RECT 215.525 72.125 215.845 72.185 ;
        RECT 222.900 72.140 223.190 72.185 ;
        RECT 207.705 71.985 208.025 72.045 ;
        RECT 198.010 71.845 203.310 71.985 ;
        RECT 198.010 71.800 198.300 71.845 ;
        RECT 199.900 71.800 200.190 71.845 ;
        RECT 203.020 71.800 203.310 71.845 ;
        RECT 203.655 71.845 208.025 71.985 ;
        RECT 175.965 71.645 176.285 71.705 ;
        RECT 179.185 71.645 179.505 71.705 ;
        RECT 175.965 71.505 179.505 71.645 ;
        RECT 175.965 71.445 176.285 71.505 ;
        RECT 179.185 71.445 179.505 71.505 ;
        RECT 191.145 71.645 191.465 71.705 ;
        RECT 203.655 71.645 203.795 71.845 ;
        RECT 207.705 71.785 208.025 71.845 ;
        RECT 215.030 71.985 215.320 72.030 ;
        RECT 216.920 71.985 217.210 72.030 ;
        RECT 220.040 71.985 220.330 72.030 ;
        RECT 230.705 71.985 231.025 72.045 ;
        RECT 215.030 71.845 220.330 71.985 ;
        RECT 215.030 71.800 215.320 71.845 ;
        RECT 216.920 71.800 217.210 71.845 ;
        RECT 220.040 71.800 220.330 71.845 ;
        RECT 225.275 71.845 231.025 71.985 ;
        RECT 191.145 71.505 203.795 71.645 ;
        RECT 191.145 71.445 191.465 71.505 ;
        RECT 205.865 71.445 206.185 71.705 ;
        RECT 206.325 71.645 206.645 71.705 ;
        RECT 225.275 71.645 225.415 71.845 ;
        RECT 230.705 71.785 231.025 71.845 ;
        RECT 256.005 71.985 256.325 72.045 ;
        RECT 256.925 71.985 257.245 72.045 ;
        RECT 256.005 71.845 257.245 71.985 ;
        RECT 256.005 71.785 256.325 71.845 ;
        RECT 256.925 71.785 257.245 71.845 ;
        RECT 206.325 71.505 225.415 71.645 ;
        RECT 237.145 71.645 237.465 71.705 ;
        RECT 247.265 71.645 247.585 71.705 ;
        RECT 258.855 71.645 258.995 72.805 ;
        RECT 260.235 72.710 260.375 73.205 ;
        RECT 261.525 73.205 265.985 73.345 ;
        RECT 261.525 73.145 261.845 73.205 ;
        RECT 259.700 72.480 259.990 72.710 ;
        RECT 260.160 72.665 260.450 72.710 ;
        RECT 260.605 72.665 260.925 72.725 ;
        RECT 260.160 72.525 260.925 72.665 ;
        RECT 260.160 72.480 260.450 72.525 ;
        RECT 259.775 72.325 259.915 72.480 ;
        RECT 260.605 72.465 260.925 72.525 ;
        RECT 262.445 72.465 262.765 72.725 ;
        RECT 262.920 72.480 263.210 72.710 ;
        RECT 263.380 72.665 263.670 72.710 ;
        RECT 263.915 72.665 264.055 73.205 ;
        RECT 265.665 73.145 265.985 73.205 ;
        RECT 267.965 73.345 268.285 73.405 ;
        RECT 277.625 73.345 277.945 73.405 ;
        RECT 267.965 73.205 277.945 73.345 ;
        RECT 267.965 73.145 268.285 73.205 ;
        RECT 277.625 73.145 277.945 73.205 ;
        RECT 278.545 73.345 278.865 73.405 ;
        RECT 290.505 73.345 290.825 73.405 ;
        RECT 302.925 73.345 303.245 73.405 ;
        RECT 278.545 73.205 290.825 73.345 ;
        RECT 278.545 73.145 278.865 73.205 ;
        RECT 290.505 73.145 290.825 73.205 ;
        RECT 298.415 73.205 303.245 73.345 ;
        RECT 279.120 73.005 279.410 73.050 ;
        RECT 282.360 73.005 283.010 73.050 ;
        RECT 283.605 73.005 283.925 73.065 ;
        RECT 279.120 72.865 283.925 73.005 ;
        RECT 279.120 72.820 279.710 72.865 ;
        RECT 282.360 72.820 283.010 72.865 ;
        RECT 263.380 72.525 264.055 72.665 ;
        RECT 264.300 72.665 264.590 72.710 ;
        RECT 264.745 72.665 265.065 72.725 ;
        RECT 264.300 72.525 265.065 72.665 ;
        RECT 263.380 72.480 263.670 72.525 ;
        RECT 264.300 72.480 264.590 72.525 ;
        RECT 262.995 72.325 263.135 72.480 ;
        RECT 264.745 72.465 265.065 72.525 ;
        RECT 275.340 72.665 275.630 72.710 ;
        RECT 276.245 72.665 276.565 72.725 ;
        RECT 275.340 72.525 276.565 72.665 ;
        RECT 275.340 72.480 275.630 72.525 ;
        RECT 276.245 72.465 276.565 72.525 ;
        RECT 277.165 72.465 277.485 72.725 ;
        RECT 279.420 72.505 279.710 72.820 ;
        RECT 283.605 72.805 283.925 72.865 ;
        RECT 284.525 73.005 284.845 73.065 ;
        RECT 290.045 73.005 290.365 73.065 ;
        RECT 291.885 73.005 292.205 73.065 ;
        RECT 298.415 73.050 298.555 73.205 ;
        RECT 302.925 73.145 303.245 73.205 ;
        RECT 305.700 73.345 305.990 73.390 ;
        RECT 306.605 73.345 306.925 73.405 ;
        RECT 305.700 73.205 306.925 73.345 ;
        RECT 305.700 73.160 305.990 73.205 ;
        RECT 306.605 73.145 306.925 73.205 ;
        RECT 301.085 73.050 301.405 73.065 ;
        RECT 284.525 72.865 289.815 73.005 ;
        RECT 284.525 72.805 284.845 72.865 ;
        RECT 280.500 72.665 280.790 72.710 ;
        RECT 284.080 72.665 284.370 72.710 ;
        RECT 285.915 72.665 286.205 72.710 ;
        RECT 280.500 72.525 286.205 72.665 ;
        RECT 280.500 72.480 280.790 72.525 ;
        RECT 284.080 72.480 284.370 72.525 ;
        RECT 285.915 72.480 286.205 72.525 ;
        RECT 286.365 72.465 286.685 72.725 ;
        RECT 288.665 72.465 288.985 72.725 ;
        RECT 263.825 72.325 264.145 72.385 ;
        RECT 272.105 72.325 272.425 72.385 ;
        RECT 275.800 72.325 276.090 72.370 ;
        RECT 259.775 72.185 262.700 72.325 ;
        RECT 262.995 72.185 272.425 72.325 ;
        RECT 260.145 71.985 260.465 72.045 ;
        RECT 261.540 71.985 261.830 72.030 ;
        RECT 260.145 71.845 261.830 71.985 ;
        RECT 262.560 71.985 262.700 72.185 ;
        RECT 263.825 72.125 264.145 72.185 ;
        RECT 272.105 72.125 272.425 72.185 ;
        RECT 275.415 72.185 276.090 72.325 ;
        RECT 275.415 72.045 275.555 72.185 ;
        RECT 275.800 72.140 276.090 72.185 ;
        RECT 276.705 72.325 277.025 72.385 ;
        RECT 283.145 72.325 283.465 72.385 ;
        RECT 284.525 72.325 284.845 72.385 ;
        RECT 289.675 72.370 289.815 72.865 ;
        RECT 290.045 72.865 292.205 73.005 ;
        RECT 290.045 72.805 290.365 72.865 ;
        RECT 291.885 72.805 292.205 72.865 ;
        RECT 298.340 72.820 298.630 73.050 ;
        RECT 300.620 73.005 301.405 73.050 ;
        RECT 304.220 73.005 304.510 73.050 ;
        RECT 300.620 72.865 304.510 73.005 ;
        RECT 300.620 72.820 301.405 72.865 ;
        RECT 301.085 72.805 301.405 72.820 ;
        RECT 303.920 72.820 304.510 72.865 ;
        RECT 297.425 72.665 297.715 72.710 ;
        RECT 299.260 72.665 299.550 72.710 ;
        RECT 302.840 72.665 303.130 72.710 ;
        RECT 297.425 72.525 303.130 72.665 ;
        RECT 297.425 72.480 297.715 72.525 ;
        RECT 299.260 72.480 299.550 72.525 ;
        RECT 302.840 72.480 303.130 72.525 ;
        RECT 303.920 72.505 304.210 72.820 ;
        RECT 306.605 72.665 306.925 72.725 ;
        RECT 307.080 72.665 307.370 72.710 ;
        RECT 306.605 72.525 307.370 72.665 ;
        RECT 306.605 72.465 306.925 72.525 ;
        RECT 307.080 72.480 307.370 72.525 ;
        RECT 276.705 72.185 284.845 72.325 ;
        RECT 276.705 72.125 277.025 72.185 ;
        RECT 283.145 72.125 283.465 72.185 ;
        RECT 284.525 72.125 284.845 72.185 ;
        RECT 285.000 72.325 285.290 72.370 ;
        RECT 289.140 72.325 289.430 72.370 ;
        RECT 285.000 72.185 287.055 72.325 ;
        RECT 285.000 72.140 285.290 72.185 ;
        RECT 269.345 71.985 269.665 72.045 ;
        RECT 262.560 71.845 269.665 71.985 ;
        RECT 260.145 71.785 260.465 71.845 ;
        RECT 261.540 71.800 261.830 71.845 ;
        RECT 269.345 71.785 269.665 71.845 ;
        RECT 275.325 71.785 275.645 72.045 ;
        RECT 286.915 72.030 287.055 72.185 ;
        RECT 287.375 72.185 289.430 72.325 ;
        RECT 280.500 71.985 280.790 72.030 ;
        RECT 283.620 71.985 283.910 72.030 ;
        RECT 285.510 71.985 285.800 72.030 ;
        RECT 280.500 71.845 285.800 71.985 ;
        RECT 280.500 71.800 280.790 71.845 ;
        RECT 283.620 71.800 283.910 71.845 ;
        RECT 285.510 71.800 285.800 71.845 ;
        RECT 286.840 71.800 287.130 72.030 ;
        RECT 237.145 71.505 258.995 71.645 ;
        RECT 259.685 71.645 260.005 71.705 ;
        RECT 261.080 71.645 261.370 71.690 ;
        RECT 259.685 71.505 261.370 71.645 ;
        RECT 206.325 71.445 206.645 71.505 ;
        RECT 237.145 71.445 237.465 71.505 ;
        RECT 247.265 71.445 247.585 71.505 ;
        RECT 259.685 71.445 260.005 71.505 ;
        RECT 261.080 71.460 261.370 71.505 ;
        RECT 262.445 71.645 262.765 71.705 ;
        RECT 270.265 71.645 270.585 71.705 ;
        RECT 262.445 71.505 270.585 71.645 ;
        RECT 262.445 71.445 262.765 71.505 ;
        RECT 270.265 71.445 270.585 71.505 ;
        RECT 277.625 71.645 277.945 71.705 ;
        RECT 287.375 71.645 287.515 72.185 ;
        RECT 289.140 72.140 289.430 72.185 ;
        RECT 289.600 72.140 289.890 72.370 ;
        RECT 290.505 72.325 290.825 72.385 ;
        RECT 296.945 72.325 297.265 72.385 ;
        RECT 290.505 72.185 297.265 72.325 ;
        RECT 290.505 72.125 290.825 72.185 ;
        RECT 296.945 72.125 297.265 72.185 ;
        RECT 297.830 71.985 298.120 72.030 ;
        RECT 299.720 71.985 300.010 72.030 ;
        RECT 302.840 71.985 303.130 72.030 ;
        RECT 297.830 71.845 303.130 71.985 ;
        RECT 297.830 71.800 298.120 71.845 ;
        RECT 299.720 71.800 300.010 71.845 ;
        RECT 302.840 71.800 303.130 71.845 ;
        RECT 303.385 71.985 303.705 72.045 ;
        RECT 308.000 71.985 308.290 72.030 ;
        RECT 303.385 71.845 308.290 71.985 ;
        RECT 303.385 71.785 303.705 71.845 ;
        RECT 308.000 71.800 308.290 71.845 ;
        RECT 277.625 71.505 287.515 71.645 ;
        RECT 290.045 71.645 290.365 71.705 ;
        RECT 300.165 71.645 300.485 71.705 ;
        RECT 290.045 71.505 300.485 71.645 ;
        RECT 277.625 71.445 277.945 71.505 ;
        RECT 290.045 71.445 290.365 71.505 ;
        RECT 300.165 71.445 300.485 71.505 ;
        RECT 301.085 71.645 301.405 71.705 ;
        RECT 303.845 71.645 304.165 71.705 ;
        RECT 301.085 71.505 304.165 71.645 ;
        RECT 301.085 71.445 301.405 71.505 ;
        RECT 303.845 71.445 304.165 71.505 ;
        RECT 162.095 70.825 311.135 71.305 ;
        RECT 173.205 70.625 173.525 70.685 ;
        RECT 190.685 70.625 191.005 70.685 ;
        RECT 173.205 70.485 186.315 70.625 ;
        RECT 173.205 70.425 173.525 70.485 ;
        RECT 170.920 70.285 171.210 70.330 ;
        RECT 174.125 70.285 174.445 70.345 ;
        RECT 170.920 70.145 174.445 70.285 ;
        RECT 170.920 70.100 171.210 70.145 ;
        RECT 174.125 70.085 174.445 70.145 ;
        RECT 174.585 70.285 174.905 70.345 ;
        RECT 177.345 70.285 177.665 70.345 ;
        RECT 174.585 70.145 177.665 70.285 ;
        RECT 174.585 70.085 174.905 70.145 ;
        RECT 177.345 70.085 177.665 70.145 ;
        RECT 173.680 69.945 173.970 69.990 ;
        RECT 178.740 69.945 179.030 69.990 ;
        RECT 179.645 69.945 179.965 70.005 ;
        RECT 173.680 69.805 179.965 69.945 ;
        RECT 173.680 69.760 173.970 69.805 ;
        RECT 178.740 69.760 179.030 69.805 ;
        RECT 179.645 69.745 179.965 69.805 ;
        RECT 172.760 69.605 173.050 69.650 ;
        RECT 175.965 69.605 176.285 69.665 ;
        RECT 172.760 69.465 176.285 69.605 ;
        RECT 172.760 69.420 173.050 69.465 ;
        RECT 175.965 69.405 176.285 69.465 ;
        RECT 183.340 69.605 183.630 69.650 ;
        RECT 185.625 69.605 185.945 69.665 ;
        RECT 186.175 69.650 186.315 70.485 ;
        RECT 190.685 70.485 194.595 70.625 ;
        RECT 190.685 70.425 191.005 70.485 ;
        RECT 187.555 70.145 194.135 70.285 ;
        RECT 183.340 69.465 185.945 69.605 ;
        RECT 183.340 69.420 183.630 69.465 ;
        RECT 185.625 69.405 185.945 69.465 ;
        RECT 186.100 69.605 186.390 69.650 ;
        RECT 187.005 69.605 187.325 69.665 ;
        RECT 187.555 69.650 187.695 70.145 ;
        RECT 188.385 69.945 188.705 70.005 ;
        RECT 188.860 69.945 189.150 69.990 ;
        RECT 192.525 69.945 192.845 70.005 ;
        RECT 188.385 69.805 192.845 69.945 ;
        RECT 188.385 69.745 188.705 69.805 ;
        RECT 188.860 69.760 189.150 69.805 ;
        RECT 192.525 69.745 192.845 69.805 ;
        RECT 193.995 69.665 194.135 70.145 ;
        RECT 194.455 70.005 194.595 70.485 ;
        RECT 201.265 70.425 201.585 70.685 ;
        RECT 205.865 70.625 206.185 70.685 ;
        RECT 219.665 70.625 219.985 70.685 ;
        RECT 230.245 70.625 230.565 70.685 ;
        RECT 205.865 70.485 214.835 70.625 ;
        RECT 205.865 70.425 206.185 70.485 ;
        RECT 205.955 70.285 206.095 70.425 ;
        RECT 203.655 70.145 206.095 70.285 ;
        RECT 194.365 69.945 194.685 70.005 ;
        RECT 203.655 69.990 203.795 70.145 ;
        RECT 213.685 70.085 214.005 70.345 ;
        RECT 194.365 69.805 198.275 69.945 ;
        RECT 194.365 69.745 194.685 69.805 ;
        RECT 186.100 69.465 187.325 69.605 ;
        RECT 186.100 69.420 186.390 69.465 ;
        RECT 187.005 69.405 187.325 69.465 ;
        RECT 187.480 69.420 187.770 69.650 ;
        RECT 189.855 69.465 193.675 69.605 ;
        RECT 164.465 69.265 164.785 69.325 ;
        RECT 177.820 69.265 178.110 69.310 ;
        RECT 189.855 69.265 189.995 69.465 ;
        RECT 164.465 69.125 189.995 69.265 ;
        RECT 190.225 69.265 190.545 69.325 ;
        RECT 192.540 69.265 192.830 69.310 ;
        RECT 190.225 69.125 192.830 69.265 ;
        RECT 193.535 69.265 193.675 69.465 ;
        RECT 193.905 69.405 194.225 69.665 ;
        RECT 196.205 69.405 196.525 69.665 ;
        RECT 197.125 69.605 197.445 69.665 ;
        RECT 197.600 69.605 197.890 69.650 ;
        RECT 197.125 69.465 197.890 69.605 ;
        RECT 198.135 69.605 198.275 69.805 ;
        RECT 203.580 69.760 203.870 69.990 ;
        RECT 204.500 69.945 204.790 69.990 ;
        RECT 206.785 69.945 207.105 70.005 ;
        RECT 204.500 69.805 207.105 69.945 ;
        RECT 204.500 69.760 204.790 69.805 ;
        RECT 206.785 69.745 207.105 69.805 ;
        RECT 208.165 69.945 208.485 70.005 ;
        RECT 213.775 69.945 213.915 70.085 ;
        RECT 208.165 69.805 213.915 69.945 ;
        RECT 208.165 69.745 208.485 69.805 ;
        RECT 211.385 69.605 211.705 69.665 ;
        RECT 198.135 69.465 211.705 69.605 ;
        RECT 197.125 69.405 197.445 69.465 ;
        RECT 197.600 69.420 197.890 69.465 ;
        RECT 211.385 69.405 211.705 69.465 ;
        RECT 211.860 69.420 212.150 69.650 ;
        RECT 212.305 69.605 212.625 69.665 ;
        RECT 213.315 69.650 213.455 69.805 ;
        RECT 212.780 69.605 213.070 69.650 ;
        RECT 212.305 69.465 213.070 69.605 ;
        RECT 210.465 69.265 210.785 69.325 ;
        RECT 211.935 69.265 212.075 69.420 ;
        RECT 212.305 69.405 212.625 69.465 ;
        RECT 212.780 69.420 213.070 69.465 ;
        RECT 213.240 69.420 213.530 69.650 ;
        RECT 213.685 69.405 214.005 69.665 ;
        RECT 214.695 69.605 214.835 70.485 ;
        RECT 219.665 70.485 230.565 70.625 ;
        RECT 219.665 70.425 219.985 70.485 ;
        RECT 230.245 70.425 230.565 70.485 ;
        RECT 233.465 70.425 233.785 70.685 ;
        RECT 241.285 70.625 241.605 70.685 ;
        RECT 256.925 70.625 257.245 70.685 ;
        RECT 261.525 70.625 261.845 70.685 ;
        RECT 241.285 70.485 257.245 70.625 ;
        RECT 241.285 70.425 241.605 70.485 ;
        RECT 217.365 70.285 217.685 70.345 ;
        RECT 228.865 70.285 229.185 70.345 ;
        RECT 231.625 70.285 231.945 70.345 ;
        RECT 217.365 70.145 220.815 70.285 ;
        RECT 217.365 70.085 217.685 70.145 ;
        RECT 215.080 69.945 215.370 69.990 ;
        RECT 220.125 69.945 220.445 70.005 ;
        RECT 215.080 69.805 220.445 69.945 ;
        RECT 220.675 69.945 220.815 70.145 ;
        RECT 228.865 70.145 231.945 70.285 ;
        RECT 228.865 70.085 229.185 70.145 ;
        RECT 231.625 70.085 231.945 70.145 ;
        RECT 235.305 70.285 235.625 70.345 ;
        RECT 244.980 70.285 245.270 70.330 ;
        RECT 245.425 70.285 245.745 70.345 ;
        RECT 235.305 70.145 245.745 70.285 ;
        RECT 235.305 70.085 235.625 70.145 ;
        RECT 244.980 70.100 245.270 70.145 ;
        RECT 245.425 70.085 245.745 70.145 ;
        RECT 220.675 69.805 247.035 69.945 ;
        RECT 215.080 69.760 215.370 69.805 ;
        RECT 220.125 69.745 220.445 69.805 ;
        RECT 241.745 69.605 242.065 69.665 ;
        RECT 214.695 69.465 245.655 69.605 ;
        RECT 241.745 69.405 242.065 69.465 ;
        RECT 229.325 69.265 229.645 69.325 ;
        RECT 193.535 69.125 211.615 69.265 ;
        RECT 211.935 69.125 229.645 69.265 ;
        RECT 164.465 69.065 164.785 69.125 ;
        RECT 177.820 69.080 178.110 69.125 ;
        RECT 190.225 69.065 190.545 69.125 ;
        RECT 192.540 69.080 192.830 69.125 ;
        RECT 210.465 69.065 210.785 69.125 ;
        RECT 172.285 68.925 172.605 68.985 ;
        RECT 173.220 68.925 173.510 68.970 ;
        RECT 172.285 68.785 173.510 68.925 ;
        RECT 172.285 68.725 172.605 68.785 ;
        RECT 173.220 68.740 173.510 68.785 ;
        RECT 175.505 68.725 175.825 68.985 ;
        RECT 177.345 68.925 177.665 68.985 ;
        RECT 182.865 68.925 183.185 68.985 ;
        RECT 177.345 68.785 183.185 68.925 ;
        RECT 177.345 68.725 177.665 68.785 ;
        RECT 182.865 68.725 183.185 68.785 ;
        RECT 183.785 68.925 184.105 68.985 ;
        RECT 186.085 68.925 186.405 68.985 ;
        RECT 183.785 68.785 186.405 68.925 ;
        RECT 183.785 68.725 184.105 68.785 ;
        RECT 186.085 68.725 186.405 68.785 ;
        RECT 187.020 68.925 187.310 68.970 ;
        RECT 192.065 68.925 192.385 68.985 ;
        RECT 187.020 68.785 192.385 68.925 ;
        RECT 187.020 68.740 187.310 68.785 ;
        RECT 192.065 68.725 192.385 68.785 ;
        RECT 197.600 68.925 197.890 68.970 ;
        RECT 202.185 68.925 202.505 68.985 ;
        RECT 197.600 68.785 202.505 68.925 ;
        RECT 197.600 68.740 197.890 68.785 ;
        RECT 202.185 68.725 202.505 68.785 ;
        RECT 203.105 68.725 203.425 68.985 ;
        RECT 211.475 68.925 211.615 69.125 ;
        RECT 229.325 69.065 229.645 69.125 ;
        RECT 234.385 69.065 234.705 69.325 ;
        RECT 235.305 69.065 235.625 69.325 ;
        RECT 236.240 69.265 236.530 69.310 ;
        RECT 236.240 69.125 242.435 69.265 ;
        RECT 236.240 69.080 236.530 69.125 ;
        RECT 213.685 68.925 214.005 68.985 ;
        RECT 211.475 68.785 214.005 68.925 ;
        RECT 213.685 68.725 214.005 68.785 ;
        RECT 218.745 68.925 219.065 68.985 ;
        RECT 233.005 68.925 233.325 68.985 ;
        RECT 218.745 68.785 233.325 68.925 ;
        RECT 218.745 68.725 219.065 68.785 ;
        RECT 233.005 68.725 233.325 68.785 ;
        RECT 234.860 68.925 235.150 68.970 ;
        RECT 240.825 68.925 241.145 68.985 ;
        RECT 234.860 68.785 241.145 68.925 ;
        RECT 234.860 68.740 235.150 68.785 ;
        RECT 240.825 68.725 241.145 68.785 ;
        RECT 241.285 68.725 241.605 68.985 ;
        RECT 242.295 68.970 242.435 69.125 ;
        RECT 242.665 69.065 242.985 69.325 ;
        RECT 244.505 69.265 244.825 69.325 ;
        RECT 243.675 69.125 244.825 69.265 ;
        RECT 242.220 68.925 242.510 68.970 ;
        RECT 243.675 68.925 243.815 69.125 ;
        RECT 244.505 69.065 244.825 69.125 ;
        RECT 244.965 69.065 245.285 69.325 ;
        RECT 245.515 69.265 245.655 69.465 ;
        RECT 245.885 69.405 246.205 69.665 ;
        RECT 246.365 69.420 246.655 69.650 ;
        RECT 246.440 69.265 246.580 69.420 ;
        RECT 245.515 69.125 246.580 69.265 ;
        RECT 246.895 69.265 247.035 69.805 ;
        RECT 247.265 69.405 247.585 69.665 ;
        RECT 247.725 69.405 248.045 69.665 ;
        RECT 248.275 69.650 248.415 70.485 ;
        RECT 256.925 70.425 257.245 70.485 ;
        RECT 260.465 70.485 261.845 70.625 ;
        RECT 258.765 70.285 259.085 70.345 ;
        RECT 260.465 70.285 260.605 70.485 ;
        RECT 261.525 70.425 261.845 70.485 ;
        RECT 264.760 70.625 265.050 70.670 ;
        RECT 265.220 70.625 265.510 70.670 ;
        RECT 264.760 70.485 265.510 70.625 ;
        RECT 264.760 70.440 265.050 70.485 ;
        RECT 265.220 70.440 265.510 70.485 ;
        RECT 277.640 70.625 277.930 70.670 ;
        RECT 290.965 70.625 291.285 70.685 ;
        RECT 294.645 70.625 294.965 70.685 ;
        RECT 277.640 70.485 294.965 70.625 ;
        RECT 277.640 70.440 277.930 70.485 ;
        RECT 290.965 70.425 291.285 70.485 ;
        RECT 294.645 70.425 294.965 70.485 ;
        RECT 304.305 70.425 304.625 70.685 ;
        RECT 258.765 70.145 260.605 70.285 ;
        RECT 261.080 70.285 261.370 70.330 ;
        RECT 265.665 70.285 265.985 70.345 ;
        RECT 278.085 70.285 278.405 70.345 ;
        RECT 261.080 70.145 265.985 70.285 ;
        RECT 258.765 70.085 259.085 70.145 ;
        RECT 256.465 69.945 256.785 70.005 ;
        RECT 256.465 69.805 258.540 69.945 ;
        RECT 256.465 69.745 256.785 69.805 ;
        RECT 248.225 69.420 248.515 69.650 ;
        RECT 256.925 69.605 257.245 69.665 ;
        RECT 258.400 69.650 258.540 69.805 ;
        RECT 259.225 69.745 259.545 70.005 ;
        RECT 257.860 69.605 258.150 69.650 ;
        RECT 256.925 69.465 258.150 69.605 ;
        RECT 256.925 69.405 257.245 69.465 ;
        RECT 257.860 69.420 258.150 69.465 ;
        RECT 258.325 69.420 258.615 69.650 ;
        RECT 259.315 69.605 259.455 69.745 ;
        RECT 260.260 69.650 260.400 70.145 ;
        RECT 261.080 70.100 261.370 70.145 ;
        RECT 265.665 70.085 265.985 70.145 ;
        RECT 266.215 70.145 278.405 70.285 ;
        RECT 260.605 69.945 260.925 70.005 ;
        RECT 266.215 69.945 266.355 70.145 ;
        RECT 278.085 70.085 278.405 70.145 ;
        RECT 279.430 70.285 279.720 70.330 ;
        RECT 281.320 70.285 281.610 70.330 ;
        RECT 284.440 70.285 284.730 70.330 ;
        RECT 279.430 70.145 284.730 70.285 ;
        RECT 279.430 70.100 279.720 70.145 ;
        RECT 281.320 70.100 281.610 70.145 ;
        RECT 284.440 70.100 284.730 70.145 ;
        RECT 285.445 70.285 285.765 70.345 ;
        RECT 288.665 70.285 288.985 70.345 ;
        RECT 292.310 70.285 292.600 70.330 ;
        RECT 294.200 70.285 294.490 70.330 ;
        RECT 297.320 70.285 297.610 70.330 ;
        RECT 305.225 70.285 305.545 70.345 ;
        RECT 285.445 70.145 292.115 70.285 ;
        RECT 285.445 70.085 285.765 70.145 ;
        RECT 288.665 70.085 288.985 70.145 ;
        RECT 260.605 69.805 266.355 69.945 ;
        RECT 266.585 69.945 266.905 70.005 ;
        RECT 272.580 69.945 272.870 69.990 ;
        RECT 275.800 69.945 276.090 69.990 ;
        RECT 266.585 69.805 276.090 69.945 ;
        RECT 260.605 69.745 260.925 69.805 ;
        RECT 259.700 69.605 259.990 69.650 ;
        RECT 258.855 69.465 259.990 69.605 ;
        RECT 256.465 69.265 256.785 69.325 ;
        RECT 258.855 69.265 258.995 69.465 ;
        RECT 259.700 69.420 259.990 69.465 ;
        RECT 260.185 69.420 260.475 69.650 ;
        RECT 261.065 69.605 261.385 69.665 ;
        RECT 262.445 69.650 262.765 69.665 ;
        RECT 262.995 69.650 263.135 69.805 ;
        RECT 266.585 69.745 266.905 69.805 ;
        RECT 272.580 69.760 272.870 69.805 ;
        RECT 275.800 69.760 276.090 69.805 ;
        RECT 278.545 69.745 278.865 70.005 ;
        RECT 290.505 69.945 290.825 70.005 ;
        RECT 291.440 69.945 291.730 69.990 ;
        RECT 290.505 69.805 291.730 69.945 ;
        RECT 291.975 69.945 292.115 70.145 ;
        RECT 292.310 70.145 297.610 70.285 ;
        RECT 292.310 70.100 292.600 70.145 ;
        RECT 294.200 70.100 294.490 70.145 ;
        RECT 297.320 70.100 297.610 70.145 ;
        RECT 303.475 70.145 305.545 70.285 ;
        RECT 303.475 69.945 303.615 70.145 ;
        RECT 305.225 70.085 305.545 70.145 ;
        RECT 291.975 69.805 303.615 69.945 ;
        RECT 303.845 69.945 304.165 70.005 ;
        RECT 307.080 69.945 307.370 69.990 ;
        RECT 303.845 69.805 307.370 69.945 ;
        RECT 290.505 69.745 290.825 69.805 ;
        RECT 291.440 69.760 291.730 69.805 ;
        RECT 303.845 69.745 304.165 69.805 ;
        RECT 307.080 69.760 307.370 69.805 ;
        RECT 264.285 69.650 264.605 69.665 ;
        RECT 261.540 69.605 261.830 69.650 ;
        RECT 261.065 69.465 261.830 69.605 ;
        RECT 261.065 69.405 261.385 69.465 ;
        RECT 261.540 69.420 261.830 69.465 ;
        RECT 262.280 69.420 262.765 69.650 ;
        RECT 262.920 69.420 263.210 69.650 ;
        RECT 264.070 69.420 264.605 69.650 ;
        RECT 262.445 69.405 262.765 69.420 ;
        RECT 264.285 69.405 264.605 69.420 ;
        RECT 265.205 69.405 265.525 69.665 ;
        RECT 265.665 69.405 265.985 69.665 ;
        RECT 269.805 69.605 270.125 69.665 ;
        RECT 270.280 69.605 270.570 69.650 ;
        RECT 269.805 69.465 270.570 69.605 ;
        RECT 269.805 69.405 270.125 69.465 ;
        RECT 270.280 69.420 270.570 69.465 ;
        RECT 270.725 69.405 271.045 69.665 ;
        RECT 275.325 69.405 275.645 69.665 ;
        RECT 276.720 69.605 277.010 69.650 ;
        RECT 277.165 69.605 277.485 69.665 ;
        RECT 276.720 69.465 277.485 69.605 ;
        RECT 276.720 69.420 277.010 69.465 ;
        RECT 277.165 69.405 277.485 69.465 ;
        RECT 279.025 69.605 279.315 69.650 ;
        RECT 280.860 69.605 281.150 69.650 ;
        RECT 284.440 69.605 284.730 69.650 ;
        RECT 279.025 69.465 284.730 69.605 ;
        RECT 279.025 69.420 279.315 69.465 ;
        RECT 280.860 69.420 281.150 69.465 ;
        RECT 284.440 69.420 284.730 69.465 ;
        RECT 246.895 69.125 256.005 69.265 ;
        RECT 242.220 68.785 243.815 68.925 ;
        RECT 242.220 68.740 242.510 68.785 ;
        RECT 249.105 68.725 249.425 68.985 ;
        RECT 255.865 68.925 256.005 69.125 ;
        RECT 256.465 69.125 258.995 69.265 ;
        RECT 256.465 69.065 256.785 69.125 ;
        RECT 259.225 69.065 259.545 69.325 ;
        RECT 263.380 69.265 263.670 69.310 ;
        RECT 267.965 69.265 268.285 69.325 ;
        RECT 263.380 69.125 268.285 69.265 ;
        RECT 263.380 69.080 263.670 69.125 ;
        RECT 267.965 69.065 268.285 69.125 ;
        RECT 273.025 69.065 273.345 69.325 ;
        RECT 279.465 69.265 279.785 69.325 ;
        RECT 279.940 69.265 280.230 69.310 ;
        RECT 279.465 69.125 280.230 69.265 ;
        RECT 279.465 69.065 279.785 69.125 ;
        RECT 279.940 69.080 280.230 69.125 ;
        RECT 282.220 69.265 282.870 69.310 ;
        RECT 283.605 69.265 283.925 69.325 ;
        RECT 285.520 69.310 285.810 69.625 ;
        RECT 291.905 69.605 292.195 69.650 ;
        RECT 293.740 69.605 294.030 69.650 ;
        RECT 297.320 69.605 297.610 69.650 ;
        RECT 291.905 69.465 297.610 69.605 ;
        RECT 291.905 69.420 292.195 69.465 ;
        RECT 293.740 69.420 294.030 69.465 ;
        RECT 297.320 69.420 297.610 69.465 ;
        RECT 285.520 69.265 286.110 69.310 ;
        RECT 282.220 69.125 286.110 69.265 ;
        RECT 282.220 69.080 282.870 69.125 ;
        RECT 283.605 69.065 283.925 69.125 ;
        RECT 285.820 69.080 286.110 69.125 ;
        RECT 291.425 69.265 291.745 69.325 ;
        RECT 298.400 69.310 298.690 69.625 ;
        RECT 300.165 69.605 300.485 69.665 ;
        RECT 302.940 69.605 303.230 69.650 ;
        RECT 303.385 69.605 303.705 69.665 ;
        RECT 300.165 69.465 301.775 69.605 ;
        RECT 300.165 69.405 300.485 69.465 ;
        RECT 292.820 69.265 293.110 69.310 ;
        RECT 291.425 69.125 293.110 69.265 ;
        RECT 291.425 69.065 291.745 69.125 ;
        RECT 292.820 69.080 293.110 69.125 ;
        RECT 295.100 69.265 295.750 69.310 ;
        RECT 298.400 69.265 298.990 69.310 ;
        RECT 301.085 69.265 301.405 69.325 ;
        RECT 295.100 69.125 301.405 69.265 ;
        RECT 301.635 69.265 301.775 69.465 ;
        RECT 302.940 69.465 303.705 69.605 ;
        RECT 302.940 69.420 303.230 69.465 ;
        RECT 303.385 69.405 303.705 69.465 ;
        RECT 304.765 69.605 305.085 69.665 ;
        RECT 306.160 69.605 306.450 69.650 ;
        RECT 304.765 69.465 306.450 69.605 ;
        RECT 304.765 69.405 305.085 69.465 ;
        RECT 306.160 69.420 306.450 69.465 ;
        RECT 306.620 69.265 306.910 69.310 ;
        RECT 301.635 69.125 306.910 69.265 ;
        RECT 295.100 69.080 295.750 69.125 ;
        RECT 298.700 69.080 298.990 69.125 ;
        RECT 301.085 69.065 301.405 69.125 ;
        RECT 306.620 69.080 306.910 69.125 ;
        RECT 267.060 68.925 267.350 68.970 ;
        RECT 255.865 68.785 267.350 68.925 ;
        RECT 267.060 68.740 267.350 68.785 ;
        RECT 281.765 68.925 282.085 68.985 ;
        RECT 287.300 68.925 287.590 68.970 ;
        RECT 281.765 68.785 287.590 68.925 ;
        RECT 281.765 68.725 282.085 68.785 ;
        RECT 287.300 68.740 287.590 68.785 ;
        RECT 293.265 68.925 293.585 68.985 ;
        RECT 300.180 68.925 300.470 68.970 ;
        RECT 293.265 68.785 300.470 68.925 ;
        RECT 293.265 68.725 293.585 68.785 ;
        RECT 300.180 68.740 300.470 68.785 ;
        RECT 162.095 68.105 311.135 68.585 ;
        RECT 166.780 67.905 167.070 67.950 ;
        RECT 167.225 67.905 167.545 67.965 ;
        RECT 172.285 67.905 172.605 67.965 ;
        RECT 166.780 67.765 172.605 67.905 ;
        RECT 166.780 67.720 167.070 67.765 ;
        RECT 167.225 67.705 167.545 67.765 ;
        RECT 172.285 67.705 172.605 67.765 ;
        RECT 195.285 67.905 195.605 67.965 ;
        RECT 199.425 67.905 199.745 67.965 ;
        RECT 210.020 67.905 210.310 67.950 ;
        RECT 212.765 67.905 213.085 67.965 ;
        RECT 195.285 67.765 207.705 67.905 ;
        RECT 195.285 67.705 195.605 67.765 ;
        RECT 199.425 67.705 199.745 67.765 ;
        RECT 168.260 67.565 168.550 67.610 ;
        RECT 171.500 67.565 172.150 67.610 ;
        RECT 172.745 67.565 173.065 67.625 ;
        RECT 168.260 67.425 173.065 67.565 ;
        RECT 168.260 67.380 168.850 67.425 ;
        RECT 171.500 67.380 172.150 67.425 ;
        RECT 168.560 67.065 168.850 67.380 ;
        RECT 172.745 67.365 173.065 67.425 ;
        RECT 174.125 67.365 174.445 67.625 ;
        RECT 181.025 67.610 181.345 67.625 ;
        RECT 180.560 67.565 181.345 67.610 ;
        RECT 184.160 67.565 184.450 67.610 ;
        RECT 180.560 67.425 184.450 67.565 ;
        RECT 180.560 67.380 181.345 67.425 ;
        RECT 181.025 67.365 181.345 67.380 ;
        RECT 183.860 67.380 184.450 67.425 ;
        RECT 185.165 67.565 185.485 67.625 ;
        RECT 189.305 67.565 189.625 67.625 ;
        RECT 191.620 67.565 191.910 67.610 ;
        RECT 185.165 67.425 189.075 67.565 ;
        RECT 169.640 67.225 169.930 67.270 ;
        RECT 173.220 67.225 173.510 67.270 ;
        RECT 175.055 67.225 175.345 67.270 ;
        RECT 169.640 67.085 175.345 67.225 ;
        RECT 169.640 67.040 169.930 67.085 ;
        RECT 173.220 67.040 173.510 67.085 ;
        RECT 175.055 67.040 175.345 67.085 ;
        RECT 175.520 67.225 175.810 67.270 ;
        RECT 176.885 67.225 177.205 67.285 ;
        RECT 175.520 67.085 177.205 67.225 ;
        RECT 175.520 67.040 175.810 67.085 ;
        RECT 176.885 67.025 177.205 67.085 ;
        RECT 177.365 67.225 177.655 67.270 ;
        RECT 179.200 67.225 179.490 67.270 ;
        RECT 182.780 67.225 183.070 67.270 ;
        RECT 177.365 67.085 183.070 67.225 ;
        RECT 177.365 67.040 177.655 67.085 ;
        RECT 179.200 67.040 179.490 67.085 ;
        RECT 182.780 67.040 183.070 67.085 ;
        RECT 183.860 67.065 184.150 67.380 ;
        RECT 185.165 67.365 185.485 67.425 ;
        RECT 188.400 67.040 188.690 67.270 ;
        RECT 188.935 67.225 189.075 67.425 ;
        RECT 189.305 67.425 191.910 67.565 ;
        RECT 189.305 67.365 189.625 67.425 ;
        RECT 191.620 67.380 191.910 67.425 ;
        RECT 192.525 67.365 192.845 67.625 ;
        RECT 196.665 67.565 196.985 67.625 ;
        RECT 207.565 67.565 207.705 67.765 ;
        RECT 210.020 67.765 213.085 67.905 ;
        RECT 210.020 67.720 210.310 67.765 ;
        RECT 212.765 67.705 213.085 67.765 ;
        RECT 213.240 67.905 213.530 67.950 ;
        RECT 215.065 67.905 215.385 67.965 ;
        RECT 213.240 67.765 215.385 67.905 ;
        RECT 213.240 67.720 213.530 67.765 ;
        RECT 215.065 67.705 215.385 67.765 ;
        RECT 218.285 67.905 218.605 67.965 ;
        RECT 230.705 67.905 231.025 67.965 ;
        RECT 256.005 67.905 256.325 67.965 ;
        RECT 259.225 67.905 259.545 67.965 ;
        RECT 218.285 67.765 221.505 67.905 ;
        RECT 218.285 67.705 218.605 67.765 ;
        RECT 212.305 67.565 212.625 67.625 ;
        RECT 220.585 67.565 220.905 67.625 ;
        RECT 196.665 67.425 199.195 67.565 ;
        RECT 207.565 67.425 212.625 67.565 ;
        RECT 196.665 67.365 196.985 67.425 ;
        RECT 199.055 67.285 199.195 67.425 ;
        RECT 190.240 67.225 190.530 67.270 ;
        RECT 188.935 67.085 190.530 67.225 ;
        RECT 190.240 67.040 190.530 67.085 ;
        RECT 191.160 67.225 191.450 67.270 ;
        RECT 194.365 67.225 194.685 67.285 ;
        RECT 191.160 67.085 194.685 67.225 ;
        RECT 191.160 67.040 191.450 67.085 ;
        RECT 169.640 66.545 169.930 66.590 ;
        RECT 172.760 66.545 173.050 66.590 ;
        RECT 174.650 66.545 174.940 66.590 ;
        RECT 169.640 66.405 174.940 66.545 ;
        RECT 169.640 66.360 169.930 66.405 ;
        RECT 172.760 66.360 173.050 66.405 ;
        RECT 174.650 66.360 174.940 66.405 ;
        RECT 177.770 66.545 178.060 66.590 ;
        RECT 179.660 66.545 179.950 66.590 ;
        RECT 182.780 66.545 183.070 66.590 ;
        RECT 188.475 66.545 188.615 67.040 ;
        RECT 189.305 66.885 189.625 66.945 ;
        RECT 191.235 66.885 191.375 67.040 ;
        RECT 194.365 67.025 194.685 67.085 ;
        RECT 197.585 67.270 197.905 67.285 ;
        RECT 197.585 67.040 198.120 67.270 ;
        RECT 198.520 67.040 198.810 67.270 ;
        RECT 198.980 67.055 199.270 67.285 ;
        RECT 197.585 67.025 197.905 67.040 ;
        RECT 189.305 66.745 191.375 66.885 ;
        RECT 189.305 66.685 189.625 66.745 ;
        RECT 191.145 66.545 191.465 66.605 ;
        RECT 177.770 66.405 183.070 66.545 ;
        RECT 177.770 66.360 178.060 66.405 ;
        RECT 179.660 66.360 179.950 66.405 ;
        RECT 182.780 66.360 183.070 66.405 ;
        RECT 185.255 66.405 186.775 66.545 ;
        RECT 188.475 66.405 191.465 66.545 ;
        RECT 198.595 66.545 198.735 67.040 ;
        RECT 199.885 67.025 200.205 67.285 ;
        RECT 200.345 67.225 200.665 67.285 ;
        RECT 200.345 67.085 201.035 67.225 ;
        RECT 200.345 67.025 200.665 67.085 ;
        RECT 200.895 66.885 201.035 67.085 ;
        RECT 207.705 67.025 208.025 67.285 ;
        RECT 208.165 67.025 208.485 67.285 ;
        RECT 209.175 67.270 209.315 67.425 ;
        RECT 212.305 67.365 212.625 67.425 ;
        RECT 219.755 67.425 220.905 67.565 ;
        RECT 221.365 67.565 221.505 67.765 ;
        RECT 230.705 67.765 259.545 67.905 ;
        RECT 230.705 67.705 231.025 67.765 ;
        RECT 256.005 67.705 256.325 67.765 ;
        RECT 259.225 67.705 259.545 67.765 ;
        RECT 259.685 67.905 260.005 67.965 ;
        RECT 259.685 67.765 262.215 67.905 ;
        RECT 259.685 67.705 260.005 67.765 ;
        RECT 249.105 67.565 249.425 67.625 ;
        RECT 221.365 67.425 224.035 67.565 ;
        RECT 209.100 67.040 209.390 67.270 ;
        RECT 211.845 67.025 212.165 67.285 ;
        RECT 214.145 67.225 214.465 67.285 ;
        RECT 215.540 67.225 215.830 67.270 ;
        RECT 214.145 67.085 215.830 67.225 ;
        RECT 214.145 67.025 214.465 67.085 ;
        RECT 215.540 67.040 215.830 67.085 ;
        RECT 216.000 67.040 216.290 67.270 ;
        RECT 210.005 66.885 210.325 66.945 ;
        RECT 200.895 66.745 210.325 66.885 ;
        RECT 210.005 66.685 210.325 66.745 ;
        RECT 210.940 66.700 211.230 66.930 ;
        RECT 211.400 66.700 211.690 66.930 ;
        RECT 201.280 66.545 201.570 66.590 ;
        RECT 202.645 66.545 202.965 66.605 ;
        RECT 198.595 66.405 202.965 66.545 ;
        RECT 178.215 66.205 178.505 66.250 ;
        RECT 180.565 66.205 180.885 66.265 ;
        RECT 178.215 66.065 180.885 66.205 ;
        RECT 178.215 66.020 178.505 66.065 ;
        RECT 180.565 66.005 180.885 66.065 ;
        RECT 183.785 66.205 184.105 66.265 ;
        RECT 185.255 66.205 185.395 66.405 ;
        RECT 183.785 66.065 185.395 66.205 ;
        RECT 185.640 66.205 185.930 66.250 ;
        RECT 186.085 66.205 186.405 66.265 ;
        RECT 185.640 66.065 186.405 66.205 ;
        RECT 186.635 66.205 186.775 66.405 ;
        RECT 191.145 66.345 191.465 66.405 ;
        RECT 201.280 66.360 201.570 66.405 ;
        RECT 202.645 66.345 202.965 66.405 ;
        RECT 208.625 66.545 208.945 66.605 ;
        RECT 211.015 66.545 211.155 66.700 ;
        RECT 208.625 66.405 211.155 66.545 ;
        RECT 211.475 66.545 211.615 66.700 ;
        RECT 212.305 66.685 212.625 66.945 ;
        RECT 213.225 66.685 213.545 66.945 ;
        RECT 213.685 66.885 214.005 66.945 ;
        RECT 216.075 66.885 216.215 67.040 ;
        RECT 216.445 67.025 216.765 67.285 ;
        RECT 217.365 67.025 217.685 67.285 ;
        RECT 217.825 67.025 218.145 67.285 ;
        RECT 218.745 67.025 219.065 67.285 ;
        RECT 219.205 67.025 219.525 67.285 ;
        RECT 219.755 67.270 219.895 67.425 ;
        RECT 220.585 67.365 220.905 67.425 ;
        RECT 223.895 67.270 224.035 67.425 ;
        RECT 224.815 67.425 249.425 67.565 ;
        RECT 224.815 67.270 224.955 67.425 ;
        RECT 249.105 67.365 249.425 67.425 ;
        RECT 254.165 67.565 254.485 67.625 ;
        RECT 260.160 67.565 260.450 67.610 ;
        RECT 254.165 67.425 259.915 67.565 ;
        RECT 254.165 67.365 254.485 67.425 ;
        RECT 219.680 67.040 219.970 67.270 ;
        RECT 222.900 67.040 223.190 67.270 ;
        RECT 223.820 67.040 224.110 67.270 ;
        RECT 224.740 67.040 225.030 67.270 ;
        RECT 225.200 67.225 225.490 67.270 ;
        RECT 227.040 67.225 227.330 67.270 ;
        RECT 225.200 67.085 227.330 67.225 ;
        RECT 225.200 67.040 225.490 67.085 ;
        RECT 227.040 67.040 227.330 67.085 ;
        RECT 222.975 66.885 223.115 67.040 ;
        RECT 227.945 67.025 228.265 67.285 ;
        RECT 228.880 67.225 229.170 67.270 ;
        RECT 240.365 67.225 240.685 67.285 ;
        RECT 228.880 67.085 240.685 67.225 ;
        RECT 228.880 67.040 229.170 67.085 ;
        RECT 240.365 67.025 240.685 67.085 ;
        RECT 240.825 67.225 241.145 67.285 ;
        RECT 244.045 67.225 244.365 67.285 ;
        RECT 244.965 67.225 245.285 67.285 ;
        RECT 240.825 67.085 245.285 67.225 ;
        RECT 240.825 67.025 241.145 67.085 ;
        RECT 244.045 67.025 244.365 67.085 ;
        RECT 244.965 67.025 245.285 67.085 ;
        RECT 248.645 67.025 248.965 67.285 ;
        RECT 256.005 67.225 256.325 67.285 ;
        RECT 258.765 67.225 259.085 67.285 ;
        RECT 259.240 67.225 259.530 67.270 ;
        RECT 256.005 67.085 259.530 67.225 ;
        RECT 259.775 67.225 259.915 67.425 ;
        RECT 260.160 67.425 261.755 67.565 ;
        RECT 260.160 67.380 260.450 67.425 ;
        RECT 261.615 67.270 261.755 67.425 ;
        RECT 262.075 67.270 262.215 67.765 ;
        RECT 262.535 67.765 279.235 67.905 ;
        RECT 259.775 67.085 260.835 67.225 ;
        RECT 256.005 67.025 256.325 67.085 ;
        RECT 258.765 67.025 259.085 67.085 ;
        RECT 259.240 67.040 259.530 67.085 ;
        RECT 213.685 66.745 223.115 66.885 ;
        RECT 224.280 66.885 224.570 66.930 ;
        RECT 228.405 66.885 228.725 66.945 ;
        RECT 224.280 66.745 228.725 66.885 ;
        RECT 213.685 66.685 214.005 66.745 ;
        RECT 224.280 66.700 224.570 66.745 ;
        RECT 228.405 66.685 228.725 66.745 ;
        RECT 255.085 66.885 255.405 66.945 ;
        RECT 258.320 66.885 258.610 66.930 ;
        RECT 255.085 66.745 258.610 66.885 ;
        RECT 255.085 66.685 255.405 66.745 ;
        RECT 258.320 66.700 258.610 66.745 ;
        RECT 213.315 66.545 213.455 66.685 ;
        RECT 211.475 66.405 213.455 66.545 ;
        RECT 208.625 66.345 208.945 66.405 ;
        RECT 214.145 66.345 214.465 66.605 ;
        RECT 217.365 66.545 217.685 66.605 ;
        RECT 222.885 66.545 223.205 66.605 ;
        RECT 214.695 66.405 217.685 66.545 ;
        RECT 188.860 66.205 189.150 66.250 ;
        RECT 186.635 66.065 189.150 66.205 ;
        RECT 183.785 66.005 184.105 66.065 ;
        RECT 185.640 66.020 185.930 66.065 ;
        RECT 186.085 66.005 186.405 66.065 ;
        RECT 188.860 66.020 189.150 66.065 ;
        RECT 196.680 66.205 196.970 66.250 ;
        RECT 199.425 66.205 199.745 66.265 ;
        RECT 196.680 66.065 199.745 66.205 ;
        RECT 196.680 66.020 196.970 66.065 ;
        RECT 199.425 66.005 199.745 66.065 ;
        RECT 209.545 66.205 209.865 66.265 ;
        RECT 214.695 66.205 214.835 66.405 ;
        RECT 217.365 66.345 217.685 66.405 ;
        RECT 221.135 66.405 223.205 66.545 ;
        RECT 209.545 66.065 214.835 66.205 ;
        RECT 220.600 66.205 220.890 66.250 ;
        RECT 221.135 66.205 221.275 66.405 ;
        RECT 222.885 66.345 223.205 66.405 ;
        RECT 242.205 66.345 242.525 66.605 ;
        RECT 242.665 66.545 242.985 66.605 ;
        RECT 244.965 66.545 245.285 66.605 ;
        RECT 257.845 66.545 258.165 66.605 ;
        RECT 242.665 66.405 258.165 66.545 ;
        RECT 258.395 66.545 258.535 66.700 ;
        RECT 260.145 66.685 260.465 66.945 ;
        RECT 260.695 66.885 260.835 67.085 ;
        RECT 261.540 67.040 261.830 67.270 ;
        RECT 262.000 67.040 262.290 67.270 ;
        RECT 262.535 66.885 262.675 67.765 ;
        RECT 262.920 67.565 263.210 67.610 ;
        RECT 263.365 67.565 263.685 67.625 ;
        RECT 262.920 67.425 263.685 67.565 ;
        RECT 262.920 67.380 263.210 67.425 ;
        RECT 263.365 67.365 263.685 67.425 ;
        RECT 264.285 67.565 264.605 67.625 ;
        RECT 272.580 67.565 272.870 67.610 ;
        RECT 275.785 67.565 276.105 67.625 ;
        RECT 264.285 67.425 276.105 67.565 ;
        RECT 279.095 67.565 279.235 67.765 ;
        RECT 279.465 67.705 279.785 67.965 ;
        RECT 281.765 67.705 282.085 67.965 ;
        RECT 284.065 67.905 284.385 67.965 ;
        RECT 290.045 67.905 290.365 67.965 ;
        RECT 284.065 67.765 290.365 67.905 ;
        RECT 284.065 67.705 284.385 67.765 ;
        RECT 290.045 67.705 290.365 67.765 ;
        RECT 291.425 67.705 291.745 67.965 ;
        RECT 293.265 67.705 293.585 67.965 ;
        RECT 296.485 67.905 296.805 67.965 ;
        RECT 307.065 67.905 307.385 67.965 ;
        RECT 307.540 67.905 307.830 67.950 ;
        RECT 296.485 67.765 307.830 67.905 ;
        RECT 296.485 67.705 296.805 67.765 ;
        RECT 307.065 67.705 307.385 67.765 ;
        RECT 307.540 67.720 307.830 67.765 ;
        RECT 281.855 67.565 281.995 67.705 ;
        RECT 279.095 67.425 281.995 67.565 ;
        RECT 302.460 67.565 303.110 67.610 ;
        RECT 303.385 67.565 303.705 67.625 ;
        RECT 306.060 67.565 306.350 67.610 ;
        RECT 302.460 67.425 306.350 67.565 ;
        RECT 264.285 67.365 264.605 67.425 ;
        RECT 272.580 67.380 272.870 67.425 ;
        RECT 275.785 67.365 276.105 67.425 ;
        RECT 302.460 67.380 303.110 67.425 ;
        RECT 303.385 67.365 303.705 67.425 ;
        RECT 305.760 67.380 306.350 67.425 ;
        RECT 270.725 67.025 271.045 67.285 ;
        RECT 272.120 67.225 272.410 67.270 ;
        RECT 273.025 67.225 273.345 67.285 ;
        RECT 272.120 67.085 273.345 67.225 ;
        RECT 272.120 67.040 272.410 67.085 ;
        RECT 273.025 67.025 273.345 67.085 ;
        RECT 279.465 67.225 279.785 67.285 ;
        RECT 281.320 67.225 281.610 67.270 ;
        RECT 285.000 67.225 285.290 67.270 ;
        RECT 296.945 67.225 297.265 67.285 ;
        RECT 298.800 67.225 299.090 67.270 ;
        RECT 279.465 67.085 281.610 67.225 ;
        RECT 279.465 67.025 279.785 67.085 ;
        RECT 281.320 67.040 281.610 67.085 ;
        RECT 281.855 67.085 285.290 67.225 ;
        RECT 260.695 66.745 262.675 66.885 ;
        RECT 277.165 66.885 277.485 66.945 ;
        RECT 281.855 66.885 281.995 67.085 ;
        RECT 285.000 67.040 285.290 67.085 ;
        RECT 293.815 67.085 296.255 67.225 ;
        RECT 293.815 66.945 293.955 67.085 ;
        RECT 277.165 66.745 281.995 66.885 ;
        RECT 282.700 66.885 282.990 66.930 ;
        RECT 283.145 66.885 283.465 66.945 ;
        RECT 282.700 66.745 283.465 66.885 ;
        RECT 277.165 66.685 277.485 66.745 ;
        RECT 282.700 66.700 282.990 66.745 ;
        RECT 283.145 66.685 283.465 66.745 ;
        RECT 283.620 66.700 283.910 66.930 ;
        RECT 259.225 66.545 259.545 66.605 ;
        RECT 258.395 66.405 259.545 66.545 ;
        RECT 242.665 66.345 242.985 66.405 ;
        RECT 244.965 66.345 245.285 66.405 ;
        RECT 257.845 66.345 258.165 66.405 ;
        RECT 259.225 66.345 259.545 66.405 ;
        RECT 259.685 66.345 260.005 66.605 ;
        RECT 260.235 66.545 260.375 66.685 ;
        RECT 268.885 66.545 269.205 66.605 ;
        RECT 272.565 66.545 272.885 66.605 ;
        RECT 283.695 66.545 283.835 66.700 ;
        RECT 293.725 66.685 294.045 66.945 ;
        RECT 294.645 66.685 294.965 66.945 ;
        RECT 296.115 66.885 296.255 67.085 ;
        RECT 296.945 67.085 299.090 67.225 ;
        RECT 296.945 67.025 297.265 67.085 ;
        RECT 298.800 67.040 299.090 67.085 ;
        RECT 299.265 67.225 299.555 67.270 ;
        RECT 301.100 67.225 301.390 67.270 ;
        RECT 304.680 67.225 304.970 67.270 ;
        RECT 299.265 67.085 304.970 67.225 ;
        RECT 299.265 67.040 299.555 67.085 ;
        RECT 301.100 67.040 301.390 67.085 ;
        RECT 304.680 67.040 304.970 67.085 ;
        RECT 305.760 67.065 306.050 67.380 ;
        RECT 309.365 67.025 309.685 67.285 ;
        RECT 300.165 66.885 300.485 66.945 ;
        RECT 296.115 66.745 300.485 66.885 ;
        RECT 300.165 66.685 300.485 66.745 ;
        RECT 260.235 66.405 261.755 66.545 ;
        RECT 220.600 66.065 221.275 66.205 ;
        RECT 209.545 66.005 209.865 66.065 ;
        RECT 220.600 66.020 220.890 66.065 ;
        RECT 226.105 66.005 226.425 66.265 ;
        RECT 245.425 66.205 245.745 66.265 ;
        RECT 246.345 66.205 246.665 66.265 ;
        RECT 245.425 66.065 246.665 66.205 ;
        RECT 259.775 66.205 259.915 66.345 ;
        RECT 261.615 66.250 261.755 66.405 ;
        RECT 268.885 66.405 283.835 66.545 ;
        RECT 268.885 66.345 269.205 66.405 ;
        RECT 272.565 66.345 272.885 66.405 ;
        RECT 284.080 66.360 284.370 66.590 ;
        RECT 285.920 66.545 286.210 66.590 ;
        RECT 295.105 66.545 295.425 66.605 ;
        RECT 285.920 66.405 295.425 66.545 ;
        RECT 285.920 66.360 286.210 66.405 ;
        RECT 260.620 66.205 260.910 66.250 ;
        RECT 259.775 66.065 260.910 66.205 ;
        RECT 245.425 66.005 245.745 66.065 ;
        RECT 246.345 66.005 246.665 66.065 ;
        RECT 260.620 66.020 260.910 66.065 ;
        RECT 261.540 66.020 261.830 66.250 ;
        RECT 275.325 66.205 275.645 66.265 ;
        RECT 284.155 66.205 284.295 66.360 ;
        RECT 295.105 66.345 295.425 66.405 ;
        RECT 299.670 66.545 299.960 66.590 ;
        RECT 301.560 66.545 301.850 66.590 ;
        RECT 304.680 66.545 304.970 66.590 ;
        RECT 299.670 66.405 304.970 66.545 ;
        RECT 299.670 66.360 299.960 66.405 ;
        RECT 301.560 66.360 301.850 66.405 ;
        RECT 304.680 66.360 304.970 66.405 ;
        RECT 308.445 66.345 308.765 66.605 ;
        RECT 275.325 66.065 284.295 66.205 ;
        RECT 299.245 66.205 299.565 66.265 ;
        RECT 300.085 66.205 300.375 66.250 ;
        RECT 299.245 66.065 300.375 66.205 ;
        RECT 275.325 66.005 275.645 66.065 ;
        RECT 299.245 66.005 299.565 66.065 ;
        RECT 300.085 66.020 300.375 66.065 ;
        RECT 162.095 65.385 311.135 65.865 ;
        RECT 164.465 65.185 164.785 65.245 ;
        RECT 165.860 65.185 166.150 65.230 ;
        RECT 164.465 65.045 166.150 65.185 ;
        RECT 164.465 64.985 164.785 65.045 ;
        RECT 165.860 65.000 166.150 65.045 ;
        RECT 169.525 65.185 169.845 65.245 ;
        RECT 169.525 65.045 177.575 65.185 ;
        RECT 169.525 64.985 169.845 65.045 ;
        RECT 168.720 64.845 169.010 64.890 ;
        RECT 171.840 64.845 172.130 64.890 ;
        RECT 173.730 64.845 174.020 64.890 ;
        RECT 175.505 64.845 175.825 64.905 ;
        RECT 168.720 64.705 174.020 64.845 ;
        RECT 168.720 64.660 169.010 64.705 ;
        RECT 171.840 64.660 172.130 64.705 ;
        RECT 173.730 64.660 174.020 64.705 ;
        RECT 174.215 64.705 175.825 64.845 ;
        RECT 173.220 64.505 173.510 64.550 ;
        RECT 174.215 64.505 174.355 64.705 ;
        RECT 175.505 64.645 175.825 64.705 ;
        RECT 177.435 64.845 177.575 65.045 ;
        RECT 180.565 64.985 180.885 65.245 ;
        RECT 185.165 65.185 185.485 65.245 ;
        RECT 186.100 65.185 186.390 65.230 ;
        RECT 185.165 65.045 186.390 65.185 ;
        RECT 185.165 64.985 185.485 65.045 ;
        RECT 186.100 65.000 186.390 65.045 ;
        RECT 193.445 64.985 193.765 65.245 ;
        RECT 194.380 65.185 194.670 65.230 ;
        RECT 200.345 65.185 200.665 65.245 ;
        RECT 216.445 65.185 216.765 65.245 ;
        RECT 221.045 65.185 221.365 65.245 ;
        RECT 194.380 65.045 200.665 65.185 ;
        RECT 194.380 65.000 194.670 65.045 ;
        RECT 200.345 64.985 200.665 65.045 ;
        RECT 213.315 65.045 221.365 65.185 ;
        RECT 213.315 64.905 213.455 65.045 ;
        RECT 216.445 64.985 216.765 65.045 ;
        RECT 221.045 64.985 221.365 65.045 ;
        RECT 228.405 65.185 228.725 65.245 ;
        RECT 240.840 65.185 241.130 65.230 ;
        RECT 228.405 65.045 241.130 65.185 ;
        RECT 228.405 64.985 228.725 65.045 ;
        RECT 240.840 65.000 241.130 65.045 ;
        RECT 241.285 65.185 241.605 65.245 ;
        RECT 242.220 65.185 242.510 65.230 ;
        RECT 241.285 65.045 242.510 65.185 ;
        RECT 241.285 64.985 241.605 65.045 ;
        RECT 242.220 65.000 242.510 65.045 ;
        RECT 255.545 65.185 255.865 65.245 ;
        RECT 271.200 65.185 271.490 65.230 ;
        RECT 273.025 65.185 273.345 65.245 ;
        RECT 255.545 65.045 273.345 65.185 ;
        RECT 255.545 64.985 255.865 65.045 ;
        RECT 271.200 65.000 271.490 65.045 ;
        RECT 273.025 64.985 273.345 65.045 ;
        RECT 300.625 65.185 300.945 65.245 ;
        RECT 302.925 65.185 303.245 65.245 ;
        RECT 300.625 65.045 303.245 65.185 ;
        RECT 300.625 64.985 300.945 65.045 ;
        RECT 302.925 64.985 303.245 65.045 ;
        RECT 195.745 64.845 196.065 64.905 ;
        RECT 196.220 64.845 196.510 64.890 ;
        RECT 177.435 64.705 195.515 64.845 ;
        RECT 173.220 64.365 174.355 64.505 ;
        RECT 174.600 64.505 174.890 64.550 ;
        RECT 176.885 64.505 177.205 64.565 ;
        RECT 174.600 64.365 177.205 64.505 ;
        RECT 177.435 64.505 177.575 64.705 ;
        RECT 177.820 64.505 178.110 64.550 ;
        RECT 177.435 64.365 178.110 64.505 ;
        RECT 173.220 64.320 173.510 64.365 ;
        RECT 174.600 64.320 174.890 64.365 ;
        RECT 176.885 64.305 177.205 64.365 ;
        RECT 177.820 64.320 178.110 64.365 ;
        RECT 178.740 64.505 179.030 64.550 ;
        RECT 179.645 64.505 179.965 64.565 ;
        RECT 183.785 64.505 184.105 64.565 ;
        RECT 178.740 64.365 184.105 64.505 ;
        RECT 178.740 64.320 179.030 64.365 ;
        RECT 179.645 64.305 179.965 64.365 ;
        RECT 183.785 64.305 184.105 64.365 ;
        RECT 185.625 64.505 185.945 64.565 ;
        RECT 195.375 64.505 195.515 64.705 ;
        RECT 195.745 64.705 196.510 64.845 ;
        RECT 195.745 64.645 196.065 64.705 ;
        RECT 196.220 64.660 196.510 64.705 ;
        RECT 196.665 64.845 196.985 64.905 ;
        RECT 213.225 64.845 213.545 64.905 ;
        RECT 196.665 64.705 213.545 64.845 ;
        RECT 196.665 64.645 196.985 64.705 ;
        RECT 213.225 64.645 213.545 64.705 ;
        RECT 215.525 64.845 215.845 64.905 ;
        RECT 238.985 64.845 239.305 64.905 ;
        RECT 243.140 64.845 243.430 64.890 ;
        RECT 215.525 64.705 217.135 64.845 ;
        RECT 215.525 64.645 215.845 64.705 ;
        RECT 216.995 64.505 217.135 64.705 ;
        RECT 238.985 64.705 243.430 64.845 ;
        RECT 238.985 64.645 239.305 64.705 ;
        RECT 243.140 64.660 243.430 64.705 ;
        RECT 244.045 64.845 244.365 64.905 ;
        RECT 246.360 64.845 246.650 64.890 ;
        RECT 244.045 64.705 246.650 64.845 ;
        RECT 244.045 64.645 244.365 64.705 ;
        RECT 246.360 64.660 246.650 64.705 ;
        RECT 250.025 64.845 250.345 64.905 ;
        RECT 277.165 64.845 277.485 64.905 ;
        RECT 295.070 64.845 295.360 64.890 ;
        RECT 296.960 64.845 297.250 64.890 ;
        RECT 300.080 64.845 300.370 64.890 ;
        RECT 250.025 64.705 277.485 64.845 ;
        RECT 250.025 64.645 250.345 64.705 ;
        RECT 277.165 64.645 277.485 64.705 ;
        RECT 285.075 64.705 288.895 64.845 ;
        RECT 219.665 64.505 219.985 64.565 ;
        RECT 185.625 64.365 193.215 64.505 ;
        RECT 195.375 64.365 197.355 64.505 ;
        RECT 185.625 64.305 185.945 64.365 ;
        RECT 167.640 63.870 167.930 64.185 ;
        RECT 168.720 64.165 169.010 64.210 ;
        RECT 172.300 64.165 172.590 64.210 ;
        RECT 174.135 64.165 174.425 64.210 ;
        RECT 168.720 64.025 174.425 64.165 ;
        RECT 168.720 63.980 169.010 64.025 ;
        RECT 172.300 63.980 172.590 64.025 ;
        RECT 174.135 63.980 174.425 64.025 ;
        RECT 177.360 64.165 177.650 64.210 ;
        RECT 180.105 64.165 180.425 64.225 ;
        RECT 183.325 64.165 183.645 64.225 ;
        RECT 186.560 64.175 186.850 64.210 ;
        RECT 177.360 64.025 183.645 64.165 ;
        RECT 177.360 63.980 177.650 64.025 ;
        RECT 180.105 63.965 180.425 64.025 ;
        RECT 183.325 63.965 183.645 64.025 ;
        RECT 186.175 64.035 186.850 64.175 ;
        RECT 167.340 63.825 167.930 63.870 ;
        RECT 170.580 63.825 171.230 63.870 ;
        RECT 173.205 63.825 173.525 63.885 ;
        RECT 181.025 63.825 181.345 63.885 ;
        RECT 167.340 63.685 181.345 63.825 ;
        RECT 167.340 63.640 167.630 63.685 ;
        RECT 170.580 63.640 171.230 63.685 ;
        RECT 173.205 63.625 173.525 63.685 ;
        RECT 181.025 63.625 181.345 63.685 ;
        RECT 182.420 63.825 182.710 63.870 ;
        RECT 184.705 63.825 185.025 63.885 ;
        RECT 182.420 63.685 185.025 63.825 ;
        RECT 186.175 63.825 186.315 64.035 ;
        RECT 186.560 63.980 186.850 64.035 ;
        RECT 187.005 64.165 187.325 64.225 ;
        RECT 192.525 64.165 192.845 64.225 ;
        RECT 193.075 64.210 193.215 64.365 ;
        RECT 187.005 64.025 192.845 64.165 ;
        RECT 187.005 63.965 187.325 64.025 ;
        RECT 192.525 63.965 192.845 64.025 ;
        RECT 193.000 64.165 193.290 64.210 ;
        RECT 193.905 64.165 194.225 64.225 ;
        RECT 193.000 64.025 194.225 64.165 ;
        RECT 193.000 63.980 193.290 64.025 ;
        RECT 193.905 63.965 194.225 64.025 ;
        RECT 195.300 63.980 195.590 64.210 ;
        RECT 193.445 63.825 193.765 63.885 ;
        RECT 186.175 63.685 193.765 63.825 ;
        RECT 195.375 63.825 195.515 63.980 ;
        RECT 195.745 63.965 196.065 64.225 ;
        RECT 196.205 63.825 196.525 63.885 ;
        RECT 195.375 63.685 196.525 63.825 ;
        RECT 197.215 63.825 197.355 64.365 ;
        RECT 198.595 64.365 207.705 64.505 ;
        RECT 197.585 64.165 197.905 64.225 ;
        RECT 198.595 64.210 198.735 64.365 ;
        RECT 198.520 64.165 198.810 64.210 ;
        RECT 197.585 64.025 198.810 64.165 ;
        RECT 197.585 63.965 197.905 64.025 ;
        RECT 198.520 63.980 198.810 64.025 ;
        RECT 202.660 63.980 202.950 64.210 ;
        RECT 198.045 63.825 198.365 63.885 ;
        RECT 202.735 63.825 202.875 63.980 ;
        RECT 203.105 63.965 203.425 64.225 ;
        RECT 203.655 64.210 203.795 64.365 ;
        RECT 203.580 63.980 203.870 64.210 ;
        RECT 204.485 63.965 204.805 64.225 ;
        RECT 207.565 64.165 207.705 64.365 ;
        RECT 210.095 64.365 213.915 64.505 ;
        RECT 208.165 64.165 208.485 64.225 ;
        RECT 208.640 64.165 208.930 64.210 ;
        RECT 207.565 64.025 208.930 64.165 ;
        RECT 208.165 63.965 208.485 64.025 ;
        RECT 208.640 63.980 208.930 64.025 ;
        RECT 209.545 63.965 209.865 64.225 ;
        RECT 210.095 64.210 210.235 64.365 ;
        RECT 213.775 64.225 213.915 64.365 ;
        RECT 216.995 64.365 219.985 64.505 ;
        RECT 210.020 63.980 210.310 64.210 ;
        RECT 197.215 63.685 202.875 63.825 ;
        RECT 203.195 63.825 203.335 63.965 ;
        RECT 210.095 63.825 210.235 63.980 ;
        RECT 210.465 63.965 210.785 64.225 ;
        RECT 212.320 63.980 212.610 64.210 ;
        RECT 203.195 63.685 210.235 63.825 ;
        RECT 212.395 63.825 212.535 63.980 ;
        RECT 213.225 63.965 213.545 64.225 ;
        RECT 213.685 63.965 214.005 64.225 ;
        RECT 214.160 64.165 214.450 64.210 ;
        RECT 215.525 64.165 215.845 64.225 ;
        RECT 216.995 64.210 217.135 64.365 ;
        RECT 219.665 64.305 219.985 64.365 ;
        RECT 221.045 64.505 221.365 64.565 ;
        RECT 221.520 64.505 221.810 64.550 ;
        RECT 221.045 64.365 221.810 64.505 ;
        RECT 221.045 64.305 221.365 64.365 ;
        RECT 221.520 64.320 221.810 64.365 ;
        RECT 236.685 64.505 237.005 64.565 ;
        RECT 279.465 64.505 279.785 64.565 ;
        RECT 236.685 64.365 279.785 64.505 ;
        RECT 236.685 64.305 237.005 64.365 ;
        RECT 279.465 64.305 279.785 64.365 ;
        RECT 279.925 64.505 280.245 64.565 ;
        RECT 285.075 64.550 285.215 64.705 ;
        RECT 288.755 64.550 288.895 64.705 ;
        RECT 295.070 64.705 300.370 64.845 ;
        RECT 295.070 64.660 295.360 64.705 ;
        RECT 296.960 64.660 297.250 64.705 ;
        RECT 300.080 64.660 300.370 64.705 ;
        RECT 285.000 64.505 285.290 64.550 ;
        RECT 279.925 64.365 285.290 64.505 ;
        RECT 279.925 64.305 280.245 64.365 ;
        RECT 285.000 64.320 285.290 64.365 ;
        RECT 288.680 64.320 288.970 64.550 ;
        RECT 214.160 64.025 215.845 64.165 ;
        RECT 214.160 63.980 214.450 64.025 ;
        RECT 215.525 63.965 215.845 64.025 ;
        RECT 216.000 63.980 216.290 64.210 ;
        RECT 216.920 63.980 217.210 64.210 ;
        RECT 216.105 63.825 216.245 63.980 ;
        RECT 217.365 63.965 217.685 64.225 ;
        RECT 217.940 64.175 218.230 64.210 ;
        RECT 218.745 64.175 219.065 64.225 ;
        RECT 217.940 64.035 219.065 64.175 ;
        RECT 217.940 63.980 218.230 64.035 ;
        RECT 218.745 63.965 219.065 64.035 ;
        RECT 220.585 64.165 220.905 64.225 ;
        RECT 226.105 64.165 226.425 64.225 ;
        RECT 220.585 64.025 226.425 64.165 ;
        RECT 220.585 63.965 220.905 64.025 ;
        RECT 226.105 63.965 226.425 64.025 ;
        RECT 242.665 63.965 242.985 64.225 ;
        RECT 244.520 64.165 244.810 64.210 ;
        RECT 244.965 64.165 245.285 64.225 ;
        RECT 244.520 64.025 245.285 64.165 ;
        RECT 244.520 63.980 244.810 64.025 ;
        RECT 244.965 63.965 245.285 64.025 ;
        RECT 245.425 64.165 245.745 64.225 ;
        RECT 260.145 64.165 260.465 64.225 ;
        RECT 245.425 64.025 260.465 64.165 ;
        RECT 245.425 63.965 245.745 64.025 ;
        RECT 260.145 63.965 260.465 64.025 ;
        RECT 272.565 63.965 272.885 64.225 ;
        RECT 283.620 64.165 283.910 64.210 ;
        RECT 289.585 64.165 289.905 64.225 ;
        RECT 294.200 64.165 294.490 64.210 ;
        RECT 283.620 64.025 288.895 64.165 ;
        RECT 283.620 63.980 283.910 64.025 ;
        RECT 236.225 63.825 236.545 63.885 ;
        RECT 254.165 63.825 254.485 63.885 ;
        RECT 212.395 63.685 236.545 63.825 ;
        RECT 182.420 63.640 182.710 63.685 ;
        RECT 184.705 63.625 185.025 63.685 ;
        RECT 187.095 63.545 187.235 63.685 ;
        RECT 193.445 63.625 193.765 63.685 ;
        RECT 196.205 63.625 196.525 63.685 ;
        RECT 198.045 63.625 198.365 63.685 ;
        RECT 236.225 63.625 236.545 63.685 ;
        RECT 244.135 63.685 254.485 63.825 ;
        RECT 175.520 63.485 175.810 63.530 ;
        RECT 176.425 63.485 176.745 63.545 ;
        RECT 175.520 63.345 176.745 63.485 ;
        RECT 175.520 63.300 175.810 63.345 ;
        RECT 176.425 63.285 176.745 63.345 ;
        RECT 182.880 63.485 183.170 63.530 ;
        RECT 186.085 63.485 186.405 63.545 ;
        RECT 182.880 63.345 186.405 63.485 ;
        RECT 182.880 63.300 183.170 63.345 ;
        RECT 186.085 63.285 186.405 63.345 ;
        RECT 187.005 63.285 187.325 63.545 ;
        RECT 195.745 63.485 196.065 63.545 ;
        RECT 196.665 63.485 196.985 63.545 ;
        RECT 195.745 63.345 196.985 63.485 ;
        RECT 195.745 63.285 196.065 63.345 ;
        RECT 196.665 63.285 196.985 63.345 ;
        RECT 201.265 63.285 201.585 63.545 ;
        RECT 211.845 63.285 212.165 63.545 ;
        RECT 215.540 63.485 215.830 63.530 ;
        RECT 216.445 63.485 216.765 63.545 ;
        RECT 215.540 63.345 216.765 63.485 ;
        RECT 215.540 63.300 215.830 63.345 ;
        RECT 216.445 63.285 216.765 63.345 ;
        RECT 219.205 63.285 219.525 63.545 ;
        RECT 219.665 63.285 219.985 63.545 ;
        RECT 244.135 63.530 244.275 63.685 ;
        RECT 254.165 63.625 254.485 63.685 ;
        RECT 259.225 63.825 259.545 63.885 ;
        RECT 270.280 63.825 270.570 63.870 ;
        RECT 270.725 63.825 271.045 63.885 ;
        RECT 259.225 63.685 271.045 63.825 ;
        RECT 259.225 63.625 259.545 63.685 ;
        RECT 270.280 63.640 270.570 63.685 ;
        RECT 270.725 63.625 271.045 63.685 ;
        RECT 280.845 63.825 281.165 63.885 ;
        RECT 288.205 63.825 288.525 63.885 ;
        RECT 280.845 63.685 288.525 63.825 ;
        RECT 288.755 63.825 288.895 64.025 ;
        RECT 289.585 64.025 294.490 64.165 ;
        RECT 289.585 63.965 289.905 64.025 ;
        RECT 294.200 63.980 294.490 64.025 ;
        RECT 294.665 64.165 294.955 64.210 ;
        RECT 296.500 64.165 296.790 64.210 ;
        RECT 300.080 64.165 300.370 64.210 ;
        RECT 294.665 64.025 300.370 64.165 ;
        RECT 294.665 63.980 294.955 64.025 ;
        RECT 296.500 63.980 296.790 64.025 ;
        RECT 300.080 63.980 300.370 64.025 ;
        RECT 290.965 63.825 291.285 63.885 ;
        RECT 288.755 63.685 291.285 63.825 ;
        RECT 280.845 63.625 281.165 63.685 ;
        RECT 288.205 63.625 288.525 63.685 ;
        RECT 290.965 63.625 291.285 63.685 ;
        RECT 295.565 63.625 295.885 63.885 ;
        RECT 297.860 63.825 298.510 63.870 ;
        RECT 298.785 63.825 299.105 63.885 ;
        RECT 301.160 63.870 301.450 64.185 ;
        RECT 301.160 63.825 301.750 63.870 ;
        RECT 297.860 63.685 301.750 63.825 ;
        RECT 297.860 63.640 298.510 63.685 ;
        RECT 298.785 63.625 299.105 63.685 ;
        RECT 301.460 63.640 301.750 63.685 ;
        RECT 244.060 63.300 244.350 63.530 ;
        RECT 246.805 63.485 247.125 63.545 ;
        RECT 257.385 63.485 257.705 63.545 ;
        RECT 269.805 63.485 270.125 63.545 ;
        RECT 271.200 63.485 271.490 63.530 ;
        RECT 246.805 63.345 271.490 63.485 ;
        RECT 246.805 63.285 247.125 63.345 ;
        RECT 257.385 63.285 257.705 63.345 ;
        RECT 269.805 63.285 270.125 63.345 ;
        RECT 271.200 63.300 271.490 63.345 ;
        RECT 281.765 63.285 282.085 63.545 ;
        RECT 284.065 63.285 284.385 63.545 ;
        RECT 284.985 63.485 285.305 63.545 ;
        RECT 285.920 63.485 286.210 63.530 ;
        RECT 284.985 63.345 286.210 63.485 ;
        RECT 284.985 63.285 285.305 63.345 ;
        RECT 285.920 63.300 286.210 63.345 ;
        RECT 287.745 63.485 288.065 63.545 ;
        RECT 292.345 63.485 292.665 63.545 ;
        RECT 309.825 63.485 310.145 63.545 ;
        RECT 287.745 63.345 310.145 63.485 ;
        RECT 287.745 63.285 288.065 63.345 ;
        RECT 292.345 63.285 292.665 63.345 ;
        RECT 309.825 63.285 310.145 63.345 ;
        RECT 162.095 62.665 311.135 63.145 ;
        RECT 169.065 62.465 169.385 62.525 ;
        RECT 169.540 62.465 169.830 62.510 ;
        RECT 169.065 62.325 169.830 62.465 ;
        RECT 169.065 62.265 169.385 62.325 ;
        RECT 169.540 62.280 169.830 62.325 ;
        RECT 175.965 62.465 176.285 62.525 ;
        RECT 179.200 62.465 179.490 62.510 ;
        RECT 175.965 62.325 179.490 62.465 ;
        RECT 175.965 62.265 176.285 62.325 ;
        RECT 179.200 62.280 179.490 62.325 ;
        RECT 184.705 62.465 185.025 62.525 ;
        RECT 185.640 62.465 185.930 62.510 ;
        RECT 184.705 62.325 185.930 62.465 ;
        RECT 184.705 62.265 185.025 62.325 ;
        RECT 185.640 62.280 185.930 62.325 ;
        RECT 189.765 62.465 190.085 62.525 ;
        RECT 191.620 62.465 191.910 62.510 ;
        RECT 189.765 62.325 191.910 62.465 ;
        RECT 189.765 62.265 190.085 62.325 ;
        RECT 191.620 62.280 191.910 62.325 ;
        RECT 195.285 62.265 195.605 62.525 ;
        RECT 215.525 62.465 215.845 62.525 ;
        RECT 218.745 62.465 219.065 62.525 ;
        RECT 195.835 62.325 219.065 62.465 ;
        RECT 171.020 62.125 171.310 62.170 ;
        RECT 173.205 62.125 173.525 62.185 ;
        RECT 174.260 62.125 174.910 62.170 ;
        RECT 171.020 61.985 174.910 62.125 ;
        RECT 171.020 61.940 171.610 61.985 ;
        RECT 164.940 61.600 165.230 61.830 ;
        RECT 171.320 61.625 171.610 61.940 ;
        RECT 173.205 61.925 173.525 61.985 ;
        RECT 174.260 61.940 174.910 61.985 ;
        RECT 176.885 62.125 177.205 62.185 ;
        RECT 187.925 62.125 188.245 62.185 ;
        RECT 190.700 62.125 190.990 62.170 ;
        RECT 176.885 61.985 178.495 62.125 ;
        RECT 176.885 61.925 177.205 61.985 ;
        RECT 178.355 61.830 178.495 61.985 ;
        RECT 187.925 61.985 190.990 62.125 ;
        RECT 187.925 61.925 188.245 61.985 ;
        RECT 190.700 61.940 190.990 61.985 ;
        RECT 172.400 61.785 172.690 61.830 ;
        RECT 175.980 61.785 176.270 61.830 ;
        RECT 177.815 61.785 178.105 61.830 ;
        RECT 172.400 61.645 178.105 61.785 ;
        RECT 172.400 61.600 172.690 61.645 ;
        RECT 175.980 61.600 176.270 61.645 ;
        RECT 177.815 61.600 178.105 61.645 ;
        RECT 178.280 61.600 178.570 61.830 ;
        RECT 180.120 61.785 180.410 61.830 ;
        RECT 186.545 61.785 186.865 61.845 ;
        RECT 180.120 61.645 186.865 61.785 ;
        RECT 180.120 61.600 180.410 61.645 ;
        RECT 165.015 61.445 165.155 61.600 ;
        RECT 186.545 61.585 186.865 61.645 ;
        RECT 187.465 61.585 187.785 61.845 ;
        RECT 188.385 61.785 188.705 61.845 ;
        RECT 192.540 61.785 192.830 61.830 ;
        RECT 188.385 61.645 192.830 61.785 ;
        RECT 188.385 61.585 188.705 61.645 ;
        RECT 192.540 61.600 192.830 61.645 ;
        RECT 175.045 61.445 175.365 61.505 ;
        RECT 165.015 61.305 175.365 61.445 ;
        RECT 175.045 61.245 175.365 61.305 ;
        RECT 176.425 61.445 176.745 61.505 ;
        RECT 176.900 61.445 177.190 61.490 ;
        RECT 176.425 61.305 177.190 61.445 ;
        RECT 176.425 61.245 176.745 61.305 ;
        RECT 176.900 61.260 177.190 61.305 ;
        RECT 181.025 61.445 181.345 61.505 ;
        RECT 184.245 61.445 184.565 61.505 ;
        RECT 181.025 61.305 184.565 61.445 ;
        RECT 181.025 61.245 181.345 61.305 ;
        RECT 184.245 61.245 184.565 61.305 ;
        RECT 186.085 61.445 186.405 61.505 ;
        RECT 186.085 61.305 189.535 61.445 ;
        RECT 186.085 61.245 186.405 61.305 ;
        RECT 172.400 61.105 172.690 61.150 ;
        RECT 175.520 61.105 175.810 61.150 ;
        RECT 177.410 61.105 177.700 61.150 ;
        RECT 187.005 61.105 187.325 61.165 ;
        RECT 172.400 60.965 177.700 61.105 ;
        RECT 172.400 60.920 172.690 60.965 ;
        RECT 175.520 60.920 175.810 60.965 ;
        RECT 177.410 60.920 177.700 60.965 ;
        RECT 177.895 60.965 187.325 61.105 ;
        RECT 164.005 60.565 164.325 60.825 ;
        RECT 175.965 60.765 176.285 60.825 ;
        RECT 177.895 60.765 178.035 60.965 ;
        RECT 187.005 60.905 187.325 60.965 ;
        RECT 188.845 60.905 189.165 61.165 ;
        RECT 189.395 61.105 189.535 61.305 ;
        RECT 189.765 61.245 190.085 61.505 ;
        RECT 192.065 61.445 192.385 61.505 ;
        RECT 193.000 61.445 193.290 61.490 ;
        RECT 195.835 61.445 195.975 62.325 ;
        RECT 215.525 62.265 215.845 62.325 ;
        RECT 218.745 62.265 219.065 62.325 ;
        RECT 231.165 62.465 231.485 62.525 ;
        RECT 232.560 62.465 232.850 62.510 ;
        RECT 231.165 62.325 232.850 62.465 ;
        RECT 231.165 62.265 231.485 62.325 ;
        RECT 232.560 62.280 232.850 62.325 ;
        RECT 242.665 62.465 242.985 62.525 ;
        RECT 243.600 62.465 243.890 62.510 ;
        RECT 242.665 62.325 243.890 62.465 ;
        RECT 242.665 62.265 242.985 62.325 ;
        RECT 243.600 62.280 243.890 62.325 ;
        RECT 251.405 62.265 251.725 62.525 ;
        RECT 253.260 62.465 253.550 62.510 ;
        RECT 258.765 62.465 259.085 62.525 ;
        RECT 253.260 62.325 259.085 62.465 ;
        RECT 253.260 62.280 253.550 62.325 ;
        RECT 258.765 62.265 259.085 62.325 ;
        RECT 259.225 62.510 259.545 62.525 ;
        RECT 259.225 62.465 259.575 62.510 ;
        RECT 262.000 62.465 262.290 62.510 ;
        RECT 262.905 62.465 263.225 62.525 ;
        RECT 279.005 62.465 279.325 62.525 ;
        RECT 259.225 62.325 259.740 62.465 ;
        RECT 262.000 62.325 279.325 62.465 ;
        RECT 259.225 62.280 259.575 62.325 ;
        RECT 262.000 62.280 262.290 62.325 ;
        RECT 259.225 62.265 259.545 62.280 ;
        RECT 262.905 62.265 263.225 62.325 ;
        RECT 279.005 62.265 279.325 62.325 ;
        RECT 279.925 62.265 280.245 62.525 ;
        RECT 288.205 62.465 288.525 62.525 ;
        RECT 296.025 62.465 296.345 62.525 ;
        RECT 288.205 62.325 296.345 62.465 ;
        RECT 288.205 62.265 288.525 62.325 ;
        RECT 296.025 62.265 296.345 62.325 ;
        RECT 296.485 62.265 296.805 62.525 ;
        RECT 298.340 62.465 298.630 62.510 ;
        RECT 299.245 62.465 299.565 62.525 ;
        RECT 298.340 62.325 299.565 62.465 ;
        RECT 298.340 62.280 298.630 62.325 ;
        RECT 299.245 62.265 299.565 62.325 ;
        RECT 300.165 62.465 300.485 62.525 ;
        RECT 301.100 62.465 301.390 62.510 ;
        RECT 300.165 62.325 301.390 62.465 ;
        RECT 300.165 62.265 300.485 62.325 ;
        RECT 301.100 62.280 301.390 62.325 ;
        RECT 305.225 62.265 305.545 62.525 ;
        RECT 219.205 62.125 219.525 62.185 ;
        RECT 230.245 62.125 230.565 62.185 ;
        RECT 236.685 62.125 237.005 62.185 ;
        RECT 212.395 61.985 218.055 62.125 ;
        RECT 212.395 61.845 212.535 61.985 ;
        RECT 198.060 61.600 198.350 61.830 ;
        RECT 192.065 61.305 193.290 61.445 ;
        RECT 192.065 61.245 192.385 61.305 ;
        RECT 193.000 61.260 193.290 61.305 ;
        RECT 193.535 61.305 195.975 61.445 ;
        RECT 198.135 61.445 198.275 61.600 ;
        RECT 198.505 61.585 198.825 61.845 ;
        RECT 198.965 61.585 199.285 61.845 ;
        RECT 199.425 61.585 199.745 61.845 ;
        RECT 200.345 61.585 200.665 61.845 ;
        RECT 210.005 61.585 210.325 61.845 ;
        RECT 210.925 61.585 211.245 61.845 ;
        RECT 212.305 61.585 212.625 61.845 ;
        RECT 215.525 61.585 215.845 61.845 ;
        RECT 215.985 61.785 216.305 61.845 ;
        RECT 216.460 61.785 216.750 61.830 ;
        RECT 215.985 61.645 216.750 61.785 ;
        RECT 215.985 61.585 216.305 61.645 ;
        RECT 216.460 61.600 216.750 61.645 ;
        RECT 216.905 61.585 217.225 61.845 ;
        RECT 217.915 61.830 218.055 61.985 ;
        RECT 219.205 61.985 221.735 62.125 ;
        RECT 219.205 61.925 219.525 61.985 ;
        RECT 221.595 61.830 221.735 61.985 ;
        RECT 230.245 61.985 237.005 62.125 ;
        RECT 230.245 61.925 230.565 61.985 ;
        RECT 236.685 61.925 237.005 61.985 ;
        RECT 244.045 62.125 244.365 62.185 ;
        RECT 256.925 62.125 257.245 62.185 ;
        RECT 261.080 62.125 261.370 62.170 ;
        RECT 244.045 61.985 247.035 62.125 ;
        RECT 244.045 61.925 244.365 61.985 ;
        RECT 246.895 61.845 247.035 61.985 ;
        RECT 248.735 61.985 254.855 62.125 ;
        RECT 248.735 61.845 248.875 61.985 ;
        RECT 217.840 61.785 218.130 61.830 ;
        RECT 221.060 61.785 221.350 61.830 ;
        RECT 217.840 61.645 221.350 61.785 ;
        RECT 217.840 61.600 218.130 61.645 ;
        RECT 204.025 61.445 204.345 61.505 ;
        RECT 198.135 61.305 204.345 61.445 ;
        RECT 193.535 61.105 193.675 61.305 ;
        RECT 204.025 61.245 204.345 61.305 ;
        RECT 209.085 61.445 209.405 61.505 ;
        RECT 210.480 61.445 210.770 61.490 ;
        RECT 209.085 61.305 210.770 61.445 ;
        RECT 209.085 61.245 209.405 61.305 ;
        RECT 210.480 61.260 210.770 61.305 ;
        RECT 211.400 61.445 211.690 61.490 ;
        RECT 219.665 61.445 219.985 61.505 ;
        RECT 211.400 61.305 219.985 61.445 ;
        RECT 211.400 61.260 211.690 61.305 ;
        RECT 219.665 61.245 219.985 61.305 ;
        RECT 189.395 60.965 193.675 61.105 ;
        RECT 194.840 61.105 195.130 61.150 ;
        RECT 196.205 61.105 196.525 61.165 ;
        RECT 194.840 60.965 196.525 61.105 ;
        RECT 194.840 60.920 195.130 60.965 ;
        RECT 196.205 60.905 196.525 60.965 ;
        RECT 214.160 61.105 214.450 61.150 ;
        RECT 216.445 61.105 216.765 61.165 ;
        RECT 214.160 60.965 216.765 61.105 ;
        RECT 214.160 60.920 214.450 60.965 ;
        RECT 216.445 60.905 216.765 60.965 ;
        RECT 216.905 61.105 217.225 61.165 ;
        RECT 220.215 61.105 220.355 61.645 ;
        RECT 221.060 61.600 221.350 61.645 ;
        RECT 221.520 61.600 221.810 61.830 ;
        RECT 222.425 61.585 222.745 61.845 ;
        RECT 231.625 61.785 231.945 61.845 ;
        RECT 232.100 61.785 232.390 61.830 ;
        RECT 234.845 61.785 235.165 61.845 ;
        RECT 231.625 61.645 235.165 61.785 ;
        RECT 231.625 61.585 231.945 61.645 ;
        RECT 232.100 61.600 232.390 61.645 ;
        RECT 234.845 61.585 235.165 61.645 ;
        RECT 236.240 61.785 236.530 61.830 ;
        RECT 239.920 61.785 240.210 61.830 ;
        RECT 245.440 61.785 245.730 61.830 ;
        RECT 236.240 61.645 240.210 61.785 ;
        RECT 236.240 61.600 236.530 61.645 ;
        RECT 239.920 61.600 240.210 61.645 ;
        RECT 242.755 61.645 245.730 61.785 ;
        RECT 221.980 61.445 222.270 61.490 ;
        RECT 223.805 61.445 224.125 61.505 ;
        RECT 221.980 61.305 224.125 61.445 ;
        RECT 221.980 61.260 222.270 61.305 ;
        RECT 223.805 61.245 224.125 61.305 ;
        RECT 225.185 61.445 225.505 61.505 ;
        RECT 226.580 61.445 226.870 61.490 ;
        RECT 225.185 61.305 226.870 61.445 ;
        RECT 225.185 61.245 225.505 61.305 ;
        RECT 226.580 61.260 226.870 61.305 ;
        RECT 233.480 61.260 233.770 61.490 ;
        RECT 237.160 61.260 237.450 61.490 ;
        RECT 238.525 61.445 238.845 61.505 ;
        RECT 241.285 61.445 241.605 61.505 ;
        RECT 242.755 61.490 242.895 61.645 ;
        RECT 245.440 61.600 245.730 61.645 ;
        RECT 246.805 61.585 247.125 61.845 ;
        RECT 247.265 61.585 247.585 61.845 ;
        RECT 248.645 61.585 248.965 61.845 ;
        RECT 250.025 61.585 250.345 61.845 ;
        RECT 253.705 61.585 254.025 61.845 ;
        RECT 244.505 61.490 244.825 61.505 ;
        RECT 242.680 61.445 242.970 61.490 ;
        RECT 238.525 61.305 242.970 61.445 ;
        RECT 216.905 60.965 220.355 61.105 ;
        RECT 233.555 61.105 233.695 61.260 ;
        RECT 237.235 61.105 237.375 61.260 ;
        RECT 238.525 61.245 238.845 61.305 ;
        RECT 241.285 61.245 241.605 61.305 ;
        RECT 242.680 61.260 242.970 61.305 ;
        RECT 244.395 61.260 244.825 61.490 ;
        RECT 244.505 61.245 244.825 61.260 ;
        RECT 244.965 61.445 245.285 61.505 ;
        RECT 248.185 61.445 248.505 61.505 ;
        RECT 244.965 61.305 248.505 61.445 ;
        RECT 244.965 61.245 245.285 61.305 ;
        RECT 248.185 61.245 248.505 61.305 ;
        RECT 254.180 61.260 254.470 61.490 ;
        RECT 254.715 61.445 254.855 61.985 ;
        RECT 256.925 61.985 261.370 62.125 ;
        RECT 256.925 61.925 257.245 61.985 ;
        RECT 261.080 61.940 261.370 61.985 ;
        RECT 281.765 61.925 282.085 62.185 ;
        RECT 284.060 62.125 284.710 62.170 ;
        RECT 287.660 62.125 287.950 62.170 ;
        RECT 284.060 61.985 287.950 62.125 ;
        RECT 284.060 61.940 284.710 61.985 ;
        RECT 287.360 61.940 287.950 61.985 ;
        RECT 300.640 62.125 300.930 62.170 ;
        RECT 302.925 62.125 303.245 62.185 ;
        RECT 300.640 61.985 303.245 62.125 ;
        RECT 300.640 61.940 300.930 61.985 ;
        RECT 287.360 61.845 287.650 61.940 ;
        RECT 302.925 61.925 303.245 61.985 ;
        RECT 257.385 61.585 257.705 61.845 ;
        RECT 260.145 61.785 260.465 61.845 ;
        RECT 262.445 61.785 262.765 61.845 ;
        RECT 260.145 61.645 262.765 61.785 ;
        RECT 260.145 61.585 260.465 61.645 ;
        RECT 262.445 61.585 262.765 61.645 ;
        RECT 262.905 61.785 263.225 61.845 ;
        RECT 269.345 61.785 269.665 61.845 ;
        RECT 262.905 61.645 269.665 61.785 ;
        RECT 262.905 61.585 263.225 61.645 ;
        RECT 269.345 61.585 269.665 61.645 ;
        RECT 277.165 61.785 277.485 61.845 ;
        RECT 279.020 61.785 279.310 61.830 ;
        RECT 277.165 61.645 279.310 61.785 ;
        RECT 277.165 61.585 277.485 61.645 ;
        RECT 279.020 61.600 279.310 61.645 ;
        RECT 280.865 61.785 281.155 61.830 ;
        RECT 282.700 61.785 282.990 61.830 ;
        RECT 286.280 61.785 286.570 61.830 ;
        RECT 280.865 61.645 286.570 61.785 ;
        RECT 280.865 61.600 281.155 61.645 ;
        RECT 282.700 61.600 282.990 61.645 ;
        RECT 286.280 61.600 286.570 61.645 ;
        RECT 287.285 61.625 287.650 61.845 ;
        RECT 304.765 61.785 305.085 61.845 ;
        RECT 306.145 61.785 306.465 61.845 ;
        RECT 304.765 61.645 306.465 61.785 ;
        RECT 287.285 61.585 287.605 61.625 ;
        RECT 304.765 61.585 305.085 61.645 ;
        RECT 306.145 61.585 306.465 61.645 ;
        RECT 275.325 61.445 275.645 61.505 ;
        RECT 277.640 61.445 277.930 61.490 ;
        RECT 254.715 61.305 277.930 61.445 ;
        RECT 249.565 61.105 249.885 61.165 ;
        RECT 250.960 61.105 251.250 61.150 ;
        RECT 254.255 61.105 254.395 61.260 ;
        RECT 275.325 61.245 275.645 61.305 ;
        RECT 277.640 61.260 277.930 61.305 ;
        RECT 278.085 61.245 278.405 61.505 ;
        RECT 280.400 61.445 280.690 61.490 ;
        RECT 289.140 61.445 289.430 61.490 ;
        RECT 290.965 61.445 291.285 61.505 ;
        RECT 280.400 61.305 281.075 61.445 ;
        RECT 280.400 61.260 280.690 61.305 ;
        RECT 256.005 61.105 256.325 61.165 ;
        RECT 260.160 61.105 260.450 61.150 ;
        RECT 233.555 60.965 254.395 61.105 ;
        RECT 254.715 60.965 260.450 61.105 ;
        RECT 216.905 60.905 217.225 60.965 ;
        RECT 249.565 60.905 249.885 60.965 ;
        RECT 250.960 60.920 251.250 60.965 ;
        RECT 175.965 60.625 178.035 60.765 ;
        RECT 180.565 60.765 180.885 60.825 ;
        RECT 184.705 60.765 185.025 60.825 ;
        RECT 180.565 60.625 185.025 60.765 ;
        RECT 175.965 60.565 176.285 60.625 ;
        RECT 180.565 60.565 180.885 60.625 ;
        RECT 184.705 60.565 185.025 60.625 ;
        RECT 186.085 60.765 186.405 60.825 ;
        RECT 188.935 60.765 189.075 60.905 ;
        RECT 186.085 60.625 189.075 60.765 ;
        RECT 186.085 60.565 186.405 60.625 ;
        RECT 196.665 60.565 196.985 60.825 ;
        RECT 205.865 60.765 206.185 60.825 ;
        RECT 208.640 60.765 208.930 60.810 ;
        RECT 205.865 60.625 208.930 60.765 ;
        RECT 205.865 60.565 206.185 60.625 ;
        RECT 208.640 60.580 208.930 60.625 ;
        RECT 216.000 60.765 216.290 60.810 ;
        RECT 217.825 60.765 218.145 60.825 ;
        RECT 216.000 60.625 218.145 60.765 ;
        RECT 216.000 60.580 216.290 60.625 ;
        RECT 217.825 60.565 218.145 60.625 ;
        RECT 220.125 60.565 220.445 60.825 ;
        RECT 223.805 60.565 224.125 60.825 ;
        RECT 230.245 60.565 230.565 60.825 ;
        RECT 233.925 60.765 234.245 60.825 ;
        RECT 234.400 60.765 234.690 60.810 ;
        RECT 233.925 60.625 234.690 60.765 ;
        RECT 233.925 60.565 234.245 60.625 ;
        RECT 234.400 60.580 234.690 60.625 ;
        RECT 248.185 60.565 248.505 60.825 ;
        RECT 249.120 60.765 249.410 60.810 ;
        RECT 254.715 60.765 254.855 60.965 ;
        RECT 256.005 60.905 256.325 60.965 ;
        RECT 260.160 60.920 260.450 60.965 ;
        RECT 263.825 60.905 264.145 61.165 ;
        RECT 272.105 61.105 272.425 61.165 ;
        RECT 278.175 61.105 278.315 61.245 ;
        RECT 272.105 60.965 278.315 61.105 ;
        RECT 272.105 60.905 272.425 60.965 ;
        RECT 249.120 60.625 254.855 60.765 ;
        RECT 255.545 60.765 255.865 60.825 ;
        RECT 259.240 60.765 259.530 60.810 ;
        RECT 255.545 60.625 259.530 60.765 ;
        RECT 280.935 60.765 281.075 61.305 ;
        RECT 289.140 61.305 291.285 61.445 ;
        RECT 289.140 61.260 289.430 61.305 ;
        RECT 290.965 61.245 291.285 61.305 ;
        RECT 295.105 61.445 295.425 61.505 ;
        RECT 295.105 61.305 300.855 61.445 ;
        RECT 295.105 61.245 295.425 61.305 ;
        RECT 281.270 61.105 281.560 61.150 ;
        RECT 283.160 61.105 283.450 61.150 ;
        RECT 286.280 61.105 286.570 61.150 ;
        RECT 281.270 60.965 286.570 61.105 ;
        RECT 281.270 60.920 281.560 60.965 ;
        RECT 283.160 60.920 283.450 60.965 ;
        RECT 286.280 60.920 286.570 60.965 ;
        RECT 295.565 61.105 295.885 61.165 ;
        RECT 298.800 61.105 299.090 61.150 ;
        RECT 295.565 60.965 299.090 61.105 ;
        RECT 300.715 61.105 300.855 61.305 ;
        RECT 301.560 61.260 301.850 61.490 ;
        RECT 305.700 61.260 305.990 61.490 ;
        RECT 301.635 61.105 301.775 61.260 ;
        RECT 303.845 61.105 304.165 61.165 ;
        RECT 305.775 61.105 305.915 61.260 ;
        RECT 300.715 60.965 305.915 61.105 ;
        RECT 295.565 60.905 295.885 60.965 ;
        RECT 298.800 60.920 299.090 60.965 ;
        RECT 303.845 60.905 304.165 60.965 ;
        RECT 283.605 60.765 283.925 60.825 ;
        RECT 280.935 60.625 283.925 60.765 ;
        RECT 249.120 60.580 249.410 60.625 ;
        RECT 255.545 60.565 255.865 60.625 ;
        RECT 259.240 60.580 259.530 60.625 ;
        RECT 283.605 60.565 283.925 60.625 ;
        RECT 302.005 60.765 302.325 60.825 ;
        RECT 302.940 60.765 303.230 60.810 ;
        RECT 302.005 60.625 303.230 60.765 ;
        RECT 302.005 60.565 302.325 60.625 ;
        RECT 302.940 60.580 303.230 60.625 ;
        RECT 162.095 59.945 311.135 60.425 ;
        RECT 178.280 59.745 178.570 59.790 ;
        RECT 180.105 59.745 180.425 59.805 ;
        RECT 178.280 59.605 180.425 59.745 ;
        RECT 178.280 59.560 178.570 59.605 ;
        RECT 180.105 59.545 180.425 59.605 ;
        RECT 180.565 59.745 180.885 59.805 ;
        RECT 185.625 59.745 185.945 59.805 ;
        RECT 192.985 59.745 193.305 59.805 ;
        RECT 180.565 59.605 185.945 59.745 ;
        RECT 180.565 59.545 180.885 59.605 ;
        RECT 185.625 59.545 185.945 59.605 ;
        RECT 186.635 59.605 188.615 59.745 ;
        RECT 175.965 59.205 176.285 59.465 ;
        RECT 172.285 59.065 172.605 59.125 ;
        RECT 173.680 59.065 173.970 59.110 ;
        RECT 172.285 58.925 173.970 59.065 ;
        RECT 172.285 58.865 172.605 58.925 ;
        RECT 173.680 58.880 173.970 58.925 ;
        RECT 172.760 58.725 173.050 58.770 ;
        RECT 176.055 58.725 176.195 59.205 ;
        RECT 181.025 59.065 181.345 59.125 ;
        RECT 178.815 58.925 181.345 59.065 ;
        RECT 172.760 58.585 176.195 58.725 ;
        RECT 176.900 58.725 177.190 58.770 ;
        RECT 177.345 58.725 177.665 58.785 ;
        RECT 176.900 58.585 177.665 58.725 ;
        RECT 172.760 58.540 173.050 58.585 ;
        RECT 176.900 58.540 177.190 58.585 ;
        RECT 177.345 58.525 177.665 58.585 ;
        RECT 173.220 58.385 173.510 58.430 ;
        RECT 178.815 58.385 178.955 58.925 ;
        RECT 181.025 58.865 181.345 58.925 ;
        RECT 183.340 59.065 183.630 59.110 ;
        RECT 183.785 59.065 184.105 59.125 ;
        RECT 183.340 58.925 184.105 59.065 ;
        RECT 183.340 58.880 183.630 58.925 ;
        RECT 183.785 58.865 184.105 58.925 ;
        RECT 184.720 59.065 185.010 59.110 ;
        RECT 186.635 59.065 186.775 59.605 ;
        RECT 188.475 59.405 188.615 59.605 ;
        RECT 192.985 59.605 194.135 59.745 ;
        RECT 192.985 59.545 193.305 59.605 ;
        RECT 189.305 59.405 189.625 59.465 ;
        RECT 188.475 59.265 189.625 59.405 ;
        RECT 189.305 59.205 189.625 59.265 ;
        RECT 189.765 59.065 190.085 59.125 ;
        RECT 184.720 58.925 186.775 59.065 ;
        RECT 188.475 58.925 190.085 59.065 ;
        RECT 184.720 58.880 185.010 58.925 ;
        RECT 179.200 58.540 179.490 58.770 ;
        RECT 180.120 58.725 180.410 58.770 ;
        RECT 182.405 58.725 182.725 58.785 ;
        RECT 180.120 58.585 182.725 58.725 ;
        RECT 180.120 58.540 180.410 58.585 ;
        RECT 173.220 58.245 178.955 58.385 ;
        RECT 179.275 58.385 179.415 58.540 ;
        RECT 180.565 58.385 180.885 58.445 ;
        RECT 179.275 58.245 180.885 58.385 ;
        RECT 173.220 58.200 173.510 58.245 ;
        RECT 180.565 58.185 180.885 58.245 ;
        RECT 167.685 58.045 168.005 58.105 ;
        RECT 170.920 58.045 171.210 58.090 ;
        RECT 167.685 57.905 171.210 58.045 ;
        RECT 167.685 57.845 168.005 57.905 ;
        RECT 170.920 57.860 171.210 57.905 ;
        RECT 177.805 58.045 178.125 58.105 ;
        RECT 181.115 58.045 181.255 58.585 ;
        RECT 182.405 58.525 182.725 58.585 ;
        RECT 182.880 58.540 183.170 58.770 ;
        RECT 182.955 58.385 183.095 58.540 ;
        RECT 185.625 58.525 185.945 58.785 ;
        RECT 186.085 58.525 186.405 58.785 ;
        RECT 186.545 58.735 186.865 58.785 ;
        RECT 188.475 58.770 188.615 58.925 ;
        RECT 189.765 58.865 190.085 58.925 ;
        RECT 190.685 59.065 191.005 59.125 ;
        RECT 193.995 59.110 194.135 59.605 ;
        RECT 197.585 59.545 197.905 59.805 ;
        RECT 211.845 59.745 212.165 59.805 ;
        RECT 220.585 59.745 220.905 59.805 ;
        RECT 211.845 59.605 218.515 59.745 ;
        RECT 211.845 59.545 212.165 59.605 ;
        RECT 201.265 59.405 201.585 59.465 ;
        RECT 202.660 59.405 202.950 59.450 ;
        RECT 201.265 59.265 202.950 59.405 ;
        RECT 201.265 59.205 201.585 59.265 ;
        RECT 202.660 59.220 202.950 59.265 ;
        RECT 214.605 59.205 214.925 59.465 ;
        RECT 218.375 59.450 218.515 59.605 ;
        RECT 220.215 59.605 220.905 59.745 ;
        RECT 218.300 59.220 218.590 59.450 ;
        RECT 218.760 59.405 219.050 59.450 ;
        RECT 220.215 59.405 220.355 59.605 ;
        RECT 220.585 59.545 220.905 59.605 ;
        RECT 222.425 59.745 222.745 59.805 ;
        RECT 224.280 59.745 224.570 59.790 ;
        RECT 244.505 59.745 244.825 59.805 ;
        RECT 246.345 59.745 246.665 59.805 ;
        RECT 247.740 59.745 248.030 59.790 ;
        RECT 262.905 59.745 263.225 59.805 ;
        RECT 222.425 59.605 224.570 59.745 ;
        RECT 222.425 59.545 222.745 59.605 ;
        RECT 224.280 59.560 224.570 59.605 ;
        RECT 243.215 59.605 263.225 59.745 ;
        RECT 233.430 59.405 233.720 59.450 ;
        RECT 235.320 59.405 235.610 59.450 ;
        RECT 238.440 59.405 238.730 59.450 ;
        RECT 218.760 59.265 220.355 59.405 ;
        RECT 220.675 59.265 227.255 59.405 ;
        RECT 218.760 59.220 219.050 59.265 ;
        RECT 191.160 59.065 191.450 59.110 ;
        RECT 190.685 58.925 191.450 59.065 ;
        RECT 190.685 58.865 191.005 58.925 ;
        RECT 191.160 58.880 191.450 58.925 ;
        RECT 192.155 58.925 193.675 59.065 ;
        RECT 192.155 58.785 192.295 58.925 ;
        RECT 187.020 58.735 187.310 58.770 ;
        RECT 186.545 58.595 187.310 58.735 ;
        RECT 186.545 58.525 186.865 58.595 ;
        RECT 187.020 58.540 187.310 58.595 ;
        RECT 188.400 58.540 188.690 58.770 ;
        RECT 191.620 58.725 191.910 58.770 ;
        RECT 188.935 58.585 191.910 58.725 ;
        RECT 185.165 58.385 185.485 58.445 ;
        RECT 188.935 58.385 189.075 58.585 ;
        RECT 191.620 58.540 191.910 58.585 ;
        RECT 192.065 58.525 192.385 58.785 ;
        RECT 192.985 58.525 193.305 58.785 ;
        RECT 193.535 58.725 193.675 58.925 ;
        RECT 193.920 58.880 194.210 59.110 ;
        RECT 201.725 59.065 202.045 59.125 ;
        RECT 203.120 59.065 203.410 59.110 ;
        RECT 201.725 58.925 203.410 59.065 ;
        RECT 201.725 58.865 202.045 58.925 ;
        RECT 203.120 58.880 203.410 58.925 ;
        RECT 215.065 58.865 215.385 59.125 ;
        RECT 220.675 59.065 220.815 59.265 ;
        RECT 216.075 58.925 220.815 59.065 ;
        RECT 221.045 59.065 221.365 59.125 ;
        RECT 227.115 59.110 227.255 59.265 ;
        RECT 233.430 59.265 238.730 59.405 ;
        RECT 233.430 59.220 233.720 59.265 ;
        RECT 235.320 59.220 235.610 59.265 ;
        RECT 238.440 59.220 238.730 59.265 ;
        RECT 241.285 59.205 241.605 59.465 ;
        RECT 223.360 59.065 223.650 59.110 ;
        RECT 221.045 58.925 226.335 59.065 ;
        RECT 195.760 58.725 196.050 58.770 ;
        RECT 193.535 58.585 196.050 58.725 ;
        RECT 195.760 58.540 196.050 58.585 ;
        RECT 196.205 58.725 196.525 58.785 ;
        RECT 196.680 58.725 196.970 58.770 ;
        RECT 196.205 58.585 196.970 58.725 ;
        RECT 196.205 58.525 196.525 58.585 ;
        RECT 196.680 58.540 196.970 58.585 ;
        RECT 198.965 58.725 199.285 58.785 ;
        RECT 200.345 58.725 200.665 58.785 ;
        RECT 202.200 58.725 202.490 58.770 ;
        RECT 198.965 58.585 202.490 58.725 ;
        RECT 198.965 58.525 199.285 58.585 ;
        RECT 200.345 58.525 200.665 58.585 ;
        RECT 202.200 58.540 202.490 58.585 ;
        RECT 203.580 58.725 203.870 58.770 ;
        RECT 204.485 58.725 204.805 58.785 ;
        RECT 203.580 58.585 204.805 58.725 ;
        RECT 203.580 58.540 203.870 58.585 ;
        RECT 182.955 58.245 189.075 58.385 ;
        RECT 202.275 58.385 202.415 58.540 ;
        RECT 204.485 58.525 204.805 58.585 ;
        RECT 212.305 58.525 212.625 58.785 ;
        RECT 214.145 58.525 214.465 58.785 ;
        RECT 214.605 58.725 214.925 58.785 ;
        RECT 215.540 58.725 215.830 58.770 ;
        RECT 214.605 58.585 215.830 58.725 ;
        RECT 214.605 58.525 214.925 58.585 ;
        RECT 215.540 58.540 215.830 58.585 ;
        RECT 208.625 58.385 208.945 58.445 ;
        RECT 212.395 58.385 212.535 58.525 ;
        RECT 202.275 58.245 212.535 58.385 ;
        RECT 213.685 58.385 214.005 58.445 ;
        RECT 216.075 58.385 216.215 58.925 ;
        RECT 221.045 58.865 221.365 58.925 ;
        RECT 223.360 58.880 223.650 58.925 ;
        RECT 216.460 58.540 216.750 58.770 ;
        RECT 216.905 58.725 217.225 58.785 ;
        RECT 217.840 58.725 218.130 58.770 ;
        RECT 216.905 58.585 218.130 58.725 ;
        RECT 213.685 58.245 216.215 58.385 ;
        RECT 216.535 58.385 216.675 58.540 ;
        RECT 216.905 58.525 217.225 58.585 ;
        RECT 217.840 58.540 218.130 58.585 ;
        RECT 219.220 58.725 219.510 58.770 ;
        RECT 221.980 58.725 222.270 58.770 ;
        RECT 223.805 58.725 224.125 58.785 ;
        RECT 219.220 58.585 221.275 58.725 ;
        RECT 219.220 58.540 219.510 58.585 ;
        RECT 218.285 58.385 218.605 58.445 ;
        RECT 220.585 58.385 220.905 58.445 ;
        RECT 216.535 58.245 220.905 58.385 ;
        RECT 185.165 58.185 185.485 58.245 ;
        RECT 208.625 58.185 208.945 58.245 ;
        RECT 213.685 58.185 214.005 58.245 ;
        RECT 218.285 58.185 218.605 58.245 ;
        RECT 220.585 58.185 220.905 58.245 ;
        RECT 177.805 57.905 181.255 58.045 ;
        RECT 183.325 58.045 183.645 58.105 ;
        RECT 191.145 58.045 191.465 58.105 ;
        RECT 183.325 57.905 191.465 58.045 ;
        RECT 177.805 57.845 178.125 57.905 ;
        RECT 183.325 57.845 183.645 57.905 ;
        RECT 191.145 57.845 191.465 57.905 ;
        RECT 198.045 58.045 198.365 58.105 ;
        RECT 201.280 58.045 201.570 58.090 ;
        RECT 198.045 57.905 201.570 58.045 ;
        RECT 198.045 57.845 198.365 57.905 ;
        RECT 201.280 57.860 201.570 57.905 ;
        RECT 212.305 58.045 212.625 58.105 ;
        RECT 213.240 58.045 213.530 58.090 ;
        RECT 212.305 57.905 213.530 58.045 ;
        RECT 212.305 57.845 212.625 57.905 ;
        RECT 213.240 57.860 213.530 57.905 ;
        RECT 215.065 58.045 215.385 58.105 ;
        RECT 216.920 58.045 217.210 58.090 ;
        RECT 215.065 57.905 217.210 58.045 ;
        RECT 215.065 57.845 215.385 57.905 ;
        RECT 216.920 57.860 217.210 57.905 ;
        RECT 217.365 58.045 217.685 58.105 ;
        RECT 220.140 58.045 220.430 58.090 ;
        RECT 217.365 57.905 220.430 58.045 ;
        RECT 221.135 58.045 221.275 58.585 ;
        RECT 221.980 58.585 224.125 58.725 ;
        RECT 221.980 58.540 222.270 58.585 ;
        RECT 223.805 58.525 224.125 58.585 ;
        RECT 222.440 58.385 222.730 58.430 ;
        RECT 222.885 58.385 223.205 58.445 ;
        RECT 222.440 58.245 223.205 58.385 ;
        RECT 222.440 58.200 222.730 58.245 ;
        RECT 222.885 58.185 223.205 58.245 ;
        RECT 225.200 58.385 225.490 58.430 ;
        RECT 225.645 58.385 225.965 58.445 ;
        RECT 226.195 58.430 226.335 58.925 ;
        RECT 227.040 58.880 227.330 59.110 ;
        RECT 227.485 59.065 227.805 59.125 ;
        RECT 243.215 59.110 243.355 59.605 ;
        RECT 244.505 59.545 244.825 59.605 ;
        RECT 246.345 59.545 246.665 59.605 ;
        RECT 247.740 59.560 248.030 59.605 ;
        RECT 262.905 59.545 263.225 59.605 ;
        RECT 279.005 59.745 279.325 59.805 ;
        RECT 304.765 59.745 305.085 59.805 ;
        RECT 279.005 59.605 305.085 59.745 ;
        RECT 279.005 59.545 279.325 59.605 ;
        RECT 244.980 59.405 245.270 59.450 ;
        RECT 245.885 59.405 246.205 59.465 ;
        RECT 244.980 59.265 246.205 59.405 ;
        RECT 244.980 59.220 245.270 59.265 ;
        RECT 245.885 59.205 246.205 59.265 ;
        RECT 251.880 59.405 252.170 59.450 ;
        RECT 252.785 59.405 253.105 59.465 ;
        RECT 251.880 59.265 253.105 59.405 ;
        RECT 251.880 59.220 252.170 59.265 ;
        RECT 252.785 59.205 253.105 59.265 ;
        RECT 253.670 59.405 253.960 59.450 ;
        RECT 255.560 59.405 255.850 59.450 ;
        RECT 258.680 59.405 258.970 59.450 ;
        RECT 253.670 59.265 258.970 59.405 ;
        RECT 253.670 59.220 253.960 59.265 ;
        RECT 255.560 59.220 255.850 59.265 ;
        RECT 258.680 59.220 258.970 59.265 ;
        RECT 284.490 59.405 284.780 59.450 ;
        RECT 286.380 59.405 286.670 59.450 ;
        RECT 289.500 59.405 289.790 59.450 ;
        RECT 284.490 59.265 289.790 59.405 ;
        RECT 284.490 59.220 284.780 59.265 ;
        RECT 286.380 59.220 286.670 59.265 ;
        RECT 289.500 59.220 289.790 59.265 ;
        RECT 292.345 59.205 292.665 59.465 ;
        RECT 294.735 59.450 294.875 59.605 ;
        RECT 304.765 59.545 305.085 59.605 ;
        RECT 294.660 59.220 294.950 59.450 ;
        RECT 297.520 59.405 297.810 59.450 ;
        RECT 300.640 59.405 300.930 59.450 ;
        RECT 302.530 59.405 302.820 59.450 ;
        RECT 297.520 59.265 302.820 59.405 ;
        RECT 297.520 59.220 297.810 59.265 ;
        RECT 300.640 59.220 300.930 59.265 ;
        RECT 302.530 59.220 302.820 59.265 ;
        RECT 244.045 59.110 244.365 59.125 ;
        RECT 227.485 58.925 242.435 59.065 ;
        RECT 227.485 58.865 227.805 58.925 ;
        RECT 228.405 58.725 228.725 58.785 ;
        RECT 232.545 58.725 232.865 58.785 ;
        RECT 228.405 58.585 232.865 58.725 ;
        RECT 228.405 58.525 228.725 58.585 ;
        RECT 232.545 58.525 232.865 58.585 ;
        RECT 233.025 58.725 233.315 58.770 ;
        RECT 234.860 58.725 235.150 58.770 ;
        RECT 238.440 58.725 238.730 58.770 ;
        RECT 233.025 58.585 238.730 58.725 ;
        RECT 233.025 58.540 233.315 58.585 ;
        RECT 234.860 58.540 235.150 58.585 ;
        RECT 238.440 58.540 238.730 58.585 ;
        RECT 225.200 58.245 225.965 58.385 ;
        RECT 225.200 58.200 225.490 58.245 ;
        RECT 225.645 58.185 225.965 58.245 ;
        RECT 226.120 58.385 226.410 58.430 ;
        RECT 232.085 58.385 232.405 58.445 ;
        RECT 226.120 58.245 232.405 58.385 ;
        RECT 226.120 58.200 226.410 58.245 ;
        RECT 232.085 58.185 232.405 58.245 ;
        RECT 233.925 58.185 234.245 58.445 ;
        RECT 236.685 58.430 237.005 58.445 ;
        RECT 236.220 58.385 237.005 58.430 ;
        RECT 239.520 58.430 239.810 58.745 ;
        RECT 241.760 58.540 242.050 58.770 ;
        RECT 242.295 58.725 242.435 58.925 ;
        RECT 243.140 58.880 243.430 59.110 ;
        RECT 244.045 58.880 244.475 59.110 ;
        RECT 249.120 59.065 249.410 59.110 ;
        RECT 249.565 59.065 249.885 59.125 ;
        RECT 256.465 59.065 256.785 59.125 ;
        RECT 261.540 59.065 261.830 59.110 ;
        RECT 249.120 58.925 249.885 59.065 ;
        RECT 249.120 58.880 249.410 58.925 ;
        RECT 244.045 58.865 244.365 58.880 ;
        RECT 249.565 58.865 249.885 58.925 ;
        RECT 250.115 58.925 261.830 59.065 ;
        RECT 250.115 58.770 250.255 58.925 ;
        RECT 256.465 58.865 256.785 58.925 ;
        RECT 261.540 58.880 261.830 58.925 ;
        RECT 263.825 59.065 264.145 59.125 ;
        RECT 268.900 59.065 269.190 59.110 ;
        RECT 263.825 58.925 269.190 59.065 ;
        RECT 263.825 58.865 264.145 58.925 ;
        RECT 268.900 58.880 269.190 58.925 ;
        RECT 269.345 59.065 269.665 59.125 ;
        RECT 279.480 59.065 279.770 59.110 ;
        RECT 279.925 59.065 280.245 59.125 ;
        RECT 269.345 58.925 271.875 59.065 ;
        RECT 269.345 58.865 269.665 58.925 ;
        RECT 246.820 58.725 247.110 58.770 ;
        RECT 242.295 58.585 247.110 58.725 ;
        RECT 246.820 58.540 247.110 58.585 ;
        RECT 250.040 58.540 250.330 58.770 ;
        RECT 239.520 58.385 240.110 58.430 ;
        RECT 236.220 58.245 240.110 58.385 ;
        RECT 241.835 58.385 241.975 58.540 ;
        RECT 252.785 58.525 253.105 58.785 ;
        RECT 253.265 58.725 253.555 58.770 ;
        RECT 255.100 58.725 255.390 58.770 ;
        RECT 258.680 58.725 258.970 58.770 ;
        RECT 253.265 58.585 258.970 58.725 ;
        RECT 253.265 58.540 253.555 58.585 ;
        RECT 255.100 58.540 255.390 58.585 ;
        RECT 258.680 58.540 258.970 58.585 ;
        RECT 248.185 58.385 248.505 58.445 ;
        RECT 241.835 58.245 248.505 58.385 ;
        RECT 236.220 58.200 237.005 58.245 ;
        RECT 239.820 58.200 240.110 58.245 ;
        RECT 236.685 58.185 237.005 58.200 ;
        RECT 248.185 58.185 248.505 58.245 ;
        RECT 253.705 58.385 254.025 58.445 ;
        RECT 254.180 58.385 254.470 58.430 ;
        RECT 253.705 58.245 254.470 58.385 ;
        RECT 253.705 58.185 254.025 58.245 ;
        RECT 254.180 58.200 254.470 58.245 ;
        RECT 256.460 58.385 257.110 58.430 ;
        RECT 259.225 58.385 259.545 58.445 ;
        RECT 259.760 58.430 260.050 58.745 ;
        RECT 269.805 58.725 270.125 58.785 ;
        RECT 271.735 58.770 271.875 58.925 ;
        RECT 279.480 58.925 280.245 59.065 ;
        RECT 279.480 58.880 279.770 58.925 ;
        RECT 279.925 58.865 280.245 58.925 ;
        RECT 284.985 58.865 285.305 59.125 ;
        RECT 299.245 59.065 299.565 59.125 ;
        RECT 296.115 58.925 299.565 59.065 ;
        RECT 271.200 58.725 271.490 58.770 ;
        RECT 269.805 58.585 271.490 58.725 ;
        RECT 269.805 58.525 270.125 58.585 ;
        RECT 271.200 58.540 271.490 58.585 ;
        RECT 271.660 58.540 271.950 58.770 ;
        RECT 283.605 58.525 283.925 58.785 ;
        RECT 284.085 58.725 284.375 58.770 ;
        RECT 285.920 58.725 286.210 58.770 ;
        RECT 289.500 58.725 289.790 58.770 ;
        RECT 284.085 58.585 289.790 58.725 ;
        RECT 284.085 58.540 284.375 58.585 ;
        RECT 285.920 58.540 286.210 58.585 ;
        RECT 289.500 58.540 289.790 58.585 ;
        RECT 259.760 58.385 260.350 58.430 ;
        RECT 256.460 58.245 260.350 58.385 ;
        RECT 256.460 58.200 257.110 58.245 ;
        RECT 259.225 58.185 259.545 58.245 ;
        RECT 260.060 58.200 260.350 58.245 ;
        RECT 269.360 58.385 269.650 58.430 ;
        RECT 272.105 58.385 272.425 58.445 ;
        RECT 269.360 58.245 272.425 58.385 ;
        RECT 269.360 58.200 269.650 58.245 ;
        RECT 272.105 58.185 272.425 58.245 ;
        RECT 274.865 58.385 275.185 58.445 ;
        RECT 280.400 58.385 280.690 58.430 ;
        RECT 285.445 58.385 285.765 58.445 ;
        RECT 274.865 58.245 280.690 58.385 ;
        RECT 274.865 58.185 275.185 58.245 ;
        RECT 280.400 58.200 280.690 58.245 ;
        RECT 281.855 58.245 285.765 58.385 ;
        RECT 229.785 58.045 230.105 58.105 ;
        RECT 221.135 57.905 230.105 58.045 ;
        RECT 217.365 57.845 217.685 57.905 ;
        RECT 220.140 57.860 220.430 57.905 ;
        RECT 229.785 57.845 230.105 57.905 ;
        RECT 230.260 58.045 230.550 58.090 ;
        RECT 237.145 58.045 237.465 58.105 ;
        RECT 230.260 57.905 237.465 58.045 ;
        RECT 230.260 57.860 230.550 57.905 ;
        RECT 237.145 57.845 237.465 57.905 ;
        RECT 243.600 58.045 243.890 58.090 ;
        RECT 246.345 58.045 246.665 58.105 ;
        RECT 243.600 57.905 246.665 58.045 ;
        RECT 243.600 57.860 243.890 57.905 ;
        RECT 246.345 57.845 246.665 57.905 ;
        RECT 249.565 57.845 249.885 58.105 ;
        RECT 254.625 58.045 254.945 58.105 ;
        RECT 263.825 58.045 264.145 58.105 ;
        RECT 254.625 57.905 264.145 58.045 ;
        RECT 254.625 57.845 254.945 57.905 ;
        RECT 263.825 57.845 264.145 57.905 ;
        RECT 279.005 58.045 279.325 58.105 ;
        RECT 279.940 58.045 280.230 58.090 ;
        RECT 281.855 58.045 281.995 58.245 ;
        RECT 285.445 58.185 285.765 58.245 ;
        RECT 286.365 58.385 286.685 58.445 ;
        RECT 287.285 58.430 287.605 58.445 ;
        RECT 290.580 58.430 290.870 58.745 ;
        RECT 296.115 58.430 296.255 58.925 ;
        RECT 299.245 58.865 299.565 58.925 ;
        RECT 299.705 59.065 300.025 59.125 ;
        RECT 303.400 59.065 303.690 59.110 ;
        RECT 299.705 58.925 303.690 59.065 ;
        RECT 299.705 58.865 300.025 58.925 ;
        RECT 303.400 58.880 303.690 58.925 ;
        RECT 296.440 58.430 296.730 58.745 ;
        RECT 297.520 58.725 297.810 58.770 ;
        RECT 301.100 58.725 301.390 58.770 ;
        RECT 302.935 58.725 303.225 58.770 ;
        RECT 297.520 58.585 303.225 58.725 ;
        RECT 297.520 58.540 297.810 58.585 ;
        RECT 301.100 58.540 301.390 58.585 ;
        RECT 302.935 58.540 303.225 58.585 ;
        RECT 287.280 58.385 287.930 58.430 ;
        RECT 290.580 58.385 291.170 58.430 ;
        RECT 296.115 58.385 296.730 58.430 ;
        RECT 299.380 58.385 300.030 58.430 ;
        RECT 286.365 58.245 291.170 58.385 ;
        RECT 286.365 58.185 286.685 58.245 ;
        RECT 279.005 57.905 281.995 58.045 ;
        RECT 279.005 57.845 279.325 57.905 ;
        RECT 279.940 57.860 280.230 57.905 ;
        RECT 282.225 57.845 282.545 58.105 ;
        RECT 286.915 58.045 287.055 58.245 ;
        RECT 287.280 58.200 287.930 58.245 ;
        RECT 290.880 58.200 291.170 58.245 ;
        RECT 291.515 58.245 300.030 58.385 ;
        RECT 287.285 58.185 287.605 58.200 ;
        RECT 291.515 58.045 291.655 58.245 ;
        RECT 296.140 58.200 296.430 58.245 ;
        RECT 299.380 58.200 300.030 58.245 ;
        RECT 302.005 58.185 302.325 58.445 ;
        RECT 286.915 57.905 291.655 58.045 ;
        RECT 162.095 57.225 311.135 57.705 ;
        RECT 176.885 57.025 177.205 57.085 ;
        RECT 177.360 57.025 177.650 57.070 ;
        RECT 179.645 57.025 179.965 57.085 ;
        RECT 176.885 56.885 179.965 57.025 ;
        RECT 176.885 56.825 177.205 56.885 ;
        RECT 177.360 56.840 177.650 56.885 ;
        RECT 179.645 56.825 179.965 56.885 ;
        RECT 182.865 56.825 183.185 57.085 ;
        RECT 185.165 56.825 185.485 57.085 ;
        RECT 186.545 57.025 186.865 57.085 ;
        RECT 188.400 57.025 188.690 57.070 ;
        RECT 193.920 57.025 194.210 57.070 ;
        RECT 186.545 56.885 188.690 57.025 ;
        RECT 186.545 56.825 186.865 56.885 ;
        RECT 188.400 56.840 188.690 56.885 ;
        RECT 189.855 56.885 194.210 57.025 ;
        RECT 167.685 56.485 168.005 56.745 ;
        RECT 169.980 56.685 170.630 56.730 ;
        RECT 173.580 56.685 173.870 56.730 ;
        RECT 174.125 56.685 174.445 56.745 ;
        RECT 169.980 56.545 174.445 56.685 ;
        RECT 169.980 56.500 170.630 56.545 ;
        RECT 173.280 56.500 173.870 56.545 ;
        RECT 166.785 56.345 167.075 56.390 ;
        RECT 168.620 56.345 168.910 56.390 ;
        RECT 172.200 56.345 172.490 56.390 ;
        RECT 166.785 56.205 172.490 56.345 ;
        RECT 166.785 56.160 167.075 56.205 ;
        RECT 168.620 56.160 168.910 56.205 ;
        RECT 172.200 56.160 172.490 56.205 ;
        RECT 173.280 56.185 173.570 56.500 ;
        RECT 174.125 56.485 174.445 56.545 ;
        RECT 177.805 56.485 178.125 56.745 ;
        RECT 180.120 56.685 180.410 56.730 ;
        RECT 181.485 56.685 181.805 56.745 ;
        RECT 182.955 56.685 183.095 56.825 ;
        RECT 180.120 56.545 183.095 56.685 ;
        RECT 180.120 56.500 180.410 56.545 ;
        RECT 181.485 56.485 181.805 56.545 ;
        RECT 175.045 56.345 175.365 56.405 ;
        RECT 180.565 56.345 180.885 56.405 ;
        RECT 181.040 56.345 181.330 56.390 ;
        RECT 183.340 56.345 183.630 56.390 ;
        RECT 185.255 56.345 185.395 56.825 ;
        RECT 189.305 56.685 189.625 56.745 ;
        RECT 189.855 56.730 189.995 56.885 ;
        RECT 193.920 56.840 194.210 56.885 ;
        RECT 194.840 57.025 195.130 57.070 ;
        RECT 195.745 57.025 196.065 57.085 ;
        RECT 194.840 56.885 196.065 57.025 ;
        RECT 194.840 56.840 195.130 56.885 ;
        RECT 195.745 56.825 196.065 56.885 ;
        RECT 204.025 57.025 204.345 57.085 ;
        RECT 204.500 57.025 204.790 57.070 ;
        RECT 204.025 56.885 204.790 57.025 ;
        RECT 204.025 56.825 204.345 56.885 ;
        RECT 204.500 56.840 204.790 56.885 ;
        RECT 204.945 57.025 205.265 57.085 ;
        RECT 249.565 57.025 249.885 57.085 ;
        RECT 204.945 56.885 249.885 57.025 ;
        RECT 204.945 56.825 205.265 56.885 ;
        RECT 249.565 56.825 249.885 56.885 ;
        RECT 250.025 57.025 250.345 57.085 ;
        RECT 259.685 57.025 260.005 57.085 ;
        RECT 260.160 57.025 260.450 57.070 ;
        RECT 250.025 56.885 259.455 57.025 ;
        RECT 250.025 56.825 250.345 56.885 ;
        RECT 189.780 56.685 190.070 56.730 ;
        RECT 193.460 56.685 193.750 56.730 ;
        RECT 175.045 56.205 180.335 56.345 ;
        RECT 175.045 56.145 175.365 56.205 ;
        RECT 166.305 55.805 166.625 56.065 ;
        RECT 178.740 56.005 179.030 56.050 ;
        RECT 179.645 56.005 179.965 56.065 ;
        RECT 178.740 55.865 179.965 56.005 ;
        RECT 180.195 56.005 180.335 56.205 ;
        RECT 180.565 56.205 183.095 56.345 ;
        RECT 180.565 56.145 180.885 56.205 ;
        RECT 181.040 56.160 181.330 56.205 ;
        RECT 181.960 56.005 182.250 56.050 ;
        RECT 182.405 56.005 182.725 56.065 ;
        RECT 180.195 55.865 182.725 56.005 ;
        RECT 182.955 56.005 183.095 56.205 ;
        RECT 183.340 56.205 185.395 56.345 ;
        RECT 185.715 56.545 190.070 56.685 ;
        RECT 185.715 56.345 185.855 56.545 ;
        RECT 189.305 56.485 189.625 56.545 ;
        RECT 189.780 56.500 190.070 56.545 ;
        RECT 192.155 56.545 193.750 56.685 ;
        RECT 192.155 56.405 192.295 56.545 ;
        RECT 193.460 56.500 193.750 56.545 ;
        RECT 196.665 56.485 196.985 56.745 ;
        RECT 197.125 56.685 197.445 56.745 ;
        RECT 198.960 56.685 199.610 56.730 ;
        RECT 202.560 56.685 202.850 56.730 ;
        RECT 197.125 56.545 202.850 56.685 ;
        RECT 197.125 56.485 197.445 56.545 ;
        RECT 198.960 56.500 199.610 56.545 ;
        RECT 202.260 56.500 202.850 56.545 ;
        RECT 213.240 56.685 213.530 56.730 ;
        RECT 215.985 56.685 216.305 56.745 ;
        RECT 220.125 56.685 220.445 56.745 ;
        RECT 213.240 56.545 216.305 56.685 ;
        RECT 213.240 56.500 213.530 56.545 ;
        RECT 187.005 56.390 187.325 56.405 ;
        RECT 186.400 56.345 186.690 56.390 ;
        RECT 185.715 56.205 186.690 56.345 ;
        RECT 183.340 56.160 183.630 56.205 ;
        RECT 186.400 56.160 186.690 56.205 ;
        RECT 186.895 56.160 187.325 56.390 ;
        RECT 190.240 56.345 190.530 56.390 ;
        RECT 192.065 56.345 192.385 56.405 ;
        RECT 190.240 56.205 192.385 56.345 ;
        RECT 190.240 56.160 190.530 56.205 ;
        RECT 187.005 56.145 187.325 56.160 ;
        RECT 192.065 56.145 192.385 56.205 ;
        RECT 193.000 56.160 193.290 56.390 ;
        RECT 195.765 56.345 196.055 56.390 ;
        RECT 197.600 56.345 197.890 56.390 ;
        RECT 201.180 56.345 201.470 56.390 ;
        RECT 195.765 56.205 201.470 56.345 ;
        RECT 195.765 56.160 196.055 56.205 ;
        RECT 197.600 56.160 197.890 56.205 ;
        RECT 201.180 56.160 201.470 56.205 ;
        RECT 202.260 56.185 202.550 56.500 ;
        RECT 215.985 56.485 216.305 56.545 ;
        RECT 219.295 56.545 220.445 56.685 ;
        RECT 205.420 56.160 205.710 56.390 ;
        RECT 206.340 56.345 206.630 56.390 ;
        RECT 208.625 56.345 208.945 56.405 ;
        RECT 211.400 56.345 211.690 56.390 ;
        RECT 206.340 56.205 211.690 56.345 ;
        RECT 206.340 56.160 206.630 56.205 ;
        RECT 184.705 56.005 185.025 56.065 ;
        RECT 185.625 56.005 185.945 56.065 ;
        RECT 189.195 56.005 189.485 56.050 ;
        RECT 182.955 55.865 184.475 56.005 ;
        RECT 178.740 55.820 179.030 55.865 ;
        RECT 179.645 55.805 179.965 55.865 ;
        RECT 181.960 55.820 182.250 55.865 ;
        RECT 182.405 55.805 182.725 55.865 ;
        RECT 167.190 55.665 167.480 55.710 ;
        RECT 169.080 55.665 169.370 55.710 ;
        RECT 172.200 55.665 172.490 55.710 ;
        RECT 167.190 55.525 172.490 55.665 ;
        RECT 167.190 55.480 167.480 55.525 ;
        RECT 169.080 55.480 169.370 55.525 ;
        RECT 172.200 55.480 172.490 55.525 ;
        RECT 175.060 55.665 175.350 55.710 ;
        RECT 177.345 55.665 177.665 55.725 ;
        RECT 183.325 55.665 183.645 55.725 ;
        RECT 175.060 55.525 183.645 55.665 ;
        RECT 175.060 55.480 175.350 55.525 ;
        RECT 177.345 55.465 177.665 55.525 ;
        RECT 183.325 55.465 183.645 55.525 ;
        RECT 183.785 55.465 184.105 55.725 ;
        RECT 184.335 55.665 184.475 55.865 ;
        RECT 184.705 55.865 189.485 56.005 ;
        RECT 184.705 55.805 185.025 55.865 ;
        RECT 185.625 55.805 185.945 55.865 ;
        RECT 189.195 55.820 189.485 55.865 ;
        RECT 191.605 56.005 191.925 56.065 ;
        RECT 193.075 56.005 193.215 56.160 ;
        RECT 191.605 55.865 193.215 56.005 ;
        RECT 186.545 55.665 186.865 55.725 ;
        RECT 184.335 55.525 186.865 55.665 ;
        RECT 189.270 55.665 189.410 55.820 ;
        RECT 191.605 55.805 191.925 55.865 ;
        RECT 195.300 55.820 195.590 56.050 ;
        RECT 204.040 56.005 204.330 56.050 ;
        RECT 205.495 56.005 205.635 56.160 ;
        RECT 208.625 56.145 208.945 56.205 ;
        RECT 211.400 56.160 211.690 56.205 ;
        RECT 212.320 56.345 212.610 56.390 ;
        RECT 215.525 56.345 215.845 56.405 ;
        RECT 212.320 56.205 215.845 56.345 ;
        RECT 212.320 56.160 212.610 56.205 ;
        RECT 210.925 56.005 211.245 56.065 ;
        RECT 204.040 55.865 211.245 56.005 ;
        RECT 211.475 56.005 211.615 56.160 ;
        RECT 215.525 56.145 215.845 56.205 ;
        RECT 218.745 56.145 219.065 56.405 ;
        RECT 219.295 56.390 219.435 56.545 ;
        RECT 220.125 56.485 220.445 56.545 ;
        RECT 220.585 56.485 220.905 56.745 ;
        RECT 222.880 56.685 223.530 56.730 ;
        RECT 226.480 56.685 226.770 56.730 ;
        RECT 229.800 56.685 230.090 56.730 ;
        RECT 230.245 56.685 230.565 56.745 ;
        RECT 222.880 56.545 228.175 56.685 ;
        RECT 222.880 56.500 223.530 56.545 ;
        RECT 226.180 56.500 226.770 56.545 ;
        RECT 219.220 56.160 219.510 56.390 ;
        RECT 219.685 56.345 219.975 56.390 ;
        RECT 221.520 56.345 221.810 56.390 ;
        RECT 225.100 56.345 225.390 56.390 ;
        RECT 219.685 56.205 225.390 56.345 ;
        RECT 219.685 56.160 219.975 56.205 ;
        RECT 221.520 56.160 221.810 56.205 ;
        RECT 225.100 56.160 225.390 56.205 ;
        RECT 226.180 56.185 226.470 56.500 ;
        RECT 218.285 56.005 218.605 56.065 ;
        RECT 227.485 56.005 227.805 56.065 ;
        RECT 211.475 55.865 218.605 56.005 ;
        RECT 204.040 55.820 204.330 55.865 ;
        RECT 192.080 55.665 192.370 55.710 ;
        RECT 192.985 55.665 193.305 55.725 ;
        RECT 189.270 55.525 193.305 55.665 ;
        RECT 186.545 55.465 186.865 55.525 ;
        RECT 192.080 55.480 192.370 55.525 ;
        RECT 192.985 55.465 193.305 55.525 ;
        RECT 193.445 55.665 193.765 55.725 ;
        RECT 195.375 55.665 195.515 55.820 ;
        RECT 210.925 55.805 211.245 55.865 ;
        RECT 218.285 55.805 218.605 55.865 ;
        RECT 219.755 55.865 227.805 56.005 ;
        RECT 193.445 55.525 195.515 55.665 ;
        RECT 196.170 55.665 196.460 55.710 ;
        RECT 198.060 55.665 198.350 55.710 ;
        RECT 201.180 55.665 201.470 55.710 ;
        RECT 219.755 55.665 219.895 55.865 ;
        RECT 227.485 55.805 227.805 55.865 ;
        RECT 228.035 56.005 228.175 56.545 ;
        RECT 229.800 56.545 230.565 56.685 ;
        RECT 229.800 56.500 230.090 56.545 ;
        RECT 230.245 56.485 230.565 56.545 ;
        RECT 232.080 56.685 232.730 56.730 ;
        RECT 235.680 56.685 235.970 56.730 ;
        RECT 236.685 56.685 237.005 56.745 ;
        RECT 232.080 56.545 237.005 56.685 ;
        RECT 232.080 56.500 232.730 56.545 ;
        RECT 235.380 56.500 235.995 56.545 ;
        RECT 228.405 56.145 228.725 56.405 ;
        RECT 228.885 56.345 229.175 56.390 ;
        RECT 230.720 56.345 231.010 56.390 ;
        RECT 234.300 56.345 234.590 56.390 ;
        RECT 228.885 56.205 234.590 56.345 ;
        RECT 228.885 56.160 229.175 56.205 ;
        RECT 230.720 56.160 231.010 56.205 ;
        RECT 234.300 56.160 234.590 56.205 ;
        RECT 235.380 56.185 235.670 56.500 ;
        RECT 235.855 56.005 235.995 56.500 ;
        RECT 236.685 56.485 237.005 56.545 ;
        RECT 243.125 56.485 243.445 56.745 ;
        RECT 244.060 56.685 244.350 56.730 ;
        RECT 251.405 56.685 251.725 56.745 ;
        RECT 252.800 56.685 253.090 56.730 ;
        RECT 244.060 56.545 246.575 56.685 ;
        RECT 244.060 56.500 244.350 56.545 ;
        RECT 239.445 56.345 239.765 56.405 ;
        RECT 240.840 56.345 241.130 56.390 ;
        RECT 239.445 56.205 241.130 56.345 ;
        RECT 239.445 56.145 239.765 56.205 ;
        RECT 240.840 56.160 241.130 56.205 ;
        RECT 241.760 56.345 242.050 56.390 ;
        RECT 241.760 56.205 242.895 56.345 ;
        RECT 241.760 56.160 242.050 56.205 ;
        RECT 228.035 55.865 235.995 56.005 ;
        RECT 242.755 56.005 242.895 56.205 ;
        RECT 244.135 56.005 244.275 56.500 ;
        RECT 246.435 56.390 246.575 56.545 ;
        RECT 251.405 56.545 253.090 56.685 ;
        RECT 251.405 56.485 251.725 56.545 ;
        RECT 252.800 56.500 253.090 56.545 ;
        RECT 255.080 56.685 255.730 56.730 ;
        RECT 256.005 56.685 256.325 56.745 ;
        RECT 258.680 56.685 258.970 56.730 ;
        RECT 255.080 56.545 258.970 56.685 ;
        RECT 259.315 56.685 259.455 56.885 ;
        RECT 259.685 56.885 260.450 57.025 ;
        RECT 259.685 56.825 260.005 56.885 ;
        RECT 260.160 56.840 260.450 56.885 ;
        RECT 270.265 57.025 270.585 57.085 ;
        RECT 274.865 57.025 275.185 57.085 ;
        RECT 270.265 56.885 275.185 57.025 ;
        RECT 270.265 56.825 270.585 56.885 ;
        RECT 274.865 56.825 275.185 56.885 ;
        RECT 299.245 57.025 299.565 57.085 ;
        RECT 299.245 56.885 303.155 57.025 ;
        RECT 299.245 56.825 299.565 56.885 ;
        RECT 264.285 56.685 264.605 56.745 ;
        RECT 265.680 56.685 265.970 56.730 ;
        RECT 259.315 56.545 265.970 56.685 ;
        RECT 255.080 56.500 255.730 56.545 ;
        RECT 256.005 56.485 256.325 56.545 ;
        RECT 258.380 56.500 258.970 56.545 ;
        RECT 245.445 56.160 245.735 56.390 ;
        RECT 246.360 56.345 246.650 56.390 ;
        RECT 251.885 56.345 252.175 56.390 ;
        RECT 253.720 56.345 254.010 56.390 ;
        RECT 257.300 56.345 257.590 56.390 ;
        RECT 246.360 56.205 247.495 56.345 ;
        RECT 246.360 56.160 246.650 56.205 ;
        RECT 242.755 55.865 244.275 56.005 ;
        RECT 245.515 56.005 245.655 56.160 ;
        RECT 245.885 56.005 246.205 56.065 ;
        RECT 245.515 55.865 246.205 56.005 ;
        RECT 196.170 55.525 201.470 55.665 ;
        RECT 193.445 55.465 193.765 55.525 ;
        RECT 196.170 55.480 196.460 55.525 ;
        RECT 198.060 55.480 198.350 55.525 ;
        RECT 201.180 55.480 201.470 55.525 ;
        RECT 201.815 55.525 219.895 55.665 ;
        RECT 220.090 55.665 220.380 55.710 ;
        RECT 221.980 55.665 222.270 55.710 ;
        RECT 225.100 55.665 225.390 55.710 ;
        RECT 220.090 55.525 225.390 55.665 ;
        RECT 175.505 55.125 175.825 55.385 ;
        RECT 184.260 55.325 184.550 55.370 ;
        RECT 188.385 55.325 188.705 55.385 ;
        RECT 184.260 55.185 188.705 55.325 ;
        RECT 184.260 55.140 184.550 55.185 ;
        RECT 188.385 55.125 188.705 55.185 ;
        RECT 189.765 55.325 190.085 55.385 ;
        RECT 193.905 55.325 194.225 55.385 ;
        RECT 189.765 55.185 194.225 55.325 ;
        RECT 189.765 55.125 190.085 55.185 ;
        RECT 193.905 55.125 194.225 55.185 ;
        RECT 194.365 55.325 194.685 55.385 ;
        RECT 201.815 55.325 201.955 55.525 ;
        RECT 220.090 55.480 220.380 55.525 ;
        RECT 221.980 55.480 222.270 55.525 ;
        RECT 225.100 55.480 225.390 55.525 ;
        RECT 226.105 55.665 226.425 55.725 ;
        RECT 228.035 55.665 228.175 55.865 ;
        RECT 245.885 55.805 246.205 55.865 ;
        RECT 226.105 55.525 228.175 55.665 ;
        RECT 229.290 55.665 229.580 55.710 ;
        RECT 231.180 55.665 231.470 55.710 ;
        RECT 234.300 55.665 234.590 55.710 ;
        RECT 229.290 55.525 234.590 55.665 ;
        RECT 226.105 55.465 226.425 55.525 ;
        RECT 229.290 55.480 229.580 55.525 ;
        RECT 231.180 55.480 231.470 55.525 ;
        RECT 234.300 55.480 234.590 55.525 ;
        RECT 234.845 55.665 235.165 55.725 ;
        RECT 237.160 55.665 237.450 55.710 ;
        RECT 244.520 55.665 244.810 55.710 ;
        RECT 234.845 55.525 237.450 55.665 ;
        RECT 234.845 55.465 235.165 55.525 ;
        RECT 237.160 55.480 237.450 55.525 ;
        RECT 237.695 55.525 244.810 55.665 ;
        RECT 194.365 55.185 201.955 55.325 ;
        RECT 214.605 55.325 214.925 55.385 ;
        RECT 215.540 55.325 215.830 55.370 ;
        RECT 214.605 55.185 215.830 55.325 ;
        RECT 194.365 55.125 194.685 55.185 ;
        RECT 214.605 55.125 214.925 55.185 ;
        RECT 215.540 55.140 215.830 55.185 ;
        RECT 218.745 55.325 219.065 55.385 ;
        RECT 219.665 55.325 219.985 55.385 ;
        RECT 224.265 55.325 224.585 55.385 ;
        RECT 218.745 55.185 224.585 55.325 ;
        RECT 218.745 55.125 219.065 55.185 ;
        RECT 219.665 55.125 219.985 55.185 ;
        RECT 224.265 55.125 224.585 55.185 ;
        RECT 225.645 55.325 225.965 55.385 ;
        RECT 227.960 55.325 228.250 55.370 ;
        RECT 231.625 55.325 231.945 55.385 ;
        RECT 225.645 55.185 231.945 55.325 ;
        RECT 225.645 55.125 225.965 55.185 ;
        RECT 227.960 55.140 228.250 55.185 ;
        RECT 231.625 55.125 231.945 55.185 ;
        RECT 233.005 55.325 233.325 55.385 ;
        RECT 237.695 55.325 237.835 55.525 ;
        RECT 244.520 55.480 244.810 55.525 ;
        RECT 233.005 55.185 237.835 55.325 ;
        RECT 238.985 55.325 239.305 55.385 ;
        RECT 239.920 55.325 240.210 55.370 ;
        RECT 238.985 55.185 240.210 55.325 ;
        RECT 233.005 55.125 233.325 55.185 ;
        RECT 238.985 55.125 239.305 55.185 ;
        RECT 239.920 55.140 240.210 55.185 ;
        RECT 242.220 55.325 242.510 55.370 ;
        RECT 243.125 55.325 243.445 55.385 ;
        RECT 242.220 55.185 243.445 55.325 ;
        RECT 247.355 55.325 247.495 56.205 ;
        RECT 251.885 56.205 257.590 56.345 ;
        RECT 251.885 56.160 252.175 56.205 ;
        RECT 253.720 56.160 254.010 56.205 ;
        RECT 257.300 56.160 257.590 56.205 ;
        RECT 258.380 56.185 258.670 56.500 ;
        RECT 264.285 56.485 264.605 56.545 ;
        RECT 265.680 56.500 265.970 56.545 ;
        RECT 276.360 56.685 276.650 56.730 ;
        RECT 279.600 56.685 280.250 56.730 ;
        RECT 276.360 56.545 280.250 56.685 ;
        RECT 276.360 56.500 276.950 56.545 ;
        RECT 279.600 56.500 280.250 56.545 ;
        RECT 276.660 56.405 276.950 56.500 ;
        RECT 282.225 56.485 282.545 56.745 ;
        RECT 283.605 56.685 283.925 56.745 ;
        RECT 289.585 56.685 289.905 56.745 ;
        RECT 295.120 56.685 295.410 56.730 ;
        RECT 283.605 56.545 295.410 56.685 ;
        RECT 283.605 56.485 283.925 56.545 ;
        RECT 289.585 56.485 289.905 56.545 ;
        RECT 295.120 56.500 295.410 56.545 ;
        RECT 300.645 56.685 300.935 56.730 ;
        RECT 302.505 56.685 302.795 56.730 ;
        RECT 300.645 56.545 302.795 56.685 ;
        RECT 303.015 56.685 303.155 56.885 ;
        RECT 303.425 56.685 303.715 56.730 ;
        RECT 306.685 56.685 306.975 56.730 ;
        RECT 303.015 56.545 306.975 56.685 ;
        RECT 300.645 56.500 300.935 56.545 ;
        RECT 302.505 56.500 302.795 56.545 ;
        RECT 303.425 56.500 303.715 56.545 ;
        RECT 306.685 56.500 306.975 56.545 ;
        RECT 262.905 56.145 263.225 56.405 ;
        RECT 276.660 56.185 277.025 56.405 ;
        RECT 276.705 56.145 277.025 56.185 ;
        RECT 277.740 56.345 278.030 56.390 ;
        RECT 281.320 56.345 281.610 56.390 ;
        RECT 283.155 56.345 283.445 56.390 ;
        RECT 277.740 56.205 283.445 56.345 ;
        RECT 277.740 56.160 278.030 56.205 ;
        RECT 281.320 56.160 281.610 56.205 ;
        RECT 283.155 56.160 283.445 56.205 ;
        RECT 290.060 56.345 290.350 56.390 ;
        RECT 291.440 56.345 291.730 56.390 ;
        RECT 290.060 56.205 291.730 56.345 ;
        RECT 295.195 56.345 295.335 56.500 ;
        RECT 299.705 56.345 300.025 56.405 ;
        RECT 295.195 56.205 300.025 56.345 ;
        RECT 302.580 56.345 302.795 56.500 ;
        RECT 304.825 56.345 305.115 56.390 ;
        RECT 302.580 56.205 305.115 56.345 ;
        RECT 290.060 56.160 290.350 56.205 ;
        RECT 291.440 56.160 291.730 56.205 ;
        RECT 251.420 56.005 251.710 56.050 ;
        RECT 252.785 56.005 253.105 56.065 ;
        RECT 254.625 56.005 254.945 56.065 ;
        RECT 251.420 55.865 254.945 56.005 ;
        RECT 251.420 55.820 251.710 55.865 ;
        RECT 252.785 55.805 253.105 55.865 ;
        RECT 254.625 55.805 254.945 55.865 ;
        RECT 261.065 56.005 261.385 56.065 ;
        RECT 268.440 56.005 268.730 56.050 ;
        RECT 261.065 55.865 268.730 56.005 ;
        RECT 261.065 55.805 261.385 55.865 ;
        RECT 268.440 55.820 268.730 55.865 ;
        RECT 283.605 55.805 283.925 56.065 ;
        RECT 286.380 56.005 286.670 56.050 ;
        RECT 287.285 56.005 287.605 56.065 ;
        RECT 286.380 55.865 287.605 56.005 ;
        RECT 286.380 55.820 286.670 55.865 ;
        RECT 287.285 55.805 287.605 55.865 ;
        RECT 252.290 55.665 252.580 55.710 ;
        RECT 254.180 55.665 254.470 55.710 ;
        RECT 257.300 55.665 257.590 55.710 ;
        RECT 277.740 55.665 278.030 55.710 ;
        RECT 280.860 55.665 281.150 55.710 ;
        RECT 282.750 55.665 283.040 55.710 ;
        RECT 252.290 55.525 257.590 55.665 ;
        RECT 252.290 55.480 252.580 55.525 ;
        RECT 254.180 55.480 254.470 55.525 ;
        RECT 257.300 55.480 257.590 55.525 ;
        RECT 269.665 55.525 277.395 55.665 ;
        RECT 253.245 55.325 253.565 55.385 ;
        RECT 247.355 55.185 253.565 55.325 ;
        RECT 242.220 55.140 242.510 55.185 ;
        RECT 243.125 55.125 243.445 55.185 ;
        RECT 253.245 55.125 253.565 55.185 ;
        RECT 256.005 55.325 256.325 55.385 ;
        RECT 269.665 55.325 269.805 55.525 ;
        RECT 256.005 55.185 269.805 55.325 ;
        RECT 277.255 55.325 277.395 55.525 ;
        RECT 277.740 55.525 283.040 55.665 ;
        RECT 277.740 55.480 278.030 55.525 ;
        RECT 280.860 55.480 281.150 55.525 ;
        RECT 282.750 55.480 283.040 55.525 ;
        RECT 285.905 55.325 286.225 55.385 ;
        RECT 290.135 55.325 290.275 56.160 ;
        RECT 299.705 56.145 300.025 56.205 ;
        RECT 304.825 56.160 305.115 56.205 ;
        RECT 301.560 56.005 301.850 56.050 ;
        RECT 308.445 56.005 308.765 56.065 ;
        RECT 301.560 55.865 308.765 56.005 ;
        RECT 301.560 55.820 301.850 55.865 ;
        RECT 308.445 55.805 308.765 55.865 ;
        RECT 300.185 55.665 300.475 55.710 ;
        RECT 302.045 55.665 302.335 55.710 ;
        RECT 304.825 55.665 305.115 55.710 ;
        RECT 300.185 55.525 305.115 55.665 ;
        RECT 300.185 55.480 300.475 55.525 ;
        RECT 302.045 55.480 302.335 55.525 ;
        RECT 304.825 55.480 305.115 55.525 ;
        RECT 308.905 55.370 309.225 55.385 ;
        RECT 277.255 55.185 290.275 55.325 ;
        RECT 256.005 55.125 256.325 55.185 ;
        RECT 285.905 55.125 286.225 55.185 ;
        RECT 308.690 55.140 309.225 55.370 ;
        RECT 308.905 55.125 309.225 55.140 ;
        RECT 162.095 54.505 311.135 54.985 ;
        RECT 187.020 54.305 187.310 54.350 ;
        RECT 188.845 54.305 189.165 54.365 ;
        RECT 187.020 54.165 189.165 54.305 ;
        RECT 187.020 54.120 187.310 54.165 ;
        RECT 188.845 54.105 189.165 54.165 ;
        RECT 189.320 54.305 189.610 54.350 ;
        RECT 189.765 54.305 190.085 54.365 ;
        RECT 189.320 54.165 190.085 54.305 ;
        RECT 189.320 54.120 189.610 54.165 ;
        RECT 189.765 54.105 190.085 54.165 ;
        RECT 204.485 54.105 204.805 54.365 ;
        RECT 210.005 54.305 210.325 54.365 ;
        RECT 210.480 54.305 210.770 54.350 ;
        RECT 210.005 54.165 210.770 54.305 ;
        RECT 210.005 54.105 210.325 54.165 ;
        RECT 210.480 54.120 210.770 54.165 ;
        RECT 210.925 54.305 211.245 54.365 ;
        RECT 210.925 54.165 217.595 54.305 ;
        RECT 210.925 54.105 211.245 54.165 ;
        RECT 166.730 53.965 167.020 54.010 ;
        RECT 168.620 53.965 168.910 54.010 ;
        RECT 171.740 53.965 172.030 54.010 ;
        RECT 175.505 53.965 175.825 54.025 ;
        RECT 166.730 53.825 172.030 53.965 ;
        RECT 166.730 53.780 167.020 53.825 ;
        RECT 168.620 53.780 168.910 53.825 ;
        RECT 171.740 53.780 172.030 53.825 ;
        RECT 172.375 53.825 175.825 53.965 ;
        RECT 167.240 53.625 167.530 53.670 ;
        RECT 172.375 53.625 172.515 53.825 ;
        RECT 175.505 53.765 175.825 53.825 ;
        RECT 176.885 53.765 177.205 54.025 ;
        RECT 184.260 53.965 184.550 54.010 ;
        RECT 184.705 53.965 185.025 54.025 ;
        RECT 190.240 53.965 190.530 54.010 ;
        RECT 196.205 53.965 196.525 54.025 ;
        RECT 184.260 53.825 187.235 53.965 ;
        RECT 184.260 53.780 184.550 53.825 ;
        RECT 184.705 53.765 185.025 53.825 ;
        RECT 167.240 53.485 172.515 53.625 ;
        RECT 167.240 53.440 167.530 53.485 ;
        RECT 174.600 53.440 174.890 53.670 ;
        RECT 187.095 53.625 187.235 53.825 ;
        RECT 190.240 53.825 196.525 53.965 ;
        RECT 190.240 53.780 190.530 53.825 ;
        RECT 187.480 53.625 187.770 53.670 ;
        RECT 187.095 53.485 187.770 53.625 ;
        RECT 187.480 53.440 187.770 53.485 ;
        RECT 165.845 53.085 166.165 53.345 ;
        RECT 166.325 53.285 166.615 53.330 ;
        RECT 168.160 53.285 168.450 53.330 ;
        RECT 171.740 53.285 172.030 53.330 ;
        RECT 166.325 53.145 172.030 53.285 ;
        RECT 166.325 53.100 166.615 53.145 ;
        RECT 168.160 53.100 168.450 53.145 ;
        RECT 171.740 53.100 172.030 53.145 ;
        RECT 172.820 52.990 173.110 53.305 ;
        RECT 174.675 53.285 174.815 53.440 ;
        RECT 187.925 53.425 188.245 53.685 ;
        RECT 191.235 53.670 191.375 53.825 ;
        RECT 196.205 53.765 196.525 53.825 ;
        RECT 211.810 53.965 212.100 54.010 ;
        RECT 213.700 53.965 213.990 54.010 ;
        RECT 216.820 53.965 217.110 54.010 ;
        RECT 211.810 53.825 217.110 53.965 ;
        RECT 217.455 53.965 217.595 54.165 ;
        RECT 219.665 54.105 219.985 54.365 ;
        RECT 229.785 54.305 230.105 54.365 ;
        RECT 233.940 54.305 234.230 54.350 ;
        RECT 229.785 54.165 234.230 54.305 ;
        RECT 229.785 54.105 230.105 54.165 ;
        RECT 233.940 54.120 234.230 54.165 ;
        RECT 234.385 54.305 234.705 54.365 ;
        RECT 255.545 54.305 255.865 54.365 ;
        RECT 234.385 54.165 255.865 54.305 ;
        RECT 234.385 54.105 234.705 54.165 ;
        RECT 255.545 54.105 255.865 54.165 ;
        RECT 261.065 54.105 261.385 54.365 ;
        RECT 299.245 54.305 299.565 54.365 ;
        RECT 302.020 54.305 302.310 54.350 ;
        RECT 299.245 54.165 302.310 54.305 ;
        RECT 299.245 54.105 299.565 54.165 ;
        RECT 302.020 54.120 302.310 54.165 ;
        RECT 227.945 53.965 228.265 54.025 ;
        RECT 233.005 53.965 233.325 54.025 ;
        RECT 217.455 53.825 228.265 53.965 ;
        RECT 211.810 53.780 212.100 53.825 ;
        RECT 213.700 53.780 213.990 53.825 ;
        RECT 216.820 53.780 217.110 53.825 ;
        RECT 227.945 53.765 228.265 53.825 ;
        RECT 229.875 53.825 233.325 53.965 ;
        RECT 229.875 53.685 230.015 53.825 ;
        RECT 233.005 53.765 233.325 53.825 ;
        RECT 233.465 53.965 233.785 54.025 ;
        RECT 247.725 53.965 248.045 54.025 ;
        RECT 233.465 53.825 248.045 53.965 ;
        RECT 233.465 53.765 233.785 53.825 ;
        RECT 247.725 53.765 248.045 53.825 ;
        RECT 250.960 53.965 251.250 54.010 ;
        RECT 263.365 53.965 263.685 54.025 ;
        RECT 250.960 53.825 263.685 53.965 ;
        RECT 250.960 53.780 251.250 53.825 ;
        RECT 263.365 53.765 263.685 53.825 ;
        RECT 263.940 53.965 264.230 54.010 ;
        RECT 267.060 53.965 267.350 54.010 ;
        RECT 268.950 53.965 269.240 54.010 ;
        RECT 263.940 53.825 269.240 53.965 ;
        RECT 263.940 53.780 264.230 53.825 ;
        RECT 267.060 53.780 267.350 53.825 ;
        RECT 268.950 53.780 269.240 53.825 ;
        RECT 290.505 53.965 290.825 54.025 ;
        RECT 304.780 53.965 305.070 54.010 ;
        RECT 290.505 53.825 305.070 53.965 ;
        RECT 290.505 53.765 290.825 53.825 ;
        RECT 304.780 53.780 305.070 53.825 ;
        RECT 191.160 53.440 191.450 53.670 ;
        RECT 193.460 53.625 193.750 53.670 ;
        RECT 196.680 53.625 196.970 53.670 ;
        RECT 207.245 53.625 207.565 53.685 ;
        RECT 210.940 53.625 211.230 53.670 ;
        RECT 220.125 53.625 220.445 53.685 ;
        RECT 193.460 53.485 195.975 53.625 ;
        RECT 193.460 53.440 193.750 53.485 ;
        RECT 175.980 53.285 176.270 53.330 ;
        RECT 174.675 53.145 176.270 53.285 ;
        RECT 175.980 53.100 176.270 53.145 ;
        RECT 182.865 53.285 183.185 53.345 ;
        RECT 185.640 53.285 185.930 53.330 ;
        RECT 187.005 53.285 187.325 53.345 ;
        RECT 182.865 53.145 187.325 53.285 ;
        RECT 188.015 53.285 188.155 53.425 ;
        RECT 188.015 53.145 188.615 53.285 ;
        RECT 182.865 53.085 183.185 53.145 ;
        RECT 185.640 53.100 185.930 53.145 ;
        RECT 187.005 53.085 187.325 53.145 ;
        RECT 169.520 52.945 170.170 52.990 ;
        RECT 172.820 52.945 173.410 52.990 ;
        RECT 174.125 52.945 174.445 53.005 ;
        RECT 169.520 52.805 174.445 52.945 ;
        RECT 169.520 52.760 170.170 52.805 ;
        RECT 173.120 52.760 173.410 52.805 ;
        RECT 174.125 52.745 174.445 52.805 ;
        RECT 183.325 52.945 183.645 53.005 ;
        RECT 186.100 52.945 186.390 52.990 ;
        RECT 187.465 52.945 187.785 53.005 ;
        RECT 183.325 52.805 187.785 52.945 ;
        RECT 183.325 52.745 183.645 52.805 ;
        RECT 186.100 52.760 186.390 52.805 ;
        RECT 187.465 52.745 187.785 52.805 ;
        RECT 183.785 52.605 184.105 52.665 ;
        RECT 185.165 52.605 185.485 52.665 ;
        RECT 183.785 52.465 185.485 52.605 ;
        RECT 188.475 52.605 188.615 53.145 ;
        RECT 191.605 53.085 191.925 53.345 ;
        RECT 192.065 53.085 192.385 53.345 ;
        RECT 195.835 53.330 195.975 53.485 ;
        RECT 196.680 53.485 202.875 53.625 ;
        RECT 196.680 53.440 196.970 53.485 ;
        RECT 192.540 53.100 192.830 53.330 ;
        RECT 195.300 53.100 195.590 53.330 ;
        RECT 195.760 53.285 196.050 53.330 ;
        RECT 197.140 53.285 197.430 53.330 ;
        RECT 195.760 53.145 197.430 53.285 ;
        RECT 195.760 53.100 196.050 53.145 ;
        RECT 197.140 53.100 197.430 53.145 ;
        RECT 189.305 52.605 189.625 52.665 ;
        RECT 192.615 52.605 192.755 53.100 ;
        RECT 193.905 52.945 194.225 53.005 ;
        RECT 195.375 52.945 195.515 53.100 ;
        RECT 198.505 53.085 198.825 53.345 ;
        RECT 198.965 53.085 199.285 53.345 ;
        RECT 202.735 53.330 202.875 53.485 ;
        RECT 207.245 53.485 220.445 53.625 ;
        RECT 207.245 53.425 207.565 53.485 ;
        RECT 210.940 53.440 211.230 53.485 ;
        RECT 220.125 53.425 220.445 53.485 ;
        RECT 229.785 53.425 230.105 53.685 ;
        RECT 230.245 53.625 230.565 53.685 ;
        RECT 231.180 53.625 231.470 53.670 ;
        RECT 232.545 53.625 232.865 53.685 ;
        RECT 242.205 53.625 242.525 53.685 ;
        RECT 254.625 53.625 254.945 53.685 ;
        RECT 259.240 53.625 259.530 53.670 ;
        RECT 267.965 53.625 268.285 53.685 ;
        RECT 269.820 53.625 270.110 53.670 ;
        RECT 230.245 53.485 232.865 53.625 ;
        RECT 230.245 53.425 230.565 53.485 ;
        RECT 231.180 53.440 231.470 53.485 ;
        RECT 232.545 53.425 232.865 53.485 ;
        RECT 235.855 53.485 242.525 53.625 ;
        RECT 202.660 53.285 202.950 53.330 ;
        RECT 208.625 53.285 208.945 53.345 ;
        RECT 202.660 53.145 208.945 53.285 ;
        RECT 202.660 53.100 202.950 53.145 ;
        RECT 208.625 53.085 208.945 53.145 ;
        RECT 211.405 53.285 211.695 53.330 ;
        RECT 213.240 53.285 213.530 53.330 ;
        RECT 216.820 53.285 217.110 53.330 ;
        RECT 211.405 53.145 217.110 53.285 ;
        RECT 211.405 53.100 211.695 53.145 ;
        RECT 213.240 53.100 213.530 53.145 ;
        RECT 216.820 53.100 217.110 53.145 ;
        RECT 198.595 52.945 198.735 53.085 ;
        RECT 193.905 52.805 198.735 52.945 ;
        RECT 193.905 52.745 194.225 52.805 ;
        RECT 203.565 52.745 203.885 53.005 ;
        RECT 209.560 52.945 209.850 52.990 ;
        RECT 210.465 52.945 210.785 53.005 ;
        RECT 209.560 52.805 210.785 52.945 ;
        RECT 209.560 52.760 209.850 52.805 ;
        RECT 210.465 52.745 210.785 52.805 ;
        RECT 212.305 52.745 212.625 53.005 ;
        RECT 217.900 52.990 218.190 53.305 ;
        RECT 218.745 53.285 219.065 53.345 ;
        RECT 227.040 53.285 227.330 53.330 ;
        RECT 235.855 53.285 235.995 53.485 ;
        RECT 242.205 53.425 242.525 53.485 ;
        RECT 247.355 53.485 270.110 53.625 ;
        RECT 218.745 53.145 235.995 53.285 ;
        RECT 218.745 53.085 219.065 53.145 ;
        RECT 227.040 53.100 227.330 53.145 ;
        RECT 236.225 53.085 236.545 53.345 ;
        RECT 237.145 53.085 237.465 53.345 ;
        RECT 237.620 53.100 237.910 53.330 ;
        RECT 214.600 52.945 215.250 52.990 ;
        RECT 217.900 52.945 218.490 52.990 ;
        RECT 223.345 52.945 223.665 53.005 ;
        RECT 226.120 52.945 226.410 52.990 ;
        RECT 214.600 52.805 223.115 52.945 ;
        RECT 214.600 52.760 215.250 52.805 ;
        RECT 218.200 52.760 218.490 52.805 ;
        RECT 188.475 52.465 192.755 52.605 ;
        RECT 214.145 52.605 214.465 52.665 ;
        RECT 218.835 52.605 218.975 52.805 ;
        RECT 214.145 52.465 218.975 52.605 ;
        RECT 222.975 52.605 223.115 52.805 ;
        RECT 223.345 52.805 226.410 52.945 ;
        RECT 223.345 52.745 223.665 52.805 ;
        RECT 226.120 52.760 226.410 52.805 ;
        RECT 232.085 52.745 232.405 53.005 ;
        RECT 233.005 52.745 233.325 53.005 ;
        RECT 235.305 52.745 235.625 53.005 ;
        RECT 237.695 52.945 237.835 53.100 ;
        RECT 238.065 53.085 238.385 53.345 ;
        RECT 238.985 53.085 239.305 53.345 ;
        RECT 242.295 52.945 242.435 53.425 ;
        RECT 243.585 53.085 243.905 53.345 ;
        RECT 247.355 53.330 247.495 53.485 ;
        RECT 254.625 53.425 254.945 53.485 ;
        RECT 259.240 53.440 259.530 53.485 ;
        RECT 267.965 53.425 268.285 53.485 ;
        RECT 269.820 53.440 270.110 53.485 ;
        RECT 279.925 53.625 280.245 53.685 ;
        RECT 284.080 53.625 284.370 53.670 ;
        RECT 279.925 53.485 284.370 53.625 ;
        RECT 279.925 53.425 280.245 53.485 ;
        RECT 284.080 53.440 284.370 53.485 ;
        RECT 308.905 53.425 309.225 53.685 ;
        RECT 247.280 53.100 247.570 53.330 ;
        RECT 247.725 53.085 248.045 53.345 ;
        RECT 255.100 53.285 255.390 53.330 ;
        RECT 256.005 53.285 256.325 53.345 ;
        RECT 248.275 53.145 256.325 53.285 ;
        RECT 248.275 52.945 248.415 53.145 ;
        RECT 255.100 53.100 255.390 53.145 ;
        RECT 256.005 53.085 256.325 53.145 ;
        RECT 237.695 52.805 241.975 52.945 ;
        RECT 242.295 52.805 248.415 52.945 ;
        RECT 252.325 52.945 252.645 53.005 ;
        RECT 253.720 52.945 254.010 52.990 ;
        RECT 252.325 52.805 254.010 52.945 ;
        RECT 225.645 52.605 225.965 52.665 ;
        RECT 222.975 52.465 225.965 52.605 ;
        RECT 183.785 52.405 184.105 52.465 ;
        RECT 185.165 52.405 185.485 52.465 ;
        RECT 189.305 52.405 189.625 52.465 ;
        RECT 214.145 52.405 214.465 52.465 ;
        RECT 225.645 52.405 225.965 52.465 ;
        RECT 240.840 52.605 241.130 52.650 ;
        RECT 241.285 52.605 241.605 52.665 ;
        RECT 240.840 52.465 241.605 52.605 ;
        RECT 241.835 52.605 241.975 52.805 ;
        RECT 252.325 52.745 252.645 52.805 ;
        RECT 253.720 52.760 254.010 52.805 ;
        RECT 254.165 52.945 254.485 53.005 ;
        RECT 254.640 52.945 254.930 52.990 ;
        RECT 254.165 52.805 254.930 52.945 ;
        RECT 254.165 52.745 254.485 52.805 ;
        RECT 254.640 52.760 254.930 52.805 ;
        RECT 259.685 52.945 260.005 53.005 ;
        RECT 262.860 52.990 263.150 53.305 ;
        RECT 263.940 53.285 264.230 53.330 ;
        RECT 267.520 53.285 267.810 53.330 ;
        RECT 269.355 53.285 269.645 53.330 ;
        RECT 263.940 53.145 269.645 53.285 ;
        RECT 263.940 53.100 264.230 53.145 ;
        RECT 267.520 53.100 267.810 53.145 ;
        RECT 269.355 53.100 269.645 53.145 ;
        RECT 270.725 53.285 271.045 53.345 ;
        RECT 273.040 53.285 273.330 53.330 ;
        RECT 270.725 53.145 273.330 53.285 ;
        RECT 270.725 53.085 271.045 53.145 ;
        RECT 273.040 53.100 273.330 53.145 ;
        RECT 279.465 53.285 279.785 53.345 ;
        RECT 283.620 53.285 283.910 53.330 ;
        RECT 279.465 53.145 283.910 53.285 ;
        RECT 279.465 53.085 279.785 53.145 ;
        RECT 283.620 53.100 283.910 53.145 ;
        RECT 286.380 53.285 286.670 53.330 ;
        RECT 287.285 53.285 287.605 53.345 ;
        RECT 286.380 53.145 287.605 53.285 ;
        RECT 286.380 53.100 286.670 53.145 ;
        RECT 287.285 53.085 287.605 53.145 ;
        RECT 301.560 53.285 301.850 53.330 ;
        RECT 303.385 53.285 303.705 53.345 ;
        RECT 301.560 53.145 303.705 53.285 ;
        RECT 301.560 53.100 301.850 53.145 ;
        RECT 303.385 53.085 303.705 53.145 ;
        RECT 305.685 53.085 306.005 53.345 ;
        RECT 262.560 52.945 263.150 52.990 ;
        RECT 265.800 52.945 266.450 52.990 ;
        RECT 259.685 52.805 266.450 52.945 ;
        RECT 259.685 52.745 260.005 52.805 ;
        RECT 262.560 52.760 262.850 52.805 ;
        RECT 265.800 52.760 266.450 52.805 ;
        RECT 268.440 52.945 268.730 52.990 ;
        RECT 270.280 52.945 270.570 52.990 ;
        RECT 268.440 52.805 270.570 52.945 ;
        RECT 268.440 52.760 268.730 52.805 ;
        RECT 270.280 52.760 270.570 52.805 ;
        RECT 278.545 52.945 278.865 53.005 ;
        RECT 300.165 52.945 300.485 53.005 ;
        RECT 278.545 52.805 300.485 52.945 ;
        RECT 278.545 52.745 278.865 52.805 ;
        RECT 300.165 52.745 300.485 52.805 ;
        RECT 250.025 52.605 250.345 52.665 ;
        RECT 241.835 52.465 250.345 52.605 ;
        RECT 240.840 52.420 241.130 52.465 ;
        RECT 241.285 52.405 241.605 52.465 ;
        RECT 250.025 52.405 250.345 52.465 ;
        RECT 251.405 52.605 251.725 52.665 ;
        RECT 252.800 52.605 253.090 52.650 ;
        RECT 251.405 52.465 253.090 52.605 ;
        RECT 251.405 52.405 251.725 52.465 ;
        RECT 252.800 52.420 253.090 52.465 ;
        RECT 255.085 52.605 255.405 52.665 ;
        RECT 256.465 52.605 256.785 52.665 ;
        RECT 255.085 52.465 256.785 52.605 ;
        RECT 255.085 52.405 255.405 52.465 ;
        RECT 256.465 52.405 256.785 52.465 ;
        RECT 280.385 52.605 280.705 52.665 ;
        RECT 281.320 52.605 281.610 52.650 ;
        RECT 280.385 52.465 281.610 52.605 ;
        RECT 280.385 52.405 280.705 52.465 ;
        RECT 281.320 52.420 281.610 52.465 ;
        RECT 283.160 52.605 283.450 52.650 ;
        RECT 284.525 52.605 284.845 52.665 ;
        RECT 287.745 52.605 288.065 52.665 ;
        RECT 283.160 52.465 288.065 52.605 ;
        RECT 283.160 52.420 283.450 52.465 ;
        RECT 284.525 52.405 284.845 52.465 ;
        RECT 287.745 52.405 288.065 52.465 ;
        RECT 306.160 52.605 306.450 52.650 ;
        RECT 307.065 52.605 307.385 52.665 ;
        RECT 306.160 52.465 307.385 52.605 ;
        RECT 306.160 52.420 306.450 52.465 ;
        RECT 307.065 52.405 307.385 52.465 ;
        RECT 162.095 51.785 311.135 52.265 ;
        RECT 172.285 51.585 172.605 51.645 ;
        RECT 179.645 51.585 179.965 51.645 ;
        RECT 184.260 51.585 184.550 51.630 ;
        RECT 172.285 51.445 184.550 51.585 ;
        RECT 172.285 51.385 172.605 51.445 ;
        RECT 179.645 51.385 179.965 51.445 ;
        RECT 184.260 51.400 184.550 51.445 ;
        RECT 188.860 51.585 189.150 51.630 ;
        RECT 192.065 51.585 192.385 51.645 ;
        RECT 188.860 51.445 192.385 51.585 ;
        RECT 188.860 51.400 189.150 51.445 ;
        RECT 192.065 51.385 192.385 51.445 ;
        RECT 197.125 51.585 197.445 51.645 ;
        RECT 210.465 51.585 210.785 51.645 ;
        RECT 213.240 51.585 213.530 51.630 ;
        RECT 213.685 51.585 214.005 51.645 ;
        RECT 252.785 51.585 253.105 51.645 ;
        RECT 283.605 51.585 283.925 51.645 ;
        RECT 197.125 51.445 198.735 51.585 ;
        RECT 197.125 51.385 197.445 51.445 ;
        RECT 169.980 51.245 170.630 51.290 ;
        RECT 173.580 51.245 173.870 51.290 ;
        RECT 174.125 51.245 174.445 51.305 ;
        RECT 176.425 51.245 176.745 51.305 ;
        RECT 169.980 51.105 176.745 51.245 ;
        RECT 169.980 51.060 170.630 51.105 ;
        RECT 173.280 51.060 173.870 51.105 ;
        RECT 166.785 50.905 167.075 50.950 ;
        RECT 168.620 50.905 168.910 50.950 ;
        RECT 172.200 50.905 172.490 50.950 ;
        RECT 166.785 50.765 172.490 50.905 ;
        RECT 166.785 50.720 167.075 50.765 ;
        RECT 168.620 50.720 168.910 50.765 ;
        RECT 172.200 50.720 172.490 50.765 ;
        RECT 173.280 50.745 173.570 51.060 ;
        RECT 174.125 51.045 174.445 51.105 ;
        RECT 176.425 51.045 176.745 51.105 ;
        RECT 177.820 51.245 178.110 51.290 ;
        RECT 180.105 51.245 180.425 51.305 ;
        RECT 185.165 51.290 185.485 51.305 ;
        RECT 177.820 51.105 180.425 51.245 ;
        RECT 177.820 51.060 178.110 51.105 ;
        RECT 175.965 50.905 176.285 50.965 ;
        RECT 175.135 50.765 176.285 50.905 ;
        RECT 166.305 50.365 166.625 50.625 ;
        RECT 167.700 50.565 167.990 50.610 ;
        RECT 170.905 50.565 171.225 50.625 ;
        RECT 175.135 50.610 175.275 50.765 ;
        RECT 175.965 50.705 176.285 50.765 ;
        RECT 167.700 50.425 171.225 50.565 ;
        RECT 167.700 50.380 167.990 50.425 ;
        RECT 170.905 50.365 171.225 50.425 ;
        RECT 175.060 50.380 175.350 50.610 ;
        RECT 167.190 50.225 167.480 50.270 ;
        RECT 169.080 50.225 169.370 50.270 ;
        RECT 172.200 50.225 172.490 50.270 ;
        RECT 167.190 50.085 172.490 50.225 ;
        RECT 167.190 50.040 167.480 50.085 ;
        RECT 169.080 50.040 169.370 50.085 ;
        RECT 172.200 50.040 172.490 50.085 ;
        RECT 172.745 49.885 173.065 49.945 ;
        RECT 177.895 49.885 178.035 51.060 ;
        RECT 180.105 51.045 180.425 51.105 ;
        RECT 185.055 51.060 185.485 51.290 ;
        RECT 186.100 51.245 186.390 51.290 ;
        RECT 189.305 51.245 189.625 51.305 ;
        RECT 193.445 51.245 193.765 51.305 ;
        RECT 193.920 51.245 194.210 51.290 ;
        RECT 186.100 51.105 189.075 51.245 ;
        RECT 186.100 51.060 186.390 51.105 ;
        RECT 185.165 51.045 185.485 51.060 ;
        RECT 182.865 50.705 183.185 50.965 ;
        RECT 183.325 50.905 183.645 50.965 ;
        RECT 183.800 50.905 184.090 50.950 ;
        RECT 188.400 50.905 188.690 50.950 ;
        RECT 183.325 50.765 184.090 50.905 ;
        RECT 183.325 50.705 183.645 50.765 ;
        RECT 183.800 50.720 184.090 50.765 ;
        RECT 185.255 50.765 188.690 50.905 ;
        RECT 182.955 50.565 183.095 50.705 ;
        RECT 185.255 50.565 185.395 50.765 ;
        RECT 188.400 50.720 188.690 50.765 ;
        RECT 182.955 50.425 185.395 50.565 ;
        RECT 185.640 50.380 185.930 50.610 ;
        RECT 187.005 50.565 187.325 50.625 ;
        RECT 187.480 50.565 187.770 50.610 ;
        RECT 187.005 50.425 187.770 50.565 ;
        RECT 183.800 50.225 184.090 50.270 ;
        RECT 185.715 50.225 185.855 50.380 ;
        RECT 187.005 50.365 187.325 50.425 ;
        RECT 187.480 50.380 187.770 50.425 ;
        RECT 183.800 50.085 185.855 50.225 ;
        RECT 188.475 50.225 188.615 50.720 ;
        RECT 188.935 50.565 189.075 51.105 ;
        RECT 189.305 51.105 194.210 51.245 ;
        RECT 189.305 51.045 189.625 51.105 ;
        RECT 193.445 51.045 193.765 51.105 ;
        RECT 193.920 51.060 194.210 51.105 ;
        RECT 196.680 51.245 196.970 51.290 ;
        RECT 198.045 51.245 198.365 51.305 ;
        RECT 196.680 51.105 198.365 51.245 ;
        RECT 198.595 51.245 198.735 51.445 ;
        RECT 210.465 51.445 214.005 51.585 ;
        RECT 210.465 51.385 210.785 51.445 ;
        RECT 213.240 51.400 213.530 51.445 ;
        RECT 213.685 51.385 214.005 51.445 ;
        RECT 247.815 51.445 253.105 51.585 ;
        RECT 198.960 51.245 199.610 51.290 ;
        RECT 202.560 51.245 202.850 51.290 ;
        RECT 207.245 51.245 207.565 51.305 ;
        RECT 198.595 51.105 202.850 51.245 ;
        RECT 196.680 51.060 196.970 51.105 ;
        RECT 198.045 51.045 198.365 51.105 ;
        RECT 198.960 51.060 199.610 51.105 ;
        RECT 202.260 51.060 202.850 51.105 ;
        RECT 204.575 51.105 207.565 51.245 ;
        RECT 190.225 50.705 190.545 50.965 ;
        RECT 195.765 50.905 196.055 50.950 ;
        RECT 197.600 50.905 197.890 50.950 ;
        RECT 201.180 50.905 201.470 50.950 ;
        RECT 195.765 50.765 201.470 50.905 ;
        RECT 195.765 50.720 196.055 50.765 ;
        RECT 197.600 50.720 197.890 50.765 ;
        RECT 201.180 50.720 201.470 50.765 ;
        RECT 202.260 50.745 202.550 51.060 ;
        RECT 204.575 50.950 204.715 51.105 ;
        RECT 207.245 51.045 207.565 51.105 ;
        RECT 208.160 51.245 208.810 51.290 ;
        RECT 211.760 51.245 212.050 51.290 ;
        RECT 212.305 51.245 212.625 51.305 ;
        RECT 214.145 51.245 214.465 51.305 ;
        RECT 208.160 51.105 214.465 51.245 ;
        RECT 208.160 51.060 208.810 51.105 ;
        RECT 211.460 51.060 212.050 51.105 ;
        RECT 204.500 50.720 204.790 50.950 ;
        RECT 204.965 50.905 205.255 50.950 ;
        RECT 206.800 50.905 207.090 50.950 ;
        RECT 210.380 50.905 210.670 50.950 ;
        RECT 204.965 50.765 210.670 50.905 ;
        RECT 204.965 50.720 205.255 50.765 ;
        RECT 206.800 50.720 207.090 50.765 ;
        RECT 210.380 50.720 210.670 50.765 ;
        RECT 211.460 50.745 211.750 51.060 ;
        RECT 212.305 51.045 212.625 51.105 ;
        RECT 214.145 51.045 214.465 51.105 ;
        RECT 214.605 51.245 214.925 51.305 ;
        RECT 217.840 51.245 218.130 51.290 ;
        RECT 218.745 51.245 219.065 51.305 ;
        RECT 214.605 51.105 219.065 51.245 ;
        RECT 214.605 51.045 214.925 51.105 ;
        RECT 217.840 51.060 218.130 51.105 ;
        RECT 218.745 51.045 219.065 51.105 ;
        RECT 219.665 51.245 219.985 51.305 ;
        RECT 221.980 51.245 222.270 51.290 ;
        RECT 223.345 51.245 223.665 51.305 ;
        RECT 219.665 51.105 223.665 51.245 ;
        RECT 219.665 51.045 219.985 51.105 ;
        RECT 221.980 51.060 222.270 51.105 ;
        RECT 223.345 51.045 223.665 51.105 ;
        RECT 220.125 50.905 220.445 50.965 ;
        RECT 223.820 50.905 224.110 50.950 ;
        RECT 230.245 50.905 230.565 50.965 ;
        RECT 220.125 50.765 230.565 50.905 ;
        RECT 220.125 50.705 220.445 50.765 ;
        RECT 223.820 50.720 224.110 50.765 ;
        RECT 230.245 50.705 230.565 50.765 ;
        RECT 236.225 50.905 236.545 50.965 ;
        RECT 247.815 50.950 247.955 51.445 ;
        RECT 252.785 51.385 253.105 51.445 ;
        RECT 279.095 51.445 288.435 51.585 ;
        RECT 256.005 51.045 256.325 51.305 ;
        RECT 260.160 51.245 260.450 51.290 ;
        RECT 262.905 51.245 263.225 51.305 ;
        RECT 267.045 51.245 267.365 51.305 ;
        RECT 260.160 51.105 267.365 51.245 ;
        RECT 260.160 51.060 260.450 51.105 ;
        RECT 262.905 51.045 263.225 51.105 ;
        RECT 267.045 51.045 267.365 51.105 ;
        RECT 271.640 51.245 272.290 51.290 ;
        RECT 275.240 51.245 275.530 51.290 ;
        RECT 276.705 51.245 277.025 51.305 ;
        RECT 271.640 51.105 277.025 51.245 ;
        RECT 271.640 51.060 272.290 51.105 ;
        RECT 274.940 51.060 275.530 51.105 ;
        RECT 247.740 50.905 248.030 50.950 ;
        RECT 236.225 50.765 248.030 50.905 ;
        RECT 236.225 50.705 236.545 50.765 ;
        RECT 247.740 50.720 248.030 50.765 ;
        RECT 249.565 50.905 249.885 50.965 ;
        RECT 250.500 50.905 250.790 50.950 ;
        RECT 251.405 50.905 251.725 50.965 ;
        RECT 249.565 50.765 250.255 50.905 ;
        RECT 249.565 50.705 249.885 50.765 ;
        RECT 193.905 50.565 194.225 50.625 ;
        RECT 188.935 50.425 194.225 50.565 ;
        RECT 193.905 50.365 194.225 50.425 ;
        RECT 195.285 50.365 195.605 50.625 ;
        RECT 205.865 50.365 206.185 50.625 ;
        RECT 238.985 50.365 239.305 50.625 ;
        RECT 244.505 50.365 244.825 50.625 ;
        RECT 248.660 50.380 248.950 50.610 ;
        RECT 249.120 50.565 249.410 50.610 ;
        RECT 250.115 50.565 250.255 50.765 ;
        RECT 250.500 50.765 251.725 50.905 ;
        RECT 250.500 50.720 250.790 50.765 ;
        RECT 251.405 50.705 251.725 50.765 ;
        RECT 252.785 50.705 253.105 50.965 ;
        RECT 253.705 50.705 254.025 50.965 ;
        RECT 254.165 50.705 254.485 50.965 ;
        RECT 254.640 50.720 254.930 50.950 ;
        RECT 255.560 50.905 255.850 50.950 ;
        RECT 256.925 50.905 257.245 50.965 ;
        RECT 255.560 50.765 257.245 50.905 ;
        RECT 255.560 50.720 255.850 50.765 ;
        RECT 254.715 50.565 254.855 50.720 ;
        RECT 256.925 50.705 257.245 50.765 ;
        RECT 266.600 50.720 266.890 50.950 ;
        RECT 255.085 50.565 255.405 50.625 ;
        RECT 249.120 50.425 249.795 50.565 ;
        RECT 250.115 50.425 255.405 50.565 ;
        RECT 249.120 50.380 249.410 50.425 ;
        RECT 189.765 50.225 190.085 50.285 ;
        RECT 188.475 50.085 190.085 50.225 ;
        RECT 183.800 50.040 184.090 50.085 ;
        RECT 189.765 50.025 190.085 50.085 ;
        RECT 196.170 50.225 196.460 50.270 ;
        RECT 198.060 50.225 198.350 50.270 ;
        RECT 201.180 50.225 201.470 50.270 ;
        RECT 196.170 50.085 201.470 50.225 ;
        RECT 196.170 50.040 196.460 50.085 ;
        RECT 198.060 50.040 198.350 50.085 ;
        RECT 201.180 50.040 201.470 50.085 ;
        RECT 205.370 50.225 205.660 50.270 ;
        RECT 207.260 50.225 207.550 50.270 ;
        RECT 210.380 50.225 210.670 50.270 ;
        RECT 205.370 50.085 210.670 50.225 ;
        RECT 205.370 50.040 205.660 50.085 ;
        RECT 207.260 50.040 207.550 50.085 ;
        RECT 210.380 50.040 210.670 50.085 ;
        RECT 225.185 50.225 225.505 50.285 ;
        RECT 248.735 50.225 248.875 50.380 ;
        RECT 225.185 50.085 248.875 50.225 ;
        RECT 249.655 50.225 249.795 50.425 ;
        RECT 255.085 50.365 255.405 50.425 ;
        RECT 256.005 50.565 256.325 50.625 ;
        RECT 263.840 50.565 264.130 50.610 ;
        RECT 256.005 50.425 264.130 50.565 ;
        RECT 256.005 50.365 256.325 50.425 ;
        RECT 263.840 50.380 264.130 50.425 ;
        RECT 261.080 50.225 261.370 50.270 ;
        RECT 249.655 50.085 261.370 50.225 ;
        RECT 225.185 50.025 225.505 50.085 ;
        RECT 261.080 50.040 261.370 50.085 ;
        RECT 262.905 50.225 263.225 50.285 ;
        RECT 266.675 50.225 266.815 50.720 ;
        RECT 267.965 50.705 268.285 50.965 ;
        RECT 268.445 50.905 268.735 50.950 ;
        RECT 270.280 50.905 270.570 50.950 ;
        RECT 273.860 50.905 274.150 50.950 ;
        RECT 268.445 50.765 274.150 50.905 ;
        RECT 268.445 50.720 268.735 50.765 ;
        RECT 270.280 50.720 270.570 50.765 ;
        RECT 273.860 50.720 274.150 50.765 ;
        RECT 274.940 50.745 275.230 51.060 ;
        RECT 276.705 51.045 277.025 51.105 ;
        RECT 269.345 50.365 269.665 50.625 ;
        RECT 276.795 50.565 276.935 51.045 ;
        RECT 279.095 50.950 279.235 51.445 ;
        RECT 283.605 51.385 283.925 51.445 ;
        RECT 280.385 51.045 280.705 51.305 ;
        RECT 288.295 51.290 288.435 51.445 ;
        RECT 282.680 51.245 283.330 51.290 ;
        RECT 286.280 51.245 286.570 51.290 ;
        RECT 282.680 51.105 286.570 51.245 ;
        RECT 282.680 51.060 283.330 51.105 ;
        RECT 285.980 51.060 286.570 51.105 ;
        RECT 288.220 51.060 288.510 51.290 ;
        RECT 299.245 51.245 299.565 51.305 ;
        RECT 302.020 51.245 302.310 51.290 ;
        RECT 305.240 51.245 305.530 51.290 ;
        RECT 299.245 51.105 305.530 51.245 ;
        RECT 279.020 50.720 279.310 50.950 ;
        RECT 279.485 50.905 279.775 50.950 ;
        RECT 281.320 50.905 281.610 50.950 ;
        RECT 284.900 50.905 285.190 50.950 ;
        RECT 279.485 50.765 285.190 50.905 ;
        RECT 279.485 50.720 279.775 50.765 ;
        RECT 281.320 50.720 281.610 50.765 ;
        RECT 284.900 50.720 285.190 50.765 ;
        RECT 285.980 50.745 286.270 51.060 ;
        RECT 299.245 51.045 299.565 51.105 ;
        RECT 302.020 51.060 302.310 51.105 ;
        RECT 305.240 51.060 305.530 51.105 ;
        RECT 306.160 51.245 306.450 51.290 ;
        RECT 308.000 51.245 308.290 51.290 ;
        RECT 306.160 51.105 308.290 51.245 ;
        RECT 306.160 51.060 306.450 51.105 ;
        RECT 308.000 51.060 308.290 51.105 ;
        RECT 303.840 50.905 304.130 50.950 ;
        RECT 306.160 50.905 306.375 51.060 ;
        RECT 308.920 50.905 309.210 50.950 ;
        RECT 303.840 50.765 306.375 50.905 ;
        RECT 306.695 50.765 309.210 50.905 ;
        RECT 283.605 50.565 283.925 50.625 ;
        RECT 285.995 50.565 286.135 50.745 ;
        RECT 303.840 50.720 304.130 50.765 ;
        RECT 286.365 50.565 286.685 50.625 ;
        RECT 276.795 50.425 286.685 50.565 ;
        RECT 283.605 50.365 283.925 50.425 ;
        RECT 286.365 50.365 286.685 50.425 ;
        RECT 287.745 50.365 288.065 50.625 ;
        RECT 305.685 50.565 306.005 50.625 ;
        RECT 306.695 50.565 306.835 50.765 ;
        RECT 308.920 50.720 309.210 50.765 ;
        RECT 305.685 50.425 306.835 50.565 ;
        RECT 305.685 50.365 306.005 50.425 ;
        RECT 307.065 50.365 307.385 50.625 ;
        RECT 267.965 50.225 268.285 50.285 ;
        RECT 262.905 50.085 268.285 50.225 ;
        RECT 262.905 50.025 263.225 50.085 ;
        RECT 267.965 50.025 268.285 50.085 ;
        RECT 268.850 50.225 269.140 50.270 ;
        RECT 270.740 50.225 271.030 50.270 ;
        RECT 273.860 50.225 274.150 50.270 ;
        RECT 268.850 50.085 274.150 50.225 ;
        RECT 268.850 50.040 269.140 50.085 ;
        RECT 270.740 50.040 271.030 50.085 ;
        RECT 273.860 50.040 274.150 50.085 ;
        RECT 279.890 50.225 280.180 50.270 ;
        RECT 281.780 50.225 282.070 50.270 ;
        RECT 284.900 50.225 285.190 50.270 ;
        RECT 279.890 50.085 285.190 50.225 ;
        RECT 279.890 50.040 280.180 50.085 ;
        RECT 281.780 50.040 282.070 50.085 ;
        RECT 284.900 50.040 285.190 50.085 ;
        RECT 303.860 50.225 304.150 50.270 ;
        RECT 306.620 50.225 306.910 50.270 ;
        RECT 308.460 50.225 308.750 50.270 ;
        RECT 303.860 50.085 308.750 50.225 ;
        RECT 303.860 50.040 304.150 50.085 ;
        RECT 306.620 50.040 306.910 50.085 ;
        RECT 308.460 50.040 308.750 50.085 ;
        RECT 172.745 49.745 178.035 49.885 ;
        RECT 203.565 49.885 203.885 49.945 ;
        RECT 204.040 49.885 204.330 49.930 ;
        RECT 210.925 49.885 211.245 49.945 ;
        RECT 203.565 49.745 211.245 49.885 ;
        RECT 172.745 49.685 173.065 49.745 ;
        RECT 203.565 49.685 203.885 49.745 ;
        RECT 204.040 49.700 204.330 49.745 ;
        RECT 210.925 49.685 211.245 49.745 ;
        RECT 211.385 49.885 211.705 49.945 ;
        RECT 220.585 49.885 220.905 49.945 ;
        RECT 211.385 49.745 220.905 49.885 ;
        RECT 211.385 49.685 211.705 49.745 ;
        RECT 220.585 49.685 220.905 49.745 ;
        RECT 231.625 49.885 231.945 49.945 ;
        RECT 235.780 49.885 236.070 49.930 ;
        RECT 231.625 49.745 236.070 49.885 ;
        RECT 231.625 49.685 231.945 49.745 ;
        RECT 235.780 49.700 236.070 49.745 ;
        RECT 241.760 49.885 242.050 49.930 ;
        RECT 242.665 49.885 242.985 49.945 ;
        RECT 241.760 49.745 242.985 49.885 ;
        RECT 241.760 49.700 242.050 49.745 ;
        RECT 242.665 49.685 242.985 49.745 ;
        RECT 246.805 49.685 247.125 49.945 ;
        RECT 251.880 49.885 252.170 49.930 ;
        RECT 260.145 49.885 260.465 49.945 ;
        RECT 251.880 49.745 260.465 49.885 ;
        RECT 251.880 49.700 252.170 49.745 ;
        RECT 260.145 49.685 260.465 49.745 ;
        RECT 266.125 49.685 266.445 49.945 ;
        RECT 276.720 49.885 277.010 49.930 ;
        RECT 277.165 49.885 277.485 49.945 ;
        RECT 276.720 49.745 277.485 49.885 ;
        RECT 276.720 49.700 277.010 49.745 ;
        RECT 277.165 49.685 277.485 49.745 ;
        RECT 277.625 49.885 277.945 49.945 ;
        RECT 300.180 49.885 300.470 49.930 ;
        RECT 277.625 49.745 300.470 49.885 ;
        RECT 277.625 49.685 277.945 49.745 ;
        RECT 300.180 49.700 300.470 49.745 ;
        RECT 162.095 49.065 311.135 49.545 ;
        RECT 170.905 48.665 171.225 48.925 ;
        RECT 190.225 48.865 190.545 48.925 ;
        RECT 214.605 48.865 214.925 48.925 ;
        RECT 190.225 48.725 214.925 48.865 ;
        RECT 190.225 48.665 190.545 48.725 ;
        RECT 172.285 48.185 172.605 48.245 ;
        RECT 173.680 48.185 173.970 48.230 ;
        RECT 172.285 48.045 173.970 48.185 ;
        RECT 172.285 47.985 172.605 48.045 ;
        RECT 173.680 48.000 173.970 48.045 ;
        RECT 179.660 48.185 179.950 48.230 ;
        RECT 184.705 48.185 185.025 48.245 ;
        RECT 179.660 48.045 185.025 48.185 ;
        RECT 179.660 48.000 179.950 48.045 ;
        RECT 184.705 47.985 185.025 48.045 ;
        RECT 173.220 47.845 173.510 47.890 ;
        RECT 175.045 47.845 175.365 47.905 ;
        RECT 173.220 47.705 175.365 47.845 ;
        RECT 173.220 47.660 173.510 47.705 ;
        RECT 175.045 47.645 175.365 47.705 ;
        RECT 180.105 47.845 180.425 47.905 ;
        RECT 199.515 47.890 199.655 48.725 ;
        RECT 214.605 48.665 214.925 48.725 ;
        RECT 215.525 48.865 215.845 48.925 ;
        RECT 222.900 48.865 223.190 48.910 ;
        RECT 236.685 48.865 237.005 48.925 ;
        RECT 215.525 48.725 237.005 48.865 ;
        RECT 215.525 48.665 215.845 48.725 ;
        RECT 222.900 48.680 223.190 48.725 ;
        RECT 236.685 48.665 237.005 48.725 ;
        RECT 239.000 48.865 239.290 48.910 ;
        RECT 245.885 48.865 246.205 48.925 ;
        RECT 239.000 48.725 246.205 48.865 ;
        RECT 239.000 48.680 239.290 48.725 ;
        RECT 245.885 48.665 246.205 48.725 ;
        RECT 254.165 48.865 254.485 48.925 ;
        RECT 263.840 48.865 264.130 48.910 ;
        RECT 254.165 48.725 264.130 48.865 ;
        RECT 254.165 48.665 254.485 48.725 ;
        RECT 263.840 48.680 264.130 48.725 ;
        RECT 269.345 48.865 269.665 48.925 ;
        RECT 270.740 48.865 271.030 48.910 ;
        RECT 269.345 48.725 271.030 48.865 ;
        RECT 269.345 48.665 269.665 48.725 ;
        RECT 270.740 48.680 271.030 48.725 ;
        RECT 278.545 48.665 278.865 48.925 ;
        RECT 207.820 48.525 208.110 48.570 ;
        RECT 210.940 48.525 211.230 48.570 ;
        RECT 212.830 48.525 213.120 48.570 ;
        RECT 214.145 48.525 214.465 48.585 ;
        RECT 207.820 48.385 213.120 48.525 ;
        RECT 207.820 48.340 208.110 48.385 ;
        RECT 210.940 48.340 211.230 48.385 ;
        RECT 212.830 48.340 213.120 48.385 ;
        RECT 213.315 48.385 214.465 48.525 ;
        RECT 212.320 48.185 212.610 48.230 ;
        RECT 213.315 48.185 213.455 48.385 ;
        RECT 214.145 48.325 214.465 48.385 ;
        RECT 215.030 48.525 215.320 48.570 ;
        RECT 216.920 48.525 217.210 48.570 ;
        RECT 220.040 48.525 220.330 48.570 ;
        RECT 215.030 48.385 220.330 48.525 ;
        RECT 215.030 48.340 215.320 48.385 ;
        RECT 216.920 48.340 217.210 48.385 ;
        RECT 220.040 48.340 220.330 48.385 ;
        RECT 231.130 48.525 231.420 48.570 ;
        RECT 233.020 48.525 233.310 48.570 ;
        RECT 236.140 48.525 236.430 48.570 ;
        RECT 231.130 48.385 236.430 48.525 ;
        RECT 231.130 48.340 231.420 48.385 ;
        RECT 233.020 48.340 233.310 48.385 ;
        RECT 236.140 48.340 236.430 48.385 ;
        RECT 242.170 48.525 242.460 48.570 ;
        RECT 244.060 48.525 244.350 48.570 ;
        RECT 247.180 48.525 247.470 48.570 ;
        RECT 242.170 48.385 247.470 48.525 ;
        RECT 242.170 48.340 242.460 48.385 ;
        RECT 244.060 48.340 244.350 48.385 ;
        RECT 247.180 48.340 247.470 48.385 ;
        RECT 250.040 48.525 250.330 48.570 ;
        RECT 255.510 48.525 255.800 48.570 ;
        RECT 257.400 48.525 257.690 48.570 ;
        RECT 260.520 48.525 260.810 48.570 ;
        RECT 250.040 48.385 255.315 48.525 ;
        RECT 250.040 48.340 250.330 48.385 ;
        RECT 212.320 48.045 213.455 48.185 ;
        RECT 213.700 48.185 213.990 48.230 ;
        RECT 219.205 48.185 219.525 48.245 ;
        RECT 213.700 48.045 219.525 48.185 ;
        RECT 212.320 48.000 212.610 48.045 ;
        RECT 213.700 48.000 213.990 48.045 ;
        RECT 219.205 47.985 219.525 48.045 ;
        RECT 230.245 47.985 230.565 48.245 ;
        RECT 242.665 47.985 242.985 48.245 ;
        RECT 181.040 47.845 181.330 47.890 ;
        RECT 180.105 47.705 181.330 47.845 ;
        RECT 180.105 47.645 180.425 47.705 ;
        RECT 181.040 47.660 181.330 47.705 ;
        RECT 193.920 47.660 194.210 47.890 ;
        RECT 199.440 47.660 199.730 47.890 ;
        RECT 178.740 47.505 179.030 47.550 ;
        RECT 182.865 47.505 183.185 47.565 ;
        RECT 178.740 47.365 183.185 47.505 ;
        RECT 193.995 47.505 194.135 47.660 ;
        RECT 195.745 47.505 196.065 47.565 ;
        RECT 193.995 47.365 196.065 47.505 ;
        RECT 178.740 47.320 179.030 47.365 ;
        RECT 182.865 47.305 183.185 47.365 ;
        RECT 195.745 47.305 196.065 47.365 ;
        RECT 204.025 47.505 204.345 47.565 ;
        RECT 206.740 47.550 207.030 47.865 ;
        RECT 207.820 47.845 208.110 47.890 ;
        RECT 211.400 47.845 211.690 47.890 ;
        RECT 213.235 47.845 213.525 47.890 ;
        RECT 207.820 47.705 213.525 47.845 ;
        RECT 207.820 47.660 208.110 47.705 ;
        RECT 211.400 47.660 211.690 47.705 ;
        RECT 213.235 47.660 213.525 47.705 ;
        RECT 214.160 47.660 214.450 47.890 ;
        RECT 214.625 47.845 214.915 47.890 ;
        RECT 216.460 47.845 216.750 47.890 ;
        RECT 220.040 47.845 220.330 47.890 ;
        RECT 214.625 47.705 220.330 47.845 ;
        RECT 214.625 47.660 214.915 47.705 ;
        RECT 216.460 47.660 216.750 47.705 ;
        RECT 220.040 47.660 220.330 47.705 ;
        RECT 221.120 47.845 221.410 47.865 ;
        RECT 226.105 47.845 226.425 47.905 ;
        RECT 221.120 47.705 226.425 47.845 ;
        RECT 206.440 47.505 207.030 47.550 ;
        RECT 209.680 47.505 210.330 47.550 ;
        RECT 212.305 47.505 212.625 47.565 ;
        RECT 204.025 47.365 205.635 47.505 ;
        RECT 204.025 47.305 204.345 47.365 ;
        RECT 170.905 47.165 171.225 47.225 ;
        RECT 172.745 47.165 173.065 47.225 ;
        RECT 170.905 47.025 173.065 47.165 ;
        RECT 170.905 46.965 171.225 47.025 ;
        RECT 172.745 46.965 173.065 47.025 ;
        RECT 176.885 46.965 177.205 47.225 ;
        RECT 179.200 47.165 179.490 47.210 ;
        RECT 179.645 47.165 179.965 47.225 ;
        RECT 179.200 47.025 179.965 47.165 ;
        RECT 179.200 46.980 179.490 47.025 ;
        RECT 179.645 46.965 179.965 47.025 ;
        RECT 183.785 47.165 184.105 47.225 ;
        RECT 184.260 47.165 184.550 47.210 ;
        RECT 183.785 47.025 184.550 47.165 ;
        RECT 183.785 46.965 184.105 47.025 ;
        RECT 184.260 46.980 184.550 47.025 ;
        RECT 204.945 46.965 205.265 47.225 ;
        RECT 205.495 47.165 205.635 47.365 ;
        RECT 206.440 47.365 212.625 47.505 ;
        RECT 206.440 47.320 206.730 47.365 ;
        RECT 209.680 47.320 210.330 47.365 ;
        RECT 212.305 47.305 212.625 47.365 ;
        RECT 211.385 47.165 211.705 47.225 ;
        RECT 205.495 47.025 211.705 47.165 ;
        RECT 214.235 47.165 214.375 47.660 ;
        RECT 215.540 47.505 215.830 47.550 ;
        RECT 215.985 47.505 216.305 47.565 ;
        RECT 221.120 47.550 221.410 47.705 ;
        RECT 226.105 47.645 226.425 47.705 ;
        RECT 230.725 47.845 231.015 47.890 ;
        RECT 232.560 47.845 232.850 47.890 ;
        RECT 236.140 47.845 236.430 47.890 ;
        RECT 230.725 47.705 236.430 47.845 ;
        RECT 230.725 47.660 231.015 47.705 ;
        RECT 232.560 47.660 232.850 47.705 ;
        RECT 236.140 47.660 236.430 47.705 ;
        RECT 215.540 47.365 216.305 47.505 ;
        RECT 215.540 47.320 215.830 47.365 ;
        RECT 215.985 47.305 216.305 47.365 ;
        RECT 217.820 47.505 218.470 47.550 ;
        RECT 221.120 47.505 221.710 47.550 ;
        RECT 227.485 47.505 227.805 47.565 ;
        RECT 237.220 47.550 237.510 47.865 ;
        RECT 240.365 47.845 240.685 47.905 ;
        RECT 241.300 47.845 241.590 47.890 ;
        RECT 240.365 47.705 241.590 47.845 ;
        RECT 240.365 47.645 240.685 47.705 ;
        RECT 241.300 47.660 241.590 47.705 ;
        RECT 241.765 47.845 242.055 47.890 ;
        RECT 243.600 47.845 243.890 47.890 ;
        RECT 247.180 47.845 247.470 47.890 ;
        RECT 241.765 47.705 247.470 47.845 ;
        RECT 241.765 47.660 242.055 47.705 ;
        RECT 243.600 47.660 243.890 47.705 ;
        RECT 247.180 47.660 247.470 47.705 ;
        RECT 217.820 47.365 221.710 47.505 ;
        RECT 217.820 47.320 218.470 47.365 ;
        RECT 221.420 47.320 221.710 47.365 ;
        RECT 222.515 47.365 227.805 47.505 ;
        RECT 216.445 47.165 216.765 47.225 ;
        RECT 220.125 47.165 220.445 47.225 ;
        RECT 214.235 47.025 220.445 47.165 ;
        RECT 211.385 46.965 211.705 47.025 ;
        RECT 216.445 46.965 216.765 47.025 ;
        RECT 220.125 46.965 220.445 47.025 ;
        RECT 220.585 47.165 220.905 47.225 ;
        RECT 222.515 47.165 222.655 47.365 ;
        RECT 227.485 47.305 227.805 47.365 ;
        RECT 231.640 47.320 231.930 47.550 ;
        RECT 233.920 47.505 234.570 47.550 ;
        RECT 237.220 47.505 237.810 47.550 ;
        RECT 238.065 47.505 238.385 47.565 ;
        RECT 233.920 47.365 238.385 47.505 ;
        RECT 233.920 47.320 234.570 47.365 ;
        RECT 237.520 47.320 237.810 47.365 ;
        RECT 220.585 47.025 222.655 47.165 ;
        RECT 226.565 47.165 226.885 47.225 ;
        RECT 231.715 47.165 231.855 47.320 ;
        RECT 238.065 47.305 238.385 47.365 ;
        RECT 242.665 47.505 242.985 47.565 ;
        RECT 244.965 47.550 245.285 47.565 ;
        RECT 248.260 47.550 248.550 47.865 ;
        RECT 244.960 47.505 245.610 47.550 ;
        RECT 248.260 47.505 248.850 47.550 ;
        RECT 242.665 47.365 248.850 47.505 ;
        RECT 242.665 47.305 242.985 47.365 ;
        RECT 244.960 47.320 245.610 47.365 ;
        RECT 248.560 47.320 248.850 47.365 ;
        RECT 244.965 47.305 245.285 47.320 ;
        RECT 226.565 47.025 231.855 47.165 ;
        RECT 238.525 47.165 238.845 47.225 ;
        RECT 250.115 47.165 250.255 48.340 ;
        RECT 254.625 47.985 254.945 48.245 ;
        RECT 255.175 48.185 255.315 48.385 ;
        RECT 255.510 48.385 260.810 48.525 ;
        RECT 255.510 48.340 255.800 48.385 ;
        RECT 257.400 48.340 257.690 48.385 ;
        RECT 260.520 48.340 260.810 48.385 ;
        RECT 281.420 48.525 281.710 48.570 ;
        RECT 284.540 48.525 284.830 48.570 ;
        RECT 286.430 48.525 286.720 48.570 ;
        RECT 281.420 48.385 286.720 48.525 ;
        RECT 281.420 48.340 281.710 48.385 ;
        RECT 284.540 48.340 284.830 48.385 ;
        RECT 286.430 48.340 286.720 48.385 ;
        RECT 288.630 48.525 288.920 48.570 ;
        RECT 290.520 48.525 290.810 48.570 ;
        RECT 293.640 48.525 293.930 48.570 ;
        RECT 288.630 48.385 293.930 48.525 ;
        RECT 288.630 48.340 288.920 48.385 ;
        RECT 290.520 48.340 290.810 48.385 ;
        RECT 293.640 48.340 293.930 48.385 ;
        RECT 256.005 48.185 256.325 48.245 ;
        RECT 255.175 48.045 256.325 48.185 ;
        RECT 256.005 47.985 256.325 48.045 ;
        RECT 256.465 48.185 256.785 48.245 ;
        RECT 263.365 48.185 263.685 48.245 ;
        RECT 256.465 48.045 262.215 48.185 ;
        RECT 256.465 47.985 256.785 48.045 ;
        RECT 255.105 47.845 255.395 47.890 ;
        RECT 256.940 47.845 257.230 47.890 ;
        RECT 260.520 47.845 260.810 47.890 ;
        RECT 255.105 47.705 260.810 47.845 ;
        RECT 255.105 47.660 255.395 47.705 ;
        RECT 256.940 47.660 257.230 47.705 ;
        RECT 260.520 47.660 260.810 47.705 ;
        RECT 256.020 47.505 256.310 47.550 ;
        RECT 257.385 47.505 257.705 47.565 ;
        RECT 261.600 47.550 261.890 47.865 ;
        RECT 262.075 47.845 262.215 48.045 ;
        RECT 263.365 48.045 269.805 48.185 ;
        RECT 263.365 47.985 263.685 48.045 ;
        RECT 266.600 47.845 266.890 47.890 ;
        RECT 262.075 47.705 266.890 47.845 ;
        RECT 266.600 47.660 266.890 47.705 ;
        RECT 267.505 47.645 267.825 47.905 ;
        RECT 267.985 47.660 268.275 47.890 ;
        RECT 269.665 47.845 269.805 48.045 ;
        RECT 277.165 47.985 277.485 48.245 ;
        RECT 287.285 48.185 287.605 48.245 ;
        RECT 287.760 48.185 288.050 48.230 ;
        RECT 289.585 48.185 289.905 48.245 ;
        RECT 287.285 48.045 289.905 48.185 ;
        RECT 287.285 47.985 287.605 48.045 ;
        RECT 287.760 48.000 288.050 48.045 ;
        RECT 289.585 47.985 289.905 48.045 ;
        RECT 296.500 48.185 296.790 48.230 ;
        RECT 297.880 48.185 298.170 48.230 ;
        RECT 296.500 48.045 298.170 48.185 ;
        RECT 296.500 48.000 296.790 48.045 ;
        RECT 297.880 48.000 298.170 48.045 ;
        RECT 270.040 47.845 270.330 47.890 ;
        RECT 269.665 47.705 270.330 47.845 ;
        RECT 270.040 47.660 270.330 47.705 ;
        RECT 258.300 47.505 258.950 47.550 ;
        RECT 261.600 47.505 262.190 47.550 ;
        RECT 256.020 47.365 257.705 47.505 ;
        RECT 256.020 47.320 256.310 47.365 ;
        RECT 257.385 47.305 257.705 47.365 ;
        RECT 257.935 47.365 262.190 47.505 ;
        RECT 238.525 47.025 250.255 47.165 ;
        RECT 251.865 47.165 252.185 47.225 ;
        RECT 257.935 47.165 258.075 47.365 ;
        RECT 258.300 47.320 258.950 47.365 ;
        RECT 261.900 47.320 262.190 47.365 ;
        RECT 266.125 47.505 266.445 47.565 ;
        RECT 268.055 47.505 268.195 47.660 ;
        RECT 266.125 47.365 268.195 47.505 ;
        RECT 266.125 47.305 266.445 47.365 ;
        RECT 268.900 47.320 269.190 47.550 ;
        RECT 269.345 47.505 269.665 47.565 ;
        RECT 277.625 47.505 277.945 47.565 ;
        RECT 280.340 47.550 280.630 47.865 ;
        RECT 281.420 47.845 281.710 47.890 ;
        RECT 285.000 47.845 285.290 47.890 ;
        RECT 286.835 47.845 287.125 47.890 ;
        RECT 281.420 47.705 287.125 47.845 ;
        RECT 281.420 47.660 281.710 47.705 ;
        RECT 285.000 47.660 285.290 47.705 ;
        RECT 286.835 47.660 287.125 47.705 ;
        RECT 288.225 47.845 288.515 47.890 ;
        RECT 290.060 47.845 290.350 47.890 ;
        RECT 293.640 47.845 293.930 47.890 ;
        RECT 288.225 47.705 293.930 47.845 ;
        RECT 288.225 47.660 288.515 47.705 ;
        RECT 290.060 47.660 290.350 47.705 ;
        RECT 293.640 47.660 293.930 47.705 ;
        RECT 283.605 47.550 283.925 47.565 ;
        RECT 269.345 47.365 277.945 47.505 ;
        RECT 259.685 47.165 260.005 47.225 ;
        RECT 251.865 47.025 260.005 47.165 ;
        RECT 220.585 46.965 220.905 47.025 ;
        RECT 226.565 46.965 226.885 47.025 ;
        RECT 238.525 46.965 238.845 47.025 ;
        RECT 251.865 46.965 252.185 47.025 ;
        RECT 259.685 46.965 260.005 47.025 ;
        RECT 263.365 46.965 263.685 47.225 ;
        RECT 268.975 47.165 269.115 47.320 ;
        RECT 269.345 47.305 269.665 47.365 ;
        RECT 277.625 47.305 277.945 47.365 ;
        RECT 280.040 47.505 280.630 47.550 ;
        RECT 283.280 47.505 283.930 47.550 ;
        RECT 280.040 47.365 283.930 47.505 ;
        RECT 280.040 47.320 280.330 47.365 ;
        RECT 283.280 47.320 283.930 47.365 ;
        RECT 283.605 47.305 283.925 47.320 ;
        RECT 285.905 47.305 286.225 47.565 ;
        RECT 289.140 47.505 289.430 47.550 ;
        RECT 290.505 47.505 290.825 47.565 ;
        RECT 294.720 47.550 295.010 47.865 ;
        RECT 289.140 47.365 290.825 47.505 ;
        RECT 289.140 47.320 289.430 47.365 ;
        RECT 290.505 47.305 290.825 47.365 ;
        RECT 291.420 47.505 292.070 47.550 ;
        RECT 294.720 47.505 295.310 47.550 ;
        RECT 297.405 47.505 297.725 47.565 ;
        RECT 303.385 47.505 303.705 47.565 ;
        RECT 291.420 47.365 303.705 47.505 ;
        RECT 291.420 47.320 292.070 47.365 ;
        RECT 295.020 47.320 295.310 47.365 ;
        RECT 297.405 47.305 297.725 47.365 ;
        RECT 303.385 47.305 303.705 47.365 ;
        RECT 274.405 47.165 274.725 47.225 ;
        RECT 268.975 47.025 274.725 47.165 ;
        RECT 274.405 46.965 274.725 47.025 ;
        RECT 298.785 47.165 299.105 47.225 ;
        RECT 301.100 47.165 301.390 47.210 ;
        RECT 298.785 47.025 301.390 47.165 ;
        RECT 298.785 46.965 299.105 47.025 ;
        RECT 301.100 46.980 301.390 47.025 ;
        RECT 162.095 46.345 311.135 46.825 ;
        RECT 176.425 46.145 176.745 46.205 ;
        RECT 180.580 46.145 180.870 46.190 ;
        RECT 183.325 46.145 183.645 46.205 ;
        RECT 204.945 46.145 205.265 46.205 ;
        RECT 233.005 46.145 233.325 46.205 ;
        RECT 242.665 46.145 242.985 46.205 ;
        RECT 176.425 46.005 179.875 46.145 ;
        RECT 176.425 45.945 176.745 46.005 ;
        RECT 175.500 45.805 176.150 45.850 ;
        RECT 179.100 45.805 179.390 45.850 ;
        RECT 175.500 45.665 179.390 45.805 ;
        RECT 179.735 45.805 179.875 46.005 ;
        RECT 180.580 46.005 183.645 46.145 ;
        RECT 180.580 45.960 180.870 46.005 ;
        RECT 183.325 45.945 183.645 46.005 ;
        RECT 183.875 46.005 197.355 46.145 ;
        RECT 183.875 45.805 184.015 46.005 ;
        RECT 179.735 45.665 184.015 45.805 ;
        RECT 192.980 45.805 193.630 45.850 ;
        RECT 196.580 45.805 196.870 45.850 ;
        RECT 192.980 45.665 196.870 45.805 ;
        RECT 197.215 45.805 197.355 46.005 ;
        RECT 204.945 46.005 233.325 46.145 ;
        RECT 204.945 45.945 205.265 46.005 ;
        RECT 233.005 45.945 233.325 46.005 ;
        RECT 239.535 46.005 242.985 46.145 ;
        RECT 208.625 45.805 208.945 45.865 ;
        RECT 197.215 45.665 208.945 45.805 ;
        RECT 175.500 45.620 176.150 45.665 ;
        RECT 178.800 45.620 179.390 45.665 ;
        RECT 192.980 45.620 193.630 45.665 ;
        RECT 196.280 45.620 196.870 45.665 ;
        RECT 172.305 45.465 172.595 45.510 ;
        RECT 174.140 45.465 174.430 45.510 ;
        RECT 177.720 45.465 178.010 45.510 ;
        RECT 172.305 45.325 178.010 45.465 ;
        RECT 172.305 45.280 172.595 45.325 ;
        RECT 174.140 45.280 174.430 45.325 ;
        RECT 177.720 45.280 178.010 45.325 ;
        RECT 178.800 45.465 179.090 45.620 ;
        RECT 184.245 45.465 184.565 45.525 ;
        RECT 178.800 45.325 184.565 45.465 ;
        RECT 178.800 45.305 179.090 45.325 ;
        RECT 184.245 45.265 184.565 45.325 ;
        RECT 189.305 45.265 189.625 45.525 ;
        RECT 189.785 45.465 190.075 45.510 ;
        RECT 191.620 45.465 191.910 45.510 ;
        RECT 195.200 45.465 195.490 45.510 ;
        RECT 189.785 45.325 195.490 45.465 ;
        RECT 189.785 45.280 190.075 45.325 ;
        RECT 191.620 45.280 191.910 45.325 ;
        RECT 195.200 45.280 195.490 45.325 ;
        RECT 196.280 45.465 196.570 45.620 ;
        RECT 208.625 45.605 208.945 45.665 ;
        RECT 220.120 45.805 220.770 45.850 ;
        RECT 223.720 45.805 224.010 45.850 ;
        RECT 226.105 45.805 226.425 45.865 ;
        RECT 220.120 45.665 226.425 45.805 ;
        RECT 220.120 45.620 220.770 45.665 ;
        RECT 223.420 45.620 224.010 45.665 ;
        RECT 197.125 45.465 197.445 45.525 ;
        RECT 196.280 45.325 197.445 45.465 ;
        RECT 196.280 45.305 196.570 45.325 ;
        RECT 197.125 45.265 197.445 45.325 ;
        RECT 203.120 45.465 203.410 45.510 ;
        RECT 205.420 45.465 205.710 45.510 ;
        RECT 203.120 45.325 205.710 45.465 ;
        RECT 203.120 45.280 203.410 45.325 ;
        RECT 205.420 45.280 205.710 45.325 ;
        RECT 211.385 45.265 211.705 45.525 ;
        RECT 216.445 45.265 216.765 45.525 ;
        RECT 216.925 45.465 217.215 45.510 ;
        RECT 218.760 45.465 219.050 45.510 ;
        RECT 222.340 45.465 222.630 45.510 ;
        RECT 216.925 45.325 222.630 45.465 ;
        RECT 216.925 45.280 217.215 45.325 ;
        RECT 218.760 45.280 219.050 45.325 ;
        RECT 222.340 45.280 222.630 45.325 ;
        RECT 223.420 45.305 223.710 45.620 ;
        RECT 226.105 45.605 226.425 45.665 ;
        RECT 233.920 45.805 234.570 45.850 ;
        RECT 237.520 45.805 237.810 45.850 ;
        RECT 233.920 45.665 237.810 45.805 ;
        RECT 233.920 45.620 234.570 45.665 ;
        RECT 237.220 45.620 237.810 45.665 ;
        RECT 227.025 45.265 227.345 45.525 ;
        RECT 227.945 45.265 228.265 45.525 ;
        RECT 228.880 45.280 229.170 45.510 ;
        RECT 166.305 45.125 166.625 45.185 ;
        RECT 171.840 45.125 172.130 45.170 ;
        RECT 166.305 44.985 172.130 45.125 ;
        RECT 166.305 44.925 166.625 44.985 ;
        RECT 171.840 44.940 172.130 44.985 ;
        RECT 173.220 45.125 173.510 45.170 ;
        RECT 173.220 44.985 181.715 45.125 ;
        RECT 173.220 44.940 173.510 44.985 ;
        RECT 171.915 44.445 172.055 44.940 ;
        RECT 181.575 44.830 181.715 44.985 ;
        RECT 183.785 44.925 184.105 45.185 ;
        RECT 184.705 45.125 185.025 45.185 ;
        RECT 190.700 45.125 190.990 45.170 ;
        RECT 197.585 45.125 197.905 45.185 ;
        RECT 184.705 44.985 197.905 45.125 ;
        RECT 184.705 44.925 185.025 44.985 ;
        RECT 190.700 44.940 190.990 44.985 ;
        RECT 197.585 44.925 197.905 44.985 ;
        RECT 199.900 44.940 200.190 45.170 ;
        RECT 172.710 44.785 173.000 44.830 ;
        RECT 174.600 44.785 174.890 44.830 ;
        RECT 177.720 44.785 178.010 44.830 ;
        RECT 172.710 44.645 178.010 44.785 ;
        RECT 172.710 44.600 173.000 44.645 ;
        RECT 174.600 44.600 174.890 44.645 ;
        RECT 177.720 44.600 178.010 44.645 ;
        RECT 181.500 44.600 181.790 44.830 ;
        RECT 190.190 44.785 190.480 44.830 ;
        RECT 192.080 44.785 192.370 44.830 ;
        RECT 195.200 44.785 195.490 44.830 ;
        RECT 199.975 44.785 200.115 44.940 ;
        RECT 205.865 44.925 206.185 45.185 ;
        RECT 206.800 45.125 207.090 45.170 ;
        RECT 210.480 45.125 210.770 45.170 ;
        RECT 206.800 44.985 210.770 45.125 ;
        RECT 206.800 44.940 207.090 44.985 ;
        RECT 210.480 44.940 210.770 44.985 ;
        RECT 210.940 45.125 211.230 45.170 ;
        RECT 214.605 45.125 214.925 45.185 ;
        RECT 210.940 44.985 214.925 45.125 ;
        RECT 210.940 44.940 211.230 44.985 ;
        RECT 190.190 44.645 195.490 44.785 ;
        RECT 190.190 44.600 190.480 44.645 ;
        RECT 192.080 44.600 192.370 44.645 ;
        RECT 195.200 44.600 195.490 44.645 ;
        RECT 197.675 44.645 200.115 44.785 ;
        RECT 175.505 44.445 175.825 44.505 ;
        RECT 171.915 44.305 175.825 44.445 ;
        RECT 175.505 44.245 175.825 44.305 ;
        RECT 188.385 44.445 188.705 44.505 ;
        RECT 197.675 44.445 197.815 44.645 ;
        RECT 188.385 44.305 197.815 44.445 ;
        RECT 188.385 44.245 188.705 44.305 ;
        RECT 198.045 44.245 198.365 44.505 ;
        RECT 199.975 44.445 200.115 44.645 ;
        RECT 202.645 44.785 202.965 44.845 ;
        RECT 203.580 44.785 203.870 44.830 ;
        RECT 202.645 44.645 203.870 44.785 ;
        RECT 210.555 44.785 210.695 44.940 ;
        RECT 214.605 44.925 214.925 44.985 ;
        RECT 217.825 44.925 218.145 45.185 ;
        RECT 225.185 44.925 225.505 45.185 ;
        RECT 228.405 44.925 228.725 45.185 ;
        RECT 212.765 44.785 213.085 44.845 ;
        RECT 210.555 44.645 213.085 44.785 ;
        RECT 202.645 44.585 202.965 44.645 ;
        RECT 203.580 44.600 203.870 44.645 ;
        RECT 212.765 44.585 213.085 44.645 ;
        RECT 217.330 44.785 217.620 44.830 ;
        RECT 219.220 44.785 219.510 44.830 ;
        RECT 222.340 44.785 222.630 44.830 ;
        RECT 217.330 44.645 222.630 44.785 ;
        RECT 217.330 44.600 217.620 44.645 ;
        RECT 219.220 44.600 219.510 44.645 ;
        RECT 222.340 44.600 222.630 44.645 ;
        RECT 210.005 44.445 210.325 44.505 ;
        RECT 199.975 44.305 210.325 44.445 ;
        RECT 210.005 44.245 210.325 44.305 ;
        RECT 213.225 44.245 213.545 44.505 ;
        RECT 226.105 44.245 226.425 44.505 ;
        RECT 228.955 44.445 229.095 45.280 ;
        RECT 229.785 45.265 230.105 45.525 ;
        RECT 230.725 45.465 231.015 45.510 ;
        RECT 232.560 45.465 232.850 45.510 ;
        RECT 236.140 45.465 236.430 45.510 ;
        RECT 230.725 45.325 236.430 45.465 ;
        RECT 230.725 45.280 231.015 45.325 ;
        RECT 232.560 45.280 232.850 45.325 ;
        RECT 236.140 45.280 236.430 45.325 ;
        RECT 237.220 45.465 237.510 45.620 ;
        RECT 239.535 45.465 239.675 46.005 ;
        RECT 242.665 45.945 242.985 46.005 ;
        RECT 243.600 46.145 243.890 46.190 ;
        RECT 244.505 46.145 244.825 46.205 ;
        RECT 243.600 46.005 244.825 46.145 ;
        RECT 243.600 45.960 243.890 46.005 ;
        RECT 244.505 45.945 244.825 46.005 ;
        RECT 252.785 46.145 253.105 46.205 ;
        RECT 264.745 46.145 265.065 46.205 ;
        RECT 252.785 46.005 265.895 46.145 ;
        RECT 252.785 45.945 253.105 46.005 ;
        RECT 264.745 45.945 265.065 46.005 ;
        RECT 240.365 45.805 240.685 45.865 ;
        RECT 244.965 45.805 245.285 45.865 ;
        RECT 251.865 45.850 252.185 45.865 ;
        RECT 251.860 45.805 252.510 45.850 ;
        RECT 255.460 45.805 255.750 45.850 ;
        RECT 240.365 45.665 244.735 45.805 ;
        RECT 240.365 45.605 240.685 45.665 ;
        RECT 237.220 45.325 239.675 45.465 ;
        RECT 237.220 45.305 237.510 45.325 ;
        RECT 239.905 45.265 240.225 45.525 ;
        RECT 240.840 45.465 241.130 45.510 ;
        RECT 242.205 45.465 242.525 45.525 ;
        RECT 240.840 45.325 242.525 45.465 ;
        RECT 240.840 45.280 241.130 45.325 ;
        RECT 230.245 44.925 230.565 45.185 ;
        RECT 231.625 44.925 231.945 45.185 ;
        RECT 231.130 44.785 231.420 44.830 ;
        RECT 233.020 44.785 233.310 44.830 ;
        RECT 236.140 44.785 236.430 44.830 ;
        RECT 240.915 44.785 241.055 45.280 ;
        RECT 242.205 45.265 242.525 45.325 ;
        RECT 242.665 45.265 242.985 45.525 ;
        RECT 244.595 45.465 244.735 45.665 ;
        RECT 244.965 45.665 255.750 45.805 ;
        RECT 244.965 45.605 245.285 45.665 ;
        RECT 251.860 45.620 252.510 45.665 ;
        RECT 255.160 45.620 255.750 45.665 ;
        RECT 251.865 45.605 252.185 45.620 ;
        RECT 248.200 45.465 248.490 45.510 ;
        RECT 244.595 45.325 248.490 45.465 ;
        RECT 248.200 45.280 248.490 45.325 ;
        RECT 248.665 45.465 248.955 45.510 ;
        RECT 250.500 45.465 250.790 45.510 ;
        RECT 254.080 45.465 254.370 45.510 ;
        RECT 248.665 45.325 254.370 45.465 ;
        RECT 248.665 45.280 248.955 45.325 ;
        RECT 250.500 45.280 250.790 45.325 ;
        RECT 254.080 45.280 254.370 45.325 ;
        RECT 255.160 45.305 255.450 45.620 ;
        RECT 257.385 45.605 257.705 45.865 ;
        RECT 262.460 45.805 262.750 45.850 ;
        RECT 265.205 45.805 265.525 45.865 ;
        RECT 265.755 45.850 265.895 46.005 ;
        RECT 267.505 45.945 267.825 46.205 ;
        RECT 268.425 46.145 268.745 46.205 ;
        RECT 274.405 46.145 274.725 46.205 ;
        RECT 280.400 46.145 280.690 46.190 ;
        RECT 268.425 46.005 270.495 46.145 ;
        RECT 268.425 45.945 268.745 46.005 ;
        RECT 262.460 45.665 265.525 45.805 ;
        RECT 262.460 45.620 262.750 45.665 ;
        RECT 265.205 45.605 265.525 45.665 ;
        RECT 265.680 45.620 265.970 45.850 ;
        RECT 266.830 45.635 267.120 45.680 ;
        RECT 267.595 45.665 269.575 45.805 ;
        RECT 267.595 45.635 267.735 45.665 ;
        RECT 260.145 45.265 260.465 45.525 ;
        RECT 262.000 45.465 262.290 45.510 ;
        RECT 260.695 45.325 262.290 45.465 ;
        RECT 241.285 44.925 241.605 45.185 ;
        RECT 241.745 44.925 242.065 45.185 ;
        RECT 245.885 45.125 246.205 45.185 ;
        RECT 246.820 45.125 247.110 45.170 ;
        RECT 245.885 44.985 247.110 45.125 ;
        RECT 245.885 44.925 246.205 44.985 ;
        RECT 246.820 44.940 247.110 44.985 ;
        RECT 249.580 45.125 249.870 45.170 ;
        RECT 251.865 45.125 252.185 45.185 ;
        RECT 249.580 44.985 252.185 45.125 ;
        RECT 249.580 44.940 249.870 44.985 ;
        RECT 251.865 44.925 252.185 44.985 ;
        RECT 256.465 45.125 256.785 45.185 ;
        RECT 256.940 45.125 257.230 45.170 ;
        RECT 256.465 44.985 257.230 45.125 ;
        RECT 256.465 44.925 256.785 44.985 ;
        RECT 256.940 44.940 257.230 44.985 ;
        RECT 243.585 44.785 243.905 44.845 ;
        RECT 231.130 44.645 236.430 44.785 ;
        RECT 231.130 44.600 231.420 44.645 ;
        RECT 233.020 44.600 233.310 44.645 ;
        RECT 236.140 44.600 236.430 44.645 ;
        RECT 238.615 44.645 241.055 44.785 ;
        RECT 241.835 44.645 243.905 44.785 ;
        RECT 237.605 44.445 237.925 44.505 ;
        RECT 238.615 44.445 238.755 44.645 ;
        RECT 228.955 44.305 238.755 44.445 ;
        RECT 239.000 44.445 239.290 44.490 ;
        RECT 241.835 44.445 241.975 44.645 ;
        RECT 243.585 44.585 243.905 44.645 ;
        RECT 249.070 44.785 249.360 44.830 ;
        RECT 250.960 44.785 251.250 44.830 ;
        RECT 254.080 44.785 254.370 44.830 ;
        RECT 249.070 44.645 254.370 44.785 ;
        RECT 249.070 44.600 249.360 44.645 ;
        RECT 250.960 44.600 251.250 44.645 ;
        RECT 254.080 44.600 254.370 44.645 ;
        RECT 255.545 44.785 255.865 44.845 ;
        RECT 260.695 44.785 260.835 45.325 ;
        RECT 262.000 45.280 262.290 45.325 ;
        RECT 262.920 45.280 263.210 45.510 ;
        RECT 263.840 45.465 264.130 45.510 ;
        RECT 266.125 45.465 266.445 45.525 ;
        RECT 263.840 45.325 266.445 45.465 ;
        RECT 266.830 45.495 267.735 45.635 ;
        RECT 266.830 45.450 267.120 45.495 ;
        RECT 263.840 45.280 264.130 45.325 ;
        RECT 262.995 45.125 263.135 45.280 ;
        RECT 266.125 45.265 266.445 45.325 ;
        RECT 267.965 45.265 268.285 45.525 ;
        RECT 268.885 45.265 269.205 45.525 ;
        RECT 269.435 45.465 269.575 45.665 ;
        RECT 269.820 45.465 270.110 45.510 ;
        RECT 269.435 45.325 270.110 45.465 ;
        RECT 270.355 45.465 270.495 46.005 ;
        RECT 274.405 46.005 280.690 46.145 ;
        RECT 274.405 45.945 274.725 46.005 ;
        RECT 280.400 45.960 280.690 46.005 ;
        RECT 285.905 45.945 286.225 46.205 ;
        RECT 278.545 45.805 278.865 45.865 ;
        RECT 279.940 45.805 280.230 45.850 ;
        RECT 278.545 45.665 280.230 45.805 ;
        RECT 278.545 45.605 278.865 45.665 ;
        RECT 279.940 45.620 280.230 45.665 ;
        RECT 292.920 45.805 293.210 45.850 ;
        RECT 296.160 45.805 296.810 45.850 ;
        RECT 297.405 45.805 297.725 45.865 ;
        RECT 292.920 45.665 297.725 45.805 ;
        RECT 292.920 45.620 293.510 45.665 ;
        RECT 296.160 45.620 296.810 45.665 ;
        RECT 270.740 45.465 271.030 45.510 ;
        RECT 272.105 45.465 272.425 45.525 ;
        RECT 270.355 45.325 271.030 45.465 ;
        RECT 269.820 45.280 270.110 45.325 ;
        RECT 270.740 45.280 271.030 45.325 ;
        RECT 271.275 45.325 272.425 45.465 ;
        RECT 264.285 45.125 264.605 45.185 ;
        RECT 262.995 44.985 264.605 45.125 ;
        RECT 269.895 45.125 270.035 45.280 ;
        RECT 271.275 45.125 271.415 45.325 ;
        RECT 272.105 45.265 272.425 45.325 ;
        RECT 293.220 45.305 293.510 45.620 ;
        RECT 297.405 45.605 297.725 45.665 ;
        RECT 298.785 45.605 299.105 45.865 ;
        RECT 294.300 45.465 294.590 45.510 ;
        RECT 297.880 45.465 298.170 45.510 ;
        RECT 299.715 45.465 300.005 45.510 ;
        RECT 294.300 45.325 300.005 45.465 ;
        RECT 294.300 45.280 294.590 45.325 ;
        RECT 297.880 45.280 298.170 45.325 ;
        RECT 299.715 45.280 300.005 45.325 ;
        RECT 279.020 45.125 279.310 45.170 ;
        RECT 269.895 44.985 271.415 45.125 ;
        RECT 271.735 44.985 279.310 45.125 ;
        RECT 264.285 44.925 264.605 44.985 ;
        RECT 255.545 44.645 260.835 44.785 ;
        RECT 261.080 44.785 261.370 44.830 ;
        RECT 270.725 44.785 271.045 44.845 ;
        RECT 261.080 44.645 271.045 44.785 ;
        RECT 255.545 44.585 255.865 44.645 ;
        RECT 261.080 44.600 261.370 44.645 ;
        RECT 270.725 44.585 271.045 44.645 ;
        RECT 271.735 44.505 271.875 44.985 ;
        RECT 279.020 44.940 279.310 44.985 ;
        RECT 282.700 44.940 282.990 45.170 ;
        RECT 300.180 45.125 300.470 45.170 ;
        RECT 305.685 45.125 306.005 45.185 ;
        RECT 300.180 44.985 306.005 45.125 ;
        RECT 300.180 44.940 300.470 44.985 ;
        RECT 282.240 44.785 282.530 44.830 ;
        RECT 282.775 44.785 282.915 44.940 ;
        RECT 305.685 44.925 306.005 44.985 ;
        RECT 282.240 44.645 282.915 44.785 ;
        RECT 294.300 44.785 294.590 44.830 ;
        RECT 297.420 44.785 297.710 44.830 ;
        RECT 299.310 44.785 299.600 44.830 ;
        RECT 294.300 44.645 299.600 44.785 ;
        RECT 282.240 44.600 282.530 44.645 ;
        RECT 294.300 44.600 294.590 44.645 ;
        RECT 297.420 44.600 297.710 44.645 ;
        RECT 299.310 44.600 299.600 44.645 ;
        RECT 239.000 44.305 241.975 44.445 ;
        RECT 242.665 44.445 242.985 44.505 ;
        RECT 244.060 44.445 244.350 44.490 ;
        RECT 242.665 44.305 244.350 44.445 ;
        RECT 237.605 44.245 237.925 44.305 ;
        RECT 239.000 44.260 239.290 44.305 ;
        RECT 242.665 44.245 242.985 44.305 ;
        RECT 244.060 44.260 244.350 44.305 ;
        RECT 263.365 44.445 263.685 44.505 ;
        RECT 266.600 44.445 266.890 44.490 ;
        RECT 263.365 44.305 266.890 44.445 ;
        RECT 263.365 44.245 263.685 44.305 ;
        RECT 266.600 44.260 266.890 44.305 ;
        RECT 271.645 44.245 271.965 44.505 ;
        RECT 289.125 44.445 289.445 44.505 ;
        RECT 291.440 44.445 291.730 44.490 ;
        RECT 289.125 44.305 291.730 44.445 ;
        RECT 289.125 44.245 289.445 44.305 ;
        RECT 291.440 44.260 291.730 44.305 ;
        RECT 162.095 43.625 311.135 44.105 ;
        RECT 174.600 43.425 174.890 43.470 ;
        RECT 180.105 43.425 180.425 43.485 ;
        RECT 174.600 43.285 180.425 43.425 ;
        RECT 174.600 43.240 174.890 43.285 ;
        RECT 180.105 43.225 180.425 43.285 ;
        RECT 182.865 43.425 183.185 43.485 ;
        RECT 184.260 43.425 184.550 43.470 ;
        RECT 182.865 43.285 184.550 43.425 ;
        RECT 182.865 43.225 183.185 43.285 ;
        RECT 184.260 43.240 184.550 43.285 ;
        RECT 197.585 43.425 197.905 43.485 ;
        RECT 212.765 43.425 213.085 43.485 ;
        RECT 197.585 43.285 213.085 43.425 ;
        RECT 197.585 43.225 197.905 43.285 ;
        RECT 212.765 43.225 213.085 43.285 ;
        RECT 213.225 43.425 213.545 43.485 ;
        RECT 214.985 43.425 215.275 43.470 ;
        RECT 213.225 43.285 215.275 43.425 ;
        RECT 213.225 43.225 213.545 43.285 ;
        RECT 214.985 43.240 215.275 43.285 ;
        RECT 222.440 43.425 222.730 43.470 ;
        RECT 222.885 43.425 223.205 43.485 ;
        RECT 222.440 43.285 223.205 43.425 ;
        RECT 222.440 43.240 222.730 43.285 ;
        RECT 222.885 43.225 223.205 43.285 ;
        RECT 226.120 43.425 226.410 43.470 ;
        RECT 226.565 43.425 226.885 43.485 ;
        RECT 226.120 43.285 226.885 43.425 ;
        RECT 226.120 43.240 226.410 43.285 ;
        RECT 226.565 43.225 226.885 43.285 ;
        RECT 227.485 43.225 227.805 43.485 ;
        RECT 228.405 43.425 228.725 43.485 ;
        RECT 238.985 43.425 239.305 43.485 ;
        RECT 239.460 43.425 239.750 43.470 ;
        RECT 228.405 43.285 236.915 43.425 ;
        RECT 228.405 43.225 228.725 43.285 ;
        RECT 166.730 43.085 167.020 43.130 ;
        RECT 168.620 43.085 168.910 43.130 ;
        RECT 171.740 43.085 172.030 43.130 ;
        RECT 166.730 42.945 172.030 43.085 ;
        RECT 166.730 42.900 167.020 42.945 ;
        RECT 168.620 42.900 168.910 42.945 ;
        RECT 171.740 42.900 172.030 42.945 ;
        RECT 176.390 43.085 176.680 43.130 ;
        RECT 178.280 43.085 178.570 43.130 ;
        RECT 181.400 43.085 181.690 43.130 ;
        RECT 176.390 42.945 181.690 43.085 ;
        RECT 176.390 42.900 176.680 42.945 ;
        RECT 178.280 42.900 178.570 42.945 ;
        RECT 181.400 42.900 181.690 42.945 ;
        RECT 185.590 43.085 185.880 43.130 ;
        RECT 187.480 43.085 187.770 43.130 ;
        RECT 190.600 43.085 190.890 43.130 ;
        RECT 185.590 42.945 190.890 43.085 ;
        RECT 185.590 42.900 185.880 42.945 ;
        RECT 187.480 42.900 187.770 42.945 ;
        RECT 190.600 42.900 190.890 42.945 ;
        RECT 175.505 42.745 175.825 42.805 ;
        RECT 184.720 42.745 185.010 42.790 ;
        RECT 189.305 42.745 189.625 42.805 ;
        RECT 193.905 42.745 194.225 42.805 ;
        RECT 197.125 42.745 197.445 42.805 ;
        RECT 197.675 42.790 197.815 43.225 ;
        RECT 202.150 43.085 202.440 43.130 ;
        RECT 204.040 43.085 204.330 43.130 ;
        RECT 207.160 43.085 207.450 43.130 ;
        RECT 202.150 42.945 207.450 43.085 ;
        RECT 202.150 42.900 202.440 42.945 ;
        RECT 204.040 42.900 204.330 42.945 ;
        RECT 207.160 42.900 207.450 42.945 ;
        RECT 210.005 42.885 210.325 43.145 ;
        RECT 211.845 42.885 212.165 43.145 ;
        RECT 214.570 43.085 214.860 43.130 ;
        RECT 216.460 43.085 216.750 43.130 ;
        RECT 219.580 43.085 219.870 43.130 ;
        RECT 214.570 42.945 219.870 43.085 ;
        RECT 214.570 42.900 214.860 42.945 ;
        RECT 216.460 42.900 216.750 42.945 ;
        RECT 219.580 42.900 219.870 42.945 ;
        RECT 231.130 43.085 231.420 43.130 ;
        RECT 233.020 43.085 233.310 43.130 ;
        RECT 236.140 43.085 236.430 43.130 ;
        RECT 231.130 42.945 236.430 43.085 ;
        RECT 236.775 43.085 236.915 43.285 ;
        RECT 238.985 43.285 239.750 43.425 ;
        RECT 238.985 43.225 239.305 43.285 ;
        RECT 239.460 43.240 239.750 43.285 ;
        RECT 251.865 43.225 252.185 43.485 ;
        RECT 256.925 43.425 257.245 43.485 ;
        RECT 257.860 43.425 258.150 43.470 ;
        RECT 269.345 43.425 269.665 43.485 ;
        RECT 256.925 43.285 258.150 43.425 ;
        RECT 256.925 43.225 257.245 43.285 ;
        RECT 257.860 43.240 258.150 43.285 ;
        RECT 266.675 43.285 269.665 43.425 ;
        RECT 243.600 43.085 243.890 43.130 ;
        RECT 236.775 42.945 243.890 43.085 ;
        RECT 231.130 42.900 231.420 42.945 ;
        RECT 233.020 42.900 233.310 42.945 ;
        RECT 236.140 42.900 236.430 42.945 ;
        RECT 243.600 42.900 243.890 42.945 ;
        RECT 255.085 43.085 255.405 43.145 ;
        RECT 263.825 43.085 264.145 43.145 ;
        RECT 255.085 42.945 264.145 43.085 ;
        RECT 255.085 42.885 255.405 42.945 ;
        RECT 263.825 42.885 264.145 42.945 ;
        RECT 264.745 42.885 265.065 43.145 ;
        RECT 175.505 42.605 189.625 42.745 ;
        RECT 175.505 42.545 175.825 42.605 ;
        RECT 184.720 42.560 185.010 42.605 ;
        RECT 189.305 42.545 189.625 42.605 ;
        RECT 191.695 42.605 197.445 42.745 ;
        RECT 165.845 42.205 166.165 42.465 ;
        RECT 166.325 42.405 166.615 42.450 ;
        RECT 168.160 42.405 168.450 42.450 ;
        RECT 171.740 42.405 172.030 42.450 ;
        RECT 166.325 42.265 172.030 42.405 ;
        RECT 166.325 42.220 166.615 42.265 ;
        RECT 168.160 42.220 168.450 42.265 ;
        RECT 171.740 42.220 172.030 42.265 ;
        RECT 167.225 41.865 167.545 42.125 ;
        RECT 172.820 42.110 173.110 42.425 ;
        RECT 175.985 42.405 176.275 42.450 ;
        RECT 177.820 42.405 178.110 42.450 ;
        RECT 181.400 42.405 181.690 42.450 ;
        RECT 175.985 42.265 181.690 42.405 ;
        RECT 175.985 42.220 176.275 42.265 ;
        RECT 177.820 42.220 178.110 42.265 ;
        RECT 181.400 42.220 181.690 42.265 ;
        RECT 169.520 42.065 170.170 42.110 ;
        RECT 172.820 42.065 173.410 42.110 ;
        RECT 169.520 41.925 173.895 42.065 ;
        RECT 169.520 41.880 170.170 41.925 ;
        RECT 173.120 41.880 173.410 41.925 ;
        RECT 172.285 41.725 172.605 41.785 ;
        RECT 173.755 41.725 173.895 41.925 ;
        RECT 176.885 41.865 177.205 42.125 ;
        RECT 182.480 42.110 182.770 42.425 ;
        RECT 185.185 42.405 185.475 42.450 ;
        RECT 187.020 42.405 187.310 42.450 ;
        RECT 190.600 42.405 190.890 42.450 ;
        RECT 191.695 42.425 191.835 42.605 ;
        RECT 193.905 42.545 194.225 42.605 ;
        RECT 197.125 42.545 197.445 42.605 ;
        RECT 197.600 42.560 197.890 42.790 ;
        RECT 202.645 42.545 202.965 42.805 ;
        RECT 213.700 42.745 213.990 42.790 ;
        RECT 218.745 42.745 219.065 42.805 ;
        RECT 213.700 42.605 219.065 42.745 ;
        RECT 213.700 42.560 213.990 42.605 ;
        RECT 218.745 42.545 219.065 42.605 ;
        RECT 223.360 42.745 223.650 42.790 ;
        RECT 226.105 42.745 226.425 42.805 ;
        RECT 223.360 42.605 226.425 42.745 ;
        RECT 223.360 42.560 223.650 42.605 ;
        RECT 226.105 42.545 226.425 42.605 ;
        RECT 231.640 42.745 231.930 42.790 ;
        RECT 235.305 42.745 235.625 42.805 ;
        RECT 231.640 42.605 235.625 42.745 ;
        RECT 231.640 42.560 231.930 42.605 ;
        RECT 235.305 42.545 235.625 42.605 ;
        RECT 236.685 42.745 237.005 42.805 ;
        RECT 241.300 42.745 241.590 42.790 ;
        RECT 236.685 42.605 241.590 42.745 ;
        RECT 236.685 42.545 237.005 42.605 ;
        RECT 241.300 42.560 241.590 42.605 ;
        RECT 241.760 42.745 242.050 42.790 ;
        RECT 242.665 42.745 242.985 42.805 ;
        RECT 241.760 42.605 242.985 42.745 ;
        RECT 241.760 42.560 242.050 42.605 ;
        RECT 242.665 42.545 242.985 42.605 ;
        RECT 246.805 42.745 247.125 42.805 ;
        RECT 248.660 42.745 248.950 42.790 ;
        RECT 262.905 42.745 263.225 42.805 ;
        RECT 246.805 42.605 248.950 42.745 ;
        RECT 246.805 42.545 247.125 42.605 ;
        RECT 248.660 42.560 248.950 42.605 ;
        RECT 258.400 42.605 263.225 42.745 ;
        RECT 185.185 42.265 190.890 42.405 ;
        RECT 185.185 42.220 185.475 42.265 ;
        RECT 187.020 42.220 187.310 42.265 ;
        RECT 190.600 42.220 190.890 42.265 ;
        RECT 179.180 42.065 179.830 42.110 ;
        RECT 182.480 42.065 183.070 42.110 ;
        RECT 184.245 42.065 184.565 42.125 ;
        RECT 179.180 41.925 184.565 42.065 ;
        RECT 179.180 41.880 179.830 41.925 ;
        RECT 182.780 41.880 183.070 41.925 ;
        RECT 183.415 41.725 183.555 41.925 ;
        RECT 184.245 41.865 184.565 41.925 ;
        RECT 186.085 41.865 186.405 42.125 ;
        RECT 191.680 42.110 191.970 42.425 ;
        RECT 195.745 42.405 196.065 42.465 ;
        RECT 201.280 42.405 201.570 42.450 ;
        RECT 195.745 42.265 201.570 42.405 ;
        RECT 195.745 42.205 196.065 42.265 ;
        RECT 201.280 42.220 201.570 42.265 ;
        RECT 201.745 42.405 202.035 42.450 ;
        RECT 203.580 42.405 203.870 42.450 ;
        RECT 207.160 42.405 207.450 42.450 ;
        RECT 201.745 42.265 207.450 42.405 ;
        RECT 201.745 42.220 202.035 42.265 ;
        RECT 203.580 42.220 203.870 42.265 ;
        RECT 207.160 42.220 207.450 42.265 ;
        RECT 208.165 42.425 208.485 42.465 ;
        RECT 208.165 42.405 208.530 42.425 ;
        RECT 214.165 42.405 214.455 42.450 ;
        RECT 216.000 42.405 216.290 42.450 ;
        RECT 219.580 42.405 219.870 42.450 ;
        RECT 208.165 42.265 212.535 42.405 ;
        RECT 208.165 42.205 208.530 42.265 ;
        RECT 188.380 42.065 189.030 42.110 ;
        RECT 191.680 42.065 192.270 42.110 ;
        RECT 188.380 41.925 192.270 42.065 ;
        RECT 188.380 41.880 189.030 41.925 ;
        RECT 191.980 41.880 192.270 41.925 ;
        RECT 192.525 42.065 192.845 42.125 ;
        RECT 208.240 42.110 208.530 42.205 ;
        RECT 196.680 42.065 196.970 42.110 ;
        RECT 192.525 41.925 196.970 42.065 ;
        RECT 192.525 41.865 192.845 41.925 ;
        RECT 196.680 41.880 196.970 41.925 ;
        RECT 204.940 42.065 205.590 42.110 ;
        RECT 208.240 42.065 208.830 42.110 ;
        RECT 210.480 42.065 210.770 42.110 ;
        RECT 204.940 41.925 208.830 42.065 ;
        RECT 204.940 41.880 205.590 41.925 ;
        RECT 208.540 41.880 208.830 41.925 ;
        RECT 209.175 41.925 210.770 42.065 ;
        RECT 212.395 42.065 212.535 42.265 ;
        RECT 214.165 42.265 219.870 42.405 ;
        RECT 214.165 42.220 214.455 42.265 ;
        RECT 216.000 42.220 216.290 42.265 ;
        RECT 219.580 42.220 219.870 42.265 ;
        RECT 217.365 42.110 217.685 42.125 ;
        RECT 217.825 42.110 218.145 42.125 ;
        RECT 217.360 42.065 218.145 42.110 ;
        RECT 220.660 42.110 220.950 42.425 ;
        RECT 222.885 42.405 223.205 42.465 ;
        RECT 227.025 42.405 227.345 42.465 ;
        RECT 230.245 42.405 230.565 42.465 ;
        RECT 222.885 42.265 226.795 42.405 ;
        RECT 222.885 42.205 223.205 42.265 ;
        RECT 220.660 42.065 221.250 42.110 ;
        RECT 212.395 41.925 221.250 42.065 ;
        RECT 226.655 42.065 226.795 42.265 ;
        RECT 227.025 42.265 230.565 42.405 ;
        RECT 227.025 42.205 227.345 42.265 ;
        RECT 230.245 42.205 230.565 42.265 ;
        RECT 230.725 42.405 231.015 42.450 ;
        RECT 232.560 42.405 232.850 42.450 ;
        RECT 236.140 42.405 236.430 42.450 ;
        RECT 230.725 42.265 236.430 42.405 ;
        RECT 230.725 42.220 231.015 42.265 ;
        RECT 232.560 42.220 232.850 42.265 ;
        RECT 236.140 42.220 236.430 42.265 ;
        RECT 237.220 42.110 237.510 42.425 ;
        RECT 240.365 42.205 240.685 42.465 ;
        RECT 242.205 42.205 242.525 42.465 ;
        RECT 243.125 42.205 243.445 42.465 ;
        RECT 246.360 42.220 246.650 42.450 ;
        RECT 228.880 42.065 229.170 42.110 ;
        RECT 226.655 41.925 229.170 42.065 ;
        RECT 172.285 41.585 183.555 41.725 ;
        RECT 190.225 41.725 190.545 41.785 ;
        RECT 192.985 41.725 193.305 41.785 ;
        RECT 193.460 41.725 193.750 41.770 ;
        RECT 190.225 41.585 193.750 41.725 ;
        RECT 172.285 41.525 172.605 41.585 ;
        RECT 190.225 41.525 190.545 41.585 ;
        RECT 192.985 41.525 193.305 41.585 ;
        RECT 193.460 41.540 193.750 41.585 ;
        RECT 194.365 41.525 194.685 41.785 ;
        RECT 196.205 41.525 196.525 41.785 ;
        RECT 198.045 41.725 198.365 41.785 ;
        RECT 209.175 41.725 209.315 41.925 ;
        RECT 210.480 41.880 210.770 41.925 ;
        RECT 217.360 41.880 218.145 41.925 ;
        RECT 220.960 41.880 221.250 41.925 ;
        RECT 228.880 41.880 229.170 41.925 ;
        RECT 233.920 42.065 234.570 42.110 ;
        RECT 237.220 42.065 237.810 42.110 ;
        RECT 238.065 42.065 238.385 42.125 ;
        RECT 246.435 42.065 246.575 42.220 ;
        RECT 233.920 41.925 238.385 42.065 ;
        RECT 233.920 41.880 234.570 41.925 ;
        RECT 237.520 41.880 237.810 41.925 ;
        RECT 217.365 41.865 217.685 41.880 ;
        RECT 217.825 41.865 218.145 41.880 ;
        RECT 238.065 41.865 238.385 41.925 ;
        RECT 239.535 41.925 246.575 42.065 ;
        RECT 249.105 42.065 249.425 42.125 ;
        RECT 253.260 42.065 253.550 42.110 ;
        RECT 249.105 41.925 253.550 42.065 ;
        RECT 239.535 41.785 239.675 41.925 ;
        RECT 249.105 41.865 249.425 41.925 ;
        RECT 253.260 41.880 253.550 41.925 ;
        RECT 253.705 42.065 254.025 42.125 ;
        RECT 258.400 42.065 258.540 42.605 ;
        RECT 262.905 42.545 263.225 42.605 ;
        RECT 258.780 42.405 259.070 42.450 ;
        RECT 263.365 42.405 263.685 42.465 ;
        RECT 258.780 42.265 263.685 42.405 ;
        RECT 258.780 42.220 259.070 42.265 ;
        RECT 263.365 42.205 263.685 42.265 ;
        RECT 264.300 42.405 264.590 42.450 ;
        RECT 265.205 42.405 265.525 42.465 ;
        RECT 266.675 42.405 266.815 43.285 ;
        RECT 269.345 43.225 269.665 43.285 ;
        RECT 272.105 43.425 272.425 43.485 ;
        RECT 276.720 43.425 277.010 43.470 ;
        RECT 272.105 43.285 277.010 43.425 ;
        RECT 272.105 43.225 272.425 43.285 ;
        RECT 276.720 43.240 277.010 43.285 ;
        RECT 267.930 43.085 268.220 43.130 ;
        RECT 269.820 43.085 270.110 43.130 ;
        RECT 272.940 43.085 273.230 43.130 ;
        RECT 279.940 43.085 280.230 43.130 ;
        RECT 267.930 42.945 273.230 43.085 ;
        RECT 267.930 42.900 268.220 42.945 ;
        RECT 269.820 42.900 270.110 42.945 ;
        RECT 272.940 42.900 273.230 42.945 ;
        RECT 273.575 42.945 280.230 43.085 ;
        RECT 267.045 42.545 267.365 42.805 ;
        RECT 272.105 42.745 272.425 42.805 ;
        RECT 273.575 42.745 273.715 42.945 ;
        RECT 279.940 42.900 280.230 42.945 ;
        RECT 280.385 43.085 280.705 43.145 ;
        RECT 280.385 42.945 289.355 43.085 ;
        RECT 280.385 42.885 280.705 42.945 ;
        RECT 289.215 42.805 289.355 42.945 ;
        RECT 272.105 42.605 273.715 42.745 ;
        RECT 275.800 42.745 276.090 42.790 ;
        RECT 276.260 42.745 276.550 42.790 ;
        RECT 275.800 42.605 276.550 42.745 ;
        RECT 272.105 42.545 272.425 42.605 ;
        RECT 275.800 42.560 276.090 42.605 ;
        RECT 276.260 42.560 276.550 42.605 ;
        RECT 277.180 42.745 277.470 42.790 ;
        RECT 285.000 42.745 285.290 42.790 ;
        RECT 277.180 42.605 285.290 42.745 ;
        RECT 277.180 42.560 277.470 42.605 ;
        RECT 264.300 42.265 266.815 42.405 ;
        RECT 267.525 42.405 267.815 42.450 ;
        RECT 269.360 42.405 269.650 42.450 ;
        RECT 272.940 42.405 273.230 42.450 ;
        RECT 267.525 42.265 273.230 42.405 ;
        RECT 264.300 42.220 264.590 42.265 ;
        RECT 265.205 42.205 265.525 42.265 ;
        RECT 267.525 42.220 267.815 42.265 ;
        RECT 269.360 42.220 269.650 42.265 ;
        RECT 272.940 42.220 273.230 42.265 ;
        RECT 273.945 42.425 274.265 42.465 ;
        RECT 273.945 42.205 274.310 42.425 ;
        RECT 277.625 42.405 277.945 42.465 ;
        RECT 278.635 42.450 278.775 42.605 ;
        RECT 285.000 42.560 285.290 42.605 ;
        RECT 289.125 42.545 289.445 42.805 ;
        RECT 277.625 42.265 278.315 42.405 ;
        RECT 277.625 42.205 277.945 42.265 ;
        RECT 259.700 42.065 259.990 42.110 ;
        RECT 253.705 41.925 259.990 42.065 ;
        RECT 253.705 41.865 254.025 41.925 ;
        RECT 259.700 41.880 259.990 41.925 ;
        RECT 260.145 41.865 260.465 42.125 ;
        RECT 261.080 41.880 261.370 42.110 ;
        RECT 262.000 42.065 262.290 42.110 ;
        RECT 267.045 42.065 267.365 42.125 ;
        RECT 262.000 41.925 267.365 42.065 ;
        RECT 262.000 41.880 262.290 41.925 ;
        RECT 198.045 41.585 209.315 41.725 ;
        RECT 212.765 41.725 213.085 41.785 ;
        RECT 226.105 41.725 226.425 41.785 ;
        RECT 212.765 41.585 226.425 41.725 ;
        RECT 198.045 41.525 198.365 41.585 ;
        RECT 212.765 41.525 213.085 41.585 ;
        RECT 226.105 41.525 226.425 41.585 ;
        RECT 239.000 41.725 239.290 41.770 ;
        RECT 239.445 41.725 239.765 41.785 ;
        RECT 239.000 41.585 239.765 41.725 ;
        RECT 239.000 41.540 239.290 41.585 ;
        RECT 239.445 41.525 239.765 41.585 ;
        RECT 241.745 41.725 242.065 41.785 ;
        RECT 253.795 41.725 253.935 41.865 ;
        RECT 241.745 41.585 253.935 41.725 ;
        RECT 241.745 41.525 242.065 41.585 ;
        RECT 254.625 41.525 254.945 41.785 ;
        RECT 256.005 41.725 256.325 41.785 ;
        RECT 261.155 41.725 261.295 41.880 ;
        RECT 267.045 41.865 267.365 41.925 ;
        RECT 268.425 41.865 268.745 42.125 ;
        RECT 274.020 42.110 274.310 42.205 ;
        RECT 270.720 42.065 271.370 42.110 ;
        RECT 274.020 42.065 274.610 42.110 ;
        RECT 270.720 41.925 274.610 42.065 ;
        RECT 278.175 42.065 278.315 42.265 ;
        RECT 278.560 42.220 278.850 42.450 ;
        RECT 279.020 42.405 279.310 42.450 ;
        RECT 280.385 42.405 280.705 42.465 ;
        RECT 279.020 42.265 280.705 42.405 ;
        RECT 279.020 42.220 279.310 42.265 ;
        RECT 279.095 42.065 279.235 42.220 ;
        RECT 280.385 42.205 280.705 42.265 ;
        RECT 281.305 42.405 281.625 42.465 ;
        RECT 283.620 42.405 283.910 42.450 ;
        RECT 281.305 42.265 283.910 42.405 ;
        RECT 281.305 42.205 281.625 42.265 ;
        RECT 283.620 42.220 283.910 42.265 ;
        RECT 284.525 42.205 284.845 42.465 ;
        RECT 306.145 42.205 306.465 42.465 ;
        RECT 278.175 41.925 279.235 42.065 ;
        RECT 279.940 42.065 280.230 42.110 ;
        RECT 280.860 42.065 281.150 42.110 ;
        RECT 285.920 42.065 286.210 42.110 ;
        RECT 279.940 41.925 281.150 42.065 ;
        RECT 270.720 41.880 271.370 41.925 ;
        RECT 274.320 41.880 274.610 41.925 ;
        RECT 279.940 41.880 280.230 41.925 ;
        RECT 280.860 41.880 281.150 41.925 ;
        RECT 281.395 41.925 286.210 42.065 ;
        RECT 256.005 41.585 261.295 41.725 ;
        RECT 264.745 41.725 265.065 41.785 ;
        RECT 268.515 41.725 268.655 41.865 ;
        RECT 264.745 41.585 268.655 41.725 ;
        RECT 279.465 41.725 279.785 41.785 ;
        RECT 281.395 41.725 281.535 41.925 ;
        RECT 285.920 41.880 286.210 41.925 ;
        RECT 279.465 41.585 281.535 41.725 ;
        RECT 256.005 41.525 256.325 41.585 ;
        RECT 264.745 41.525 265.065 41.585 ;
        RECT 279.465 41.525 279.785 41.585 ;
        RECT 307.065 41.525 307.385 41.785 ;
        RECT 162.095 40.905 311.135 41.385 ;
        RECT 167.225 40.705 167.545 40.765 ;
        RECT 176.900 40.705 177.190 40.750 ;
        RECT 167.225 40.565 177.190 40.705 ;
        RECT 167.225 40.505 167.545 40.565 ;
        RECT 176.900 40.520 177.190 40.565 ;
        RECT 178.740 40.705 179.030 40.750 ;
        RECT 183.785 40.705 184.105 40.765 ;
        RECT 178.740 40.565 184.105 40.705 ;
        RECT 178.740 40.520 179.030 40.565 ;
        RECT 183.785 40.505 184.105 40.565 ;
        RECT 186.085 40.705 186.405 40.765 ;
        RECT 188.400 40.705 188.690 40.750 ;
        RECT 186.085 40.565 188.690 40.705 ;
        RECT 186.085 40.505 186.405 40.565 ;
        RECT 188.400 40.520 188.690 40.565 ;
        RECT 190.225 40.505 190.545 40.765 ;
        RECT 191.605 40.705 191.925 40.765 ;
        RECT 193.000 40.705 193.290 40.750 ;
        RECT 196.205 40.705 196.525 40.765 ;
        RECT 191.605 40.565 196.525 40.705 ;
        RECT 191.605 40.505 191.925 40.565 ;
        RECT 193.000 40.520 193.290 40.565 ;
        RECT 196.205 40.505 196.525 40.565 ;
        RECT 197.125 40.705 197.445 40.765 ;
        RECT 204.500 40.705 204.790 40.750 ;
        RECT 211.845 40.705 212.165 40.765 ;
        RECT 197.125 40.565 198.275 40.705 ;
        RECT 197.125 40.505 197.445 40.565 ;
        RECT 172.285 40.410 172.605 40.425 ;
        RECT 169.180 40.365 169.470 40.410 ;
        RECT 172.285 40.365 173.070 40.410 ;
        RECT 169.180 40.225 173.070 40.365 ;
        RECT 169.180 40.180 169.770 40.225 ;
        RECT 169.480 39.865 169.770 40.180 ;
        RECT 172.285 40.180 173.070 40.225 ;
        RECT 184.260 40.365 184.550 40.410 ;
        RECT 185.625 40.365 185.945 40.425 ;
        RECT 190.700 40.365 190.990 40.410 ;
        RECT 197.585 40.365 197.905 40.425 ;
        RECT 184.260 40.225 190.990 40.365 ;
        RECT 184.260 40.180 184.550 40.225 ;
        RECT 172.285 40.165 172.605 40.180 ;
        RECT 185.625 40.165 185.945 40.225 ;
        RECT 190.700 40.180 190.990 40.225 ;
        RECT 195.375 40.225 197.905 40.365 ;
        RECT 198.135 40.365 198.275 40.565 ;
        RECT 204.500 40.565 212.165 40.705 ;
        RECT 204.500 40.520 204.790 40.565 ;
        RECT 211.845 40.505 212.165 40.565 ;
        RECT 219.665 40.705 219.985 40.765 ;
        RECT 224.725 40.705 225.045 40.765 ;
        RECT 227.040 40.705 227.330 40.750 ;
        RECT 227.945 40.705 228.265 40.765 ;
        RECT 219.665 40.565 223.115 40.705 ;
        RECT 219.665 40.505 219.985 40.565 ;
        RECT 198.505 40.365 198.825 40.425 ;
        RECT 199.420 40.365 200.070 40.410 ;
        RECT 203.020 40.365 203.310 40.410 ;
        RECT 198.135 40.225 203.310 40.365 ;
        RECT 170.560 40.025 170.850 40.070 ;
        RECT 174.140 40.025 174.430 40.070 ;
        RECT 175.975 40.025 176.265 40.070 ;
        RECT 170.560 39.885 176.265 40.025 ;
        RECT 170.560 39.840 170.850 39.885 ;
        RECT 174.140 39.840 174.430 39.885 ;
        RECT 175.975 39.840 176.265 39.885 ;
        RECT 187.005 40.025 187.325 40.085 ;
        RECT 193.460 40.025 193.750 40.070 ;
        RECT 187.005 39.885 189.995 40.025 ;
        RECT 187.005 39.825 187.325 39.885 ;
        RECT 164.480 39.685 164.770 39.730 ;
        RECT 167.700 39.685 167.990 39.730 ;
        RECT 164.480 39.545 167.990 39.685 ;
        RECT 164.480 39.500 164.770 39.545 ;
        RECT 167.700 39.500 167.990 39.545 ;
        RECT 175.045 39.485 175.365 39.745 ;
        RECT 176.440 39.500 176.730 39.730 ;
        RECT 176.885 39.685 177.205 39.745 ;
        RECT 179.200 39.685 179.490 39.730 ;
        RECT 176.885 39.545 179.490 39.685 ;
        RECT 170.560 39.345 170.850 39.390 ;
        RECT 173.680 39.345 173.970 39.390 ;
        RECT 175.570 39.345 175.860 39.390 ;
        RECT 170.560 39.205 175.860 39.345 ;
        RECT 176.515 39.345 176.655 39.500 ;
        RECT 176.885 39.485 177.205 39.545 ;
        RECT 179.200 39.500 179.490 39.545 ;
        RECT 179.660 39.685 179.950 39.730 ;
        RECT 180.105 39.685 180.425 39.745 ;
        RECT 179.660 39.545 180.425 39.685 ;
        RECT 179.660 39.500 179.950 39.545 ;
        RECT 180.105 39.485 180.425 39.545 ;
        RECT 187.465 39.485 187.785 39.745 ;
        RECT 189.855 39.685 189.995 39.885 ;
        RECT 190.775 39.885 193.750 40.025 ;
        RECT 190.775 39.685 190.915 39.885 ;
        RECT 193.460 39.840 193.750 39.885 ;
        RECT 189.855 39.545 190.915 39.685 ;
        RECT 191.620 39.685 191.910 39.730 ;
        RECT 195.375 39.685 195.515 40.225 ;
        RECT 197.585 40.165 197.905 40.225 ;
        RECT 198.505 40.165 198.825 40.225 ;
        RECT 199.420 40.180 200.070 40.225 ;
        RECT 202.720 40.180 203.310 40.225 ;
        RECT 215.640 40.365 215.930 40.410 ;
        RECT 217.825 40.365 218.145 40.425 ;
        RECT 218.880 40.365 219.530 40.410 ;
        RECT 215.640 40.225 219.530 40.365 ;
        RECT 215.640 40.180 216.230 40.225 ;
        RECT 196.225 40.025 196.515 40.070 ;
        RECT 198.060 40.025 198.350 40.070 ;
        RECT 201.640 40.025 201.930 40.070 ;
        RECT 196.225 39.885 201.930 40.025 ;
        RECT 196.225 39.840 196.515 39.885 ;
        RECT 198.060 39.840 198.350 39.885 ;
        RECT 201.640 39.840 201.930 39.885 ;
        RECT 202.720 39.865 203.010 40.180 ;
        RECT 215.940 39.865 216.230 40.180 ;
        RECT 217.825 40.165 218.145 40.225 ;
        RECT 218.880 40.180 219.530 40.225 ;
        RECT 222.975 40.070 223.115 40.565 ;
        RECT 224.725 40.565 228.265 40.705 ;
        RECT 224.725 40.505 225.045 40.565 ;
        RECT 227.040 40.520 227.330 40.565 ;
        RECT 227.945 40.505 228.265 40.565 ;
        RECT 239.905 40.505 240.225 40.765 ;
        RECT 244.045 40.705 244.365 40.765 ;
        RECT 249.565 40.705 249.885 40.765 ;
        RECT 258.320 40.705 258.610 40.750 ;
        RECT 244.045 40.565 249.885 40.705 ;
        RECT 244.045 40.505 244.365 40.565 ;
        RECT 249.565 40.505 249.885 40.565 ;
        RECT 251.035 40.565 258.610 40.705 ;
        RECT 226.580 40.365 226.870 40.410 ;
        RECT 231.180 40.365 231.470 40.410 ;
        RECT 235.305 40.365 235.625 40.425 ;
        RECT 226.580 40.225 235.625 40.365 ;
        RECT 226.580 40.180 226.870 40.225 ;
        RECT 231.180 40.180 231.470 40.225 ;
        RECT 235.305 40.165 235.625 40.225 ;
        RECT 235.780 40.365 236.070 40.410 ;
        RECT 248.645 40.365 248.965 40.425 ;
        RECT 235.780 40.225 248.965 40.365 ;
        RECT 235.780 40.180 236.070 40.225 ;
        RECT 248.645 40.165 248.965 40.225 ;
        RECT 217.020 40.025 217.310 40.070 ;
        RECT 220.600 40.025 220.890 40.070 ;
        RECT 222.435 40.025 222.725 40.070 ;
        RECT 217.020 39.885 222.725 40.025 ;
        RECT 217.020 39.840 217.310 39.885 ;
        RECT 220.600 39.840 220.890 39.885 ;
        RECT 222.435 39.840 222.725 39.885 ;
        RECT 222.900 40.025 223.190 40.070 ;
        RECT 227.025 40.025 227.345 40.085 ;
        RECT 222.900 39.885 227.345 40.025 ;
        RECT 222.900 39.840 223.190 39.885 ;
        RECT 227.025 39.825 227.345 39.885 ;
        RECT 231.640 40.025 231.930 40.070 ;
        RECT 234.845 40.025 235.165 40.085 ;
        RECT 231.640 39.885 235.165 40.025 ;
        RECT 231.640 39.840 231.930 39.885 ;
        RECT 234.845 39.825 235.165 39.885 ;
        RECT 238.525 40.025 238.845 40.085 ;
        RECT 240.840 40.025 241.130 40.070 ;
        RECT 238.525 39.885 241.130 40.025 ;
        RECT 238.525 39.825 238.845 39.885 ;
        RECT 240.840 39.840 241.130 39.885 ;
        RECT 241.745 39.825 242.065 40.085 ;
        RECT 244.520 40.025 244.810 40.070 ;
        RECT 248.200 40.025 248.490 40.070 ;
        RECT 250.500 40.025 250.790 40.070 ;
        RECT 244.520 39.885 250.790 40.025 ;
        RECT 244.520 39.840 244.810 39.885 ;
        RECT 248.200 39.840 248.490 39.885 ;
        RECT 250.500 39.840 250.790 39.885 ;
        RECT 191.620 39.545 195.515 39.685 ;
        RECT 191.620 39.500 191.910 39.545 ;
        RECT 195.745 39.485 196.065 39.745 ;
        RECT 197.140 39.685 197.430 39.730 ;
        RECT 197.585 39.685 197.905 39.745 ;
        RECT 197.140 39.545 197.905 39.685 ;
        RECT 197.140 39.500 197.430 39.545 ;
        RECT 197.585 39.485 197.905 39.545 ;
        RECT 207.705 39.485 208.025 39.745 ;
        RECT 213.240 39.685 213.530 39.730 ;
        RECT 214.160 39.685 214.450 39.730 ;
        RECT 213.240 39.545 214.450 39.685 ;
        RECT 213.240 39.500 213.530 39.545 ;
        RECT 214.160 39.500 214.450 39.545 ;
        RECT 221.505 39.485 221.825 39.745 ;
        RECT 226.105 39.685 226.425 39.745 ;
        RECT 231.165 39.685 231.485 39.745 ;
        RECT 232.100 39.685 232.390 39.730 ;
        RECT 226.105 39.545 230.935 39.685 ;
        RECT 226.105 39.485 226.425 39.545 ;
        RECT 195.835 39.345 195.975 39.485 ;
        RECT 176.515 39.205 195.975 39.345 ;
        RECT 196.630 39.345 196.920 39.390 ;
        RECT 198.520 39.345 198.810 39.390 ;
        RECT 201.640 39.345 201.930 39.390 ;
        RECT 196.630 39.205 201.930 39.345 ;
        RECT 170.560 39.160 170.850 39.205 ;
        RECT 173.680 39.160 173.970 39.205 ;
        RECT 175.570 39.160 175.860 39.205 ;
        RECT 196.630 39.160 196.920 39.205 ;
        RECT 198.520 39.160 198.810 39.205 ;
        RECT 201.640 39.160 201.930 39.205 ;
        RECT 202.185 39.345 202.505 39.405 ;
        RECT 204.960 39.345 205.250 39.390 ;
        RECT 202.185 39.205 205.250 39.345 ;
        RECT 202.185 39.145 202.505 39.205 ;
        RECT 204.960 39.160 205.250 39.205 ;
        RECT 217.020 39.345 217.310 39.390 ;
        RECT 220.140 39.345 220.430 39.390 ;
        RECT 222.030 39.345 222.320 39.390 ;
        RECT 217.020 39.205 222.320 39.345 ;
        RECT 217.020 39.160 217.310 39.205 ;
        RECT 220.140 39.160 220.430 39.205 ;
        RECT 222.030 39.160 222.320 39.205 ;
        RECT 227.485 39.345 227.805 39.405 ;
        RECT 229.340 39.345 229.630 39.390 ;
        RECT 227.485 39.205 229.630 39.345 ;
        RECT 230.795 39.345 230.935 39.545 ;
        RECT 231.165 39.545 232.390 39.685 ;
        RECT 231.165 39.485 231.485 39.545 ;
        RECT 232.100 39.500 232.390 39.545 ;
        RECT 235.765 39.685 236.085 39.745 ;
        RECT 236.240 39.685 236.530 39.730 ;
        RECT 235.765 39.545 236.530 39.685 ;
        RECT 235.765 39.485 236.085 39.545 ;
        RECT 236.240 39.500 236.530 39.545 ;
        RECT 236.685 39.485 237.005 39.745 ;
        RECT 244.980 39.500 245.270 39.730 ;
        RECT 245.055 39.345 245.195 39.500 ;
        RECT 248.645 39.485 248.965 39.745 ;
        RECT 249.120 39.685 249.410 39.730 ;
        RECT 251.035 39.685 251.175 40.565 ;
        RECT 258.320 40.520 258.610 40.565 ;
        RECT 258.765 40.705 259.085 40.765 ;
        RECT 265.205 40.705 265.525 40.765 ;
        RECT 258.765 40.565 265.525 40.705 ;
        RECT 258.765 40.505 259.085 40.565 ;
        RECT 259.315 40.070 259.455 40.565 ;
        RECT 265.205 40.505 265.525 40.565 ;
        RECT 271.660 40.705 271.950 40.750 ;
        RECT 283.605 40.705 283.925 40.765 ;
        RECT 289.585 40.705 289.905 40.765 ;
        RECT 303.385 40.705 303.705 40.765 ;
        RECT 308.000 40.705 308.290 40.750 ;
        RECT 271.660 40.565 280.155 40.705 ;
        RECT 271.660 40.520 271.950 40.565 ;
        RECT 269.345 40.365 269.665 40.425 ;
        RECT 270.265 40.365 270.585 40.425 ;
        RECT 269.345 40.225 270.585 40.365 ;
        RECT 269.345 40.165 269.665 40.225 ;
        RECT 270.265 40.165 270.585 40.225 ;
        RECT 273.600 40.365 273.890 40.410 ;
        RECT 276.840 40.365 277.490 40.410 ;
        RECT 273.600 40.225 277.490 40.365 ;
        RECT 273.600 40.180 274.190 40.225 ;
        RECT 276.840 40.180 277.490 40.225 ;
        RECT 273.900 40.085 274.190 40.180 ;
        RECT 279.465 40.165 279.785 40.425 ;
        RECT 280.015 40.365 280.155 40.565 ;
        RECT 283.605 40.565 289.905 40.705 ;
        RECT 283.605 40.505 283.925 40.565 ;
        RECT 289.585 40.505 289.905 40.565 ;
        RECT 293.355 40.565 308.290 40.705 ;
        RECT 286.365 40.410 286.685 40.425 ;
        RECT 282.800 40.365 283.090 40.410 ;
        RECT 286.040 40.365 286.690 40.410 ;
        RECT 293.355 40.365 293.495 40.565 ;
        RECT 303.385 40.505 303.705 40.565 ;
        RECT 308.000 40.520 308.290 40.565 ;
        RECT 280.015 40.225 281.995 40.365 ;
        RECT 256.480 39.840 256.770 40.070 ;
        RECT 257.400 40.025 257.690 40.070 ;
        RECT 257.400 39.885 258.995 40.025 ;
        RECT 257.400 39.840 257.690 39.885 ;
        RECT 249.120 39.545 251.175 39.685 ;
        RECT 249.120 39.500 249.410 39.545 ;
        RECT 230.795 39.205 245.195 39.345 ;
        RECT 248.185 39.345 248.505 39.405 ;
        RECT 249.195 39.345 249.335 39.500 ;
        RECT 253.245 39.485 253.565 39.745 ;
        RECT 256.555 39.685 256.695 39.840 ;
        RECT 258.305 39.685 258.625 39.745 ;
        RECT 256.555 39.545 258.625 39.685 ;
        RECT 258.855 39.685 258.995 39.885 ;
        RECT 259.240 39.840 259.530 40.070 ;
        RECT 260.145 39.825 260.465 40.085 ;
        RECT 262.920 39.840 263.210 40.070 ;
        RECT 271.660 40.025 271.950 40.070 ;
        RECT 272.105 40.025 272.425 40.085 ;
        RECT 271.660 39.885 272.425 40.025 ;
        RECT 271.660 39.840 271.950 39.885 ;
        RECT 259.685 39.685 260.005 39.745 ;
        RECT 258.855 39.545 260.005 39.685 ;
        RECT 258.305 39.485 258.625 39.545 ;
        RECT 259.685 39.485 260.005 39.545 ;
        RECT 248.185 39.205 249.335 39.345 ;
        RECT 256.925 39.345 257.245 39.405 ;
        RECT 262.000 39.345 262.290 39.390 ;
        RECT 256.925 39.205 262.290 39.345 ;
        RECT 227.485 39.145 227.805 39.205 ;
        RECT 229.340 39.160 229.630 39.205 ;
        RECT 248.185 39.145 248.505 39.205 ;
        RECT 256.925 39.145 257.245 39.205 ;
        RECT 262.000 39.160 262.290 39.205 ;
        RECT 167.240 39.005 167.530 39.050 ;
        RECT 179.645 39.005 179.965 39.065 ;
        RECT 167.240 38.865 179.965 39.005 ;
        RECT 167.240 38.820 167.530 38.865 ;
        RECT 179.645 38.805 179.965 38.865 ;
        RECT 210.020 39.005 210.310 39.050 ;
        RECT 214.605 39.005 214.925 39.065 ;
        RECT 216.445 39.005 216.765 39.065 ;
        RECT 210.020 38.865 216.765 39.005 ;
        RECT 210.020 38.820 210.310 38.865 ;
        RECT 214.605 38.805 214.925 38.865 ;
        RECT 216.445 38.805 216.765 38.865 ;
        RECT 228.880 39.005 229.170 39.050 ;
        RECT 231.625 39.005 231.945 39.065 ;
        RECT 228.880 38.865 231.945 39.005 ;
        RECT 228.880 38.820 229.170 38.865 ;
        RECT 231.625 38.805 231.945 38.865 ;
        RECT 232.085 39.005 232.405 39.065 ;
        RECT 233.940 39.005 234.230 39.050 ;
        RECT 232.085 38.865 234.230 39.005 ;
        RECT 232.085 38.805 232.405 38.865 ;
        RECT 233.940 38.820 234.230 38.865 ;
        RECT 242.205 38.805 242.525 39.065 ;
        RECT 243.125 39.005 243.445 39.065 ;
        RECT 246.360 39.005 246.650 39.050 ;
        RECT 243.125 38.865 246.650 39.005 ;
        RECT 243.125 38.805 243.445 38.865 ;
        RECT 246.360 38.820 246.650 38.865 ;
        RECT 257.400 39.005 257.690 39.050 ;
        RECT 262.995 39.005 263.135 39.840 ;
        RECT 272.105 39.825 272.425 39.885 ;
        RECT 273.900 39.865 274.265 40.085 ;
        RECT 273.945 39.825 274.265 39.865 ;
        RECT 274.980 40.025 275.270 40.070 ;
        RECT 278.560 40.025 278.850 40.070 ;
        RECT 280.395 40.025 280.685 40.070 ;
        RECT 274.980 39.885 280.685 40.025 ;
        RECT 274.980 39.840 275.270 39.885 ;
        RECT 278.560 39.840 278.850 39.885 ;
        RECT 280.395 39.840 280.685 39.885 ;
        RECT 264.300 39.685 264.590 39.730 ;
        RECT 265.680 39.685 265.970 39.730 ;
        RECT 264.300 39.545 265.970 39.685 ;
        RECT 264.300 39.500 264.590 39.545 ;
        RECT 265.680 39.500 265.970 39.545 ;
        RECT 267.505 39.685 267.825 39.745 ;
        RECT 268.440 39.685 268.730 39.730 ;
        RECT 267.505 39.545 268.730 39.685 ;
        RECT 274.035 39.685 274.175 39.825 ;
        RECT 274.035 39.545 280.615 39.685 ;
        RECT 267.505 39.485 267.825 39.545 ;
        RECT 268.440 39.500 268.730 39.545 ;
        RECT 263.840 39.345 264.130 39.390 ;
        RECT 269.805 39.345 270.125 39.405 ;
        RECT 271.200 39.345 271.490 39.390 ;
        RECT 263.840 39.205 271.490 39.345 ;
        RECT 263.840 39.160 264.130 39.205 ;
        RECT 269.805 39.145 270.125 39.205 ;
        RECT 271.200 39.160 271.490 39.205 ;
        RECT 274.980 39.345 275.270 39.390 ;
        RECT 278.100 39.345 278.390 39.390 ;
        RECT 279.990 39.345 280.280 39.390 ;
        RECT 274.980 39.205 280.280 39.345 ;
        RECT 274.980 39.160 275.270 39.205 ;
        RECT 278.100 39.160 278.390 39.205 ;
        RECT 279.990 39.160 280.280 39.205 ;
        RECT 257.400 38.865 263.135 39.005 ;
        RECT 257.400 38.820 257.690 38.865 ;
        RECT 272.105 38.805 272.425 39.065 ;
        RECT 280.475 39.005 280.615 39.545 ;
        RECT 280.860 39.500 281.150 39.730 ;
        RECT 280.935 39.345 281.075 39.500 ;
        RECT 281.305 39.485 281.625 39.745 ;
        RECT 281.855 39.685 281.995 40.225 ;
        RECT 282.800 40.225 293.495 40.365 ;
        RECT 301.540 40.365 302.190 40.410 ;
        RECT 302.925 40.365 303.245 40.425 ;
        RECT 305.140 40.365 305.430 40.410 ;
        RECT 301.540 40.225 305.430 40.365 ;
        RECT 282.800 40.180 283.390 40.225 ;
        RECT 286.040 40.180 286.690 40.225 ;
        RECT 301.540 40.180 302.190 40.225 ;
        RECT 283.100 39.865 283.390 40.180 ;
        RECT 286.365 40.165 286.685 40.180 ;
        RECT 302.925 40.165 303.245 40.225 ;
        RECT 304.840 40.180 305.430 40.225 ;
        RECT 284.180 40.025 284.470 40.070 ;
        RECT 287.760 40.025 288.050 40.070 ;
        RECT 289.595 40.025 289.885 40.070 ;
        RECT 284.180 39.885 289.885 40.025 ;
        RECT 284.180 39.840 284.470 39.885 ;
        RECT 287.760 39.840 288.050 39.885 ;
        RECT 289.595 39.840 289.885 39.885 ;
        RECT 298.345 40.025 298.635 40.070 ;
        RECT 300.180 40.025 300.470 40.070 ;
        RECT 303.760 40.025 304.050 40.070 ;
        RECT 298.345 39.885 304.050 40.025 ;
        RECT 298.345 39.840 298.635 39.885 ;
        RECT 300.180 39.840 300.470 39.885 ;
        RECT 303.760 39.840 304.050 39.885 ;
        RECT 304.840 39.865 305.130 40.180 ;
        RECT 307.065 39.825 307.385 40.085 ;
        RECT 288.680 39.685 288.970 39.730 ;
        RECT 281.855 39.545 288.970 39.685 ;
        RECT 288.680 39.500 288.970 39.545 ;
        RECT 290.045 39.685 290.365 39.745 ;
        RECT 297.880 39.685 298.170 39.730 ;
        RECT 299.260 39.685 299.550 39.730 ;
        RECT 307.525 39.685 307.845 39.745 ;
        RECT 290.045 39.545 298.555 39.685 ;
        RECT 290.045 39.485 290.365 39.545 ;
        RECT 297.880 39.500 298.170 39.545 ;
        RECT 283.605 39.345 283.925 39.405 ;
        RECT 280.935 39.205 283.925 39.345 ;
        RECT 283.605 39.145 283.925 39.205 ;
        RECT 284.180 39.345 284.470 39.390 ;
        RECT 287.300 39.345 287.590 39.390 ;
        RECT 289.190 39.345 289.480 39.390 ;
        RECT 284.180 39.205 289.480 39.345 ;
        RECT 284.180 39.160 284.470 39.205 ;
        RECT 287.300 39.160 287.590 39.205 ;
        RECT 289.190 39.160 289.480 39.205 ;
        RECT 286.365 39.005 286.685 39.065 ;
        RECT 280.475 38.865 286.685 39.005 ;
        RECT 298.415 39.005 298.555 39.545 ;
        RECT 299.260 39.545 307.845 39.685 ;
        RECT 299.260 39.500 299.550 39.545 ;
        RECT 307.525 39.485 307.845 39.545 ;
        RECT 298.750 39.345 299.040 39.390 ;
        RECT 300.640 39.345 300.930 39.390 ;
        RECT 303.760 39.345 304.050 39.390 ;
        RECT 298.750 39.205 304.050 39.345 ;
        RECT 298.750 39.160 299.040 39.205 ;
        RECT 300.640 39.160 300.930 39.205 ;
        RECT 303.760 39.160 304.050 39.205 ;
        RECT 305.685 39.005 306.005 39.065 ;
        RECT 298.415 38.865 306.005 39.005 ;
        RECT 286.365 38.805 286.685 38.865 ;
        RECT 305.685 38.805 306.005 38.865 ;
        RECT 306.605 38.805 306.925 39.065 ;
        RECT 162.095 38.185 311.135 38.665 ;
        RECT 170.920 37.985 171.210 38.030 ;
        RECT 175.045 37.985 175.365 38.045 ;
        RECT 170.920 37.845 175.365 37.985 ;
        RECT 170.920 37.800 171.210 37.845 ;
        RECT 175.045 37.785 175.365 37.845 ;
        RECT 185.640 37.985 185.930 38.030 ;
        RECT 187.005 37.985 187.325 38.045 ;
        RECT 185.640 37.845 187.325 37.985 ;
        RECT 185.640 37.800 185.930 37.845 ;
        RECT 187.005 37.785 187.325 37.845 ;
        RECT 203.580 37.985 203.870 38.030 ;
        RECT 207.705 37.985 208.025 38.045 ;
        RECT 203.580 37.845 208.025 37.985 ;
        RECT 203.580 37.800 203.870 37.845 ;
        RECT 207.705 37.785 208.025 37.845 ;
        RECT 221.505 37.985 221.825 38.045 ;
        RECT 222.440 37.985 222.730 38.030 ;
        RECT 221.505 37.845 222.730 37.985 ;
        RECT 221.505 37.785 221.825 37.845 ;
        RECT 222.440 37.800 222.730 37.845 ;
        RECT 230.705 37.985 231.025 38.045 ;
        RECT 248.185 37.985 248.505 38.045 ;
        RECT 230.705 37.845 248.505 37.985 ;
        RECT 230.705 37.785 231.025 37.845 ;
        RECT 248.185 37.785 248.505 37.845 ;
        RECT 249.565 37.785 249.885 38.045 ;
        RECT 255.100 37.985 255.390 38.030 ;
        RECT 256.005 37.985 256.325 38.045 ;
        RECT 255.100 37.845 256.325 37.985 ;
        RECT 255.100 37.800 255.390 37.845 ;
        RECT 256.005 37.785 256.325 37.845 ;
        RECT 260.145 37.985 260.465 38.045 ;
        RECT 267.980 37.985 268.270 38.030 ;
        RECT 260.145 37.845 268.270 37.985 ;
        RECT 260.145 37.785 260.465 37.845 ;
        RECT 267.980 37.800 268.270 37.845 ;
        RECT 268.425 37.985 268.745 38.045 ;
        RECT 269.805 37.985 270.125 38.045 ;
        RECT 268.425 37.845 276.475 37.985 ;
        RECT 268.425 37.785 268.745 37.845 ;
        RECT 269.805 37.785 270.125 37.845 ;
        RECT 175.520 37.645 175.810 37.690 ;
        RECT 168.235 37.505 175.810 37.645 ;
        RECT 168.235 37.350 168.375 37.505 ;
        RECT 175.520 37.460 175.810 37.505 ;
        RECT 188.500 37.645 188.790 37.690 ;
        RECT 191.620 37.645 191.910 37.690 ;
        RECT 193.510 37.645 193.800 37.690 ;
        RECT 188.500 37.505 193.800 37.645 ;
        RECT 188.500 37.460 188.790 37.505 ;
        RECT 191.620 37.460 191.910 37.505 ;
        RECT 193.510 37.460 193.800 37.505 ;
        RECT 198.505 37.645 198.825 37.705 ;
        RECT 211.860 37.645 212.150 37.690 ;
        RECT 198.505 37.505 212.150 37.645 ;
        RECT 198.505 37.445 198.825 37.505 ;
        RECT 211.860 37.460 212.150 37.505 ;
        RECT 218.300 37.645 218.590 37.690 ;
        RECT 231.130 37.645 231.420 37.690 ;
        RECT 233.020 37.645 233.310 37.690 ;
        RECT 236.140 37.645 236.430 37.690 ;
        RECT 218.300 37.505 219.435 37.645 ;
        RECT 218.300 37.460 218.590 37.505 ;
        RECT 168.160 37.120 168.450 37.350 ;
        RECT 178.725 37.305 179.045 37.365 ;
        RECT 180.105 37.305 180.425 37.365 ;
        RECT 178.725 37.165 180.425 37.305 ;
        RECT 178.725 37.105 179.045 37.165 ;
        RECT 180.105 37.105 180.425 37.165 ;
        RECT 185.180 37.305 185.470 37.350 ;
        RECT 187.005 37.305 187.325 37.365 ;
        RECT 192.525 37.305 192.845 37.365 ;
        RECT 185.180 37.165 192.845 37.305 ;
        RECT 185.180 37.120 185.470 37.165 ;
        RECT 187.005 37.105 187.325 37.165 ;
        RECT 192.525 37.105 192.845 37.165 ;
        RECT 194.380 37.305 194.670 37.350 ;
        RECT 195.745 37.305 196.065 37.365 ;
        RECT 197.125 37.305 197.445 37.365 ;
        RECT 194.380 37.165 197.445 37.305 ;
        RECT 194.380 37.120 194.670 37.165 ;
        RECT 195.745 37.105 196.065 37.165 ;
        RECT 197.125 37.105 197.445 37.165 ;
        RECT 197.585 37.305 197.905 37.365 ;
        RECT 219.295 37.350 219.435 37.505 ;
        RECT 231.130 37.505 236.430 37.645 ;
        RECT 231.130 37.460 231.420 37.505 ;
        RECT 233.020 37.460 233.310 37.505 ;
        RECT 236.140 37.460 236.430 37.505 ;
        RECT 237.145 37.645 237.465 37.705 ;
        RECT 241.710 37.645 242.000 37.690 ;
        RECT 243.600 37.645 243.890 37.690 ;
        RECT 246.720 37.645 247.010 37.690 ;
        RECT 237.145 37.505 239.675 37.645 ;
        RECT 237.145 37.445 237.465 37.505 ;
        RECT 206.800 37.305 207.090 37.350 ;
        RECT 215.540 37.305 215.830 37.350 ;
        RECT 197.585 37.165 217.135 37.305 ;
        RECT 197.585 37.105 197.905 37.165 ;
        RECT 206.800 37.120 207.090 37.165 ;
        RECT 215.540 37.120 215.830 37.165 ;
        RECT 171.365 36.765 171.685 37.025 ;
        RECT 175.045 36.965 175.365 37.025 ;
        RECT 177.820 36.965 178.110 37.010 ;
        RECT 175.045 36.825 178.110 36.965 ;
        RECT 175.045 36.765 175.365 36.825 ;
        RECT 177.820 36.780 178.110 36.825 ;
        RECT 182.420 36.965 182.710 37.010 ;
        RECT 182.865 36.965 183.185 37.025 ;
        RECT 182.420 36.825 183.185 36.965 ;
        RECT 182.420 36.780 182.710 36.825 ;
        RECT 182.865 36.765 183.185 36.825 ;
        RECT 174.600 36.625 174.890 36.670 ;
        RECT 176.885 36.625 177.205 36.685 ;
        RECT 174.600 36.485 177.205 36.625 ;
        RECT 174.600 36.440 174.890 36.485 ;
        RECT 176.885 36.425 177.205 36.485 ;
        RECT 177.360 36.625 177.650 36.670 ;
        RECT 179.645 36.625 179.965 36.685 ;
        RECT 187.420 36.670 187.710 36.985 ;
        RECT 188.500 36.965 188.790 37.010 ;
        RECT 192.080 36.965 192.370 37.010 ;
        RECT 193.915 36.965 194.205 37.010 ;
        RECT 188.500 36.825 194.205 36.965 ;
        RECT 188.500 36.780 188.790 36.825 ;
        RECT 192.080 36.780 192.370 36.825 ;
        RECT 193.915 36.780 194.205 36.825 ;
        RECT 195.285 36.765 195.605 37.025 ;
        RECT 205.420 36.965 205.710 37.010 ;
        RECT 205.865 36.965 206.185 37.025 ;
        RECT 207.720 36.965 208.010 37.010 ;
        RECT 205.420 36.825 208.010 36.965 ;
        RECT 205.420 36.780 205.710 36.825 ;
        RECT 205.865 36.765 206.185 36.825 ;
        RECT 207.720 36.780 208.010 36.825 ;
        RECT 209.085 36.965 209.405 37.025 ;
        RECT 210.480 36.965 210.770 37.010 ;
        RECT 209.085 36.825 210.770 36.965 ;
        RECT 209.085 36.765 209.405 36.825 ;
        RECT 210.480 36.780 210.770 36.825 ;
        RECT 216.445 36.765 216.765 37.025 ;
        RECT 216.995 36.965 217.135 37.165 ;
        RECT 219.220 37.120 219.510 37.350 ;
        RECT 223.360 37.305 223.650 37.350 ;
        RECT 227.485 37.305 227.805 37.365 ;
        RECT 223.360 37.165 227.805 37.305 ;
        RECT 223.360 37.120 223.650 37.165 ;
        RECT 227.485 37.105 227.805 37.165 ;
        RECT 227.945 37.305 228.265 37.365 ;
        RECT 239.000 37.305 239.290 37.350 ;
        RECT 227.945 37.165 239.290 37.305 ;
        RECT 227.945 37.105 228.265 37.165 ;
        RECT 239.000 37.120 239.290 37.165 ;
        RECT 227.025 36.965 227.345 37.025 ;
        RECT 230.260 36.965 230.550 37.010 ;
        RECT 216.995 36.825 226.795 36.965 ;
        RECT 177.360 36.485 179.965 36.625 ;
        RECT 177.360 36.440 177.650 36.485 ;
        RECT 179.645 36.425 179.965 36.485 ;
        RECT 187.120 36.625 187.710 36.670 ;
        RECT 190.360 36.625 191.010 36.670 ;
        RECT 193.000 36.625 193.290 36.670 ;
        RECT 194.365 36.625 194.685 36.685 ;
        RECT 187.120 36.485 192.755 36.625 ;
        RECT 187.120 36.440 187.410 36.485 ;
        RECT 190.360 36.440 191.010 36.485 ;
        RECT 192.615 36.285 192.755 36.485 ;
        RECT 193.000 36.485 194.685 36.625 ;
        RECT 193.000 36.440 193.290 36.485 ;
        RECT 194.365 36.425 194.685 36.485 ;
        RECT 208.625 36.625 208.945 36.685 ;
        RECT 213.240 36.625 213.530 36.670 ;
        RECT 225.645 36.625 225.965 36.685 ;
        RECT 208.625 36.485 225.965 36.625 ;
        RECT 226.655 36.625 226.795 36.825 ;
        RECT 227.025 36.825 230.550 36.965 ;
        RECT 227.025 36.765 227.345 36.825 ;
        RECT 230.260 36.780 230.550 36.825 ;
        RECT 230.725 36.965 231.015 37.010 ;
        RECT 232.560 36.965 232.850 37.010 ;
        RECT 236.140 36.965 236.430 37.010 ;
        RECT 230.725 36.825 236.430 36.965 ;
        RECT 230.725 36.780 231.015 36.825 ;
        RECT 232.560 36.780 232.850 36.825 ;
        RECT 236.140 36.780 236.430 36.825 ;
        RECT 231.165 36.625 231.485 36.685 ;
        RECT 226.655 36.485 231.485 36.625 ;
        RECT 208.625 36.425 208.945 36.485 ;
        RECT 213.240 36.440 213.530 36.485 ;
        RECT 225.645 36.425 225.965 36.485 ;
        RECT 231.165 36.425 231.485 36.485 ;
        RECT 231.625 36.425 231.945 36.685 ;
        RECT 237.220 36.670 237.510 36.985 ;
        RECT 233.920 36.625 234.570 36.670 ;
        RECT 237.220 36.625 237.810 36.670 ;
        RECT 239.535 36.625 239.675 37.505 ;
        RECT 241.710 37.505 247.010 37.645 ;
        RECT 241.710 37.460 242.000 37.505 ;
        RECT 243.600 37.460 243.890 37.505 ;
        RECT 246.720 37.460 247.010 37.505 ;
        RECT 257.960 37.645 258.250 37.690 ;
        RECT 261.080 37.645 261.370 37.690 ;
        RECT 262.970 37.645 263.260 37.690 ;
        RECT 267.060 37.645 267.350 37.690 ;
        RECT 276.335 37.645 276.475 37.845 ;
        RECT 278.545 37.785 278.865 38.045 ;
        RECT 281.305 37.985 281.625 38.045 ;
        RECT 283.160 37.985 283.450 38.030 ;
        RECT 281.305 37.845 283.450 37.985 ;
        RECT 281.305 37.785 281.625 37.845 ;
        RECT 283.160 37.800 283.450 37.845 ;
        RECT 305.700 37.985 305.990 38.030 ;
        RECT 306.145 37.985 306.465 38.045 ;
        RECT 305.700 37.845 306.465 37.985 ;
        RECT 305.700 37.800 305.990 37.845 ;
        RECT 306.145 37.785 306.465 37.845 ;
        RECT 282.240 37.645 282.530 37.690 ;
        RECT 257.960 37.505 263.260 37.645 ;
        RECT 257.960 37.460 258.250 37.505 ;
        RECT 261.080 37.460 261.370 37.505 ;
        RECT 262.970 37.460 263.260 37.505 ;
        RECT 263.455 37.505 267.350 37.645 ;
        RECT 240.825 37.105 241.145 37.365 ;
        RECT 242.205 37.105 242.525 37.365 ;
        RECT 244.965 37.305 245.285 37.365 ;
        RECT 262.460 37.305 262.750 37.350 ;
        RECT 263.455 37.305 263.595 37.505 ;
        RECT 267.060 37.460 267.350 37.505 ;
        RECT 269.665 37.505 276.015 37.645 ;
        RECT 276.335 37.505 282.530 37.645 ;
        RECT 244.965 37.165 257.155 37.305 ;
        RECT 244.965 37.105 245.285 37.165 ;
        RECT 241.305 36.965 241.595 37.010 ;
        RECT 243.140 36.965 243.430 37.010 ;
        RECT 246.720 36.965 247.010 37.010 ;
        RECT 257.015 36.985 257.155 37.165 ;
        RECT 262.460 37.165 263.595 37.305 ;
        RECT 263.825 37.305 264.145 37.365 ;
        RECT 266.585 37.305 266.905 37.365 ;
        RECT 263.825 37.165 266.905 37.305 ;
        RECT 262.460 37.120 262.750 37.165 ;
        RECT 263.825 37.105 264.145 37.165 ;
        RECT 266.585 37.105 266.905 37.165 ;
        RECT 241.305 36.825 247.010 36.965 ;
        RECT 241.305 36.780 241.595 36.825 ;
        RECT 243.140 36.780 243.430 36.825 ;
        RECT 246.720 36.780 247.010 36.825 ;
        RECT 241.745 36.625 242.065 36.685 ;
        RECT 244.965 36.670 245.285 36.685 ;
        RECT 233.920 36.485 242.065 36.625 ;
        RECT 233.920 36.440 234.570 36.485 ;
        RECT 237.520 36.440 237.810 36.485 ;
        RECT 241.745 36.425 242.065 36.485 ;
        RECT 244.500 36.625 245.285 36.670 ;
        RECT 247.800 36.670 248.090 36.985 ;
        RECT 256.880 36.965 257.170 36.985 ;
        RECT 257.385 36.965 257.705 37.025 ;
        RECT 256.880 36.825 257.705 36.965 ;
        RECT 256.880 36.670 257.170 36.825 ;
        RECT 257.385 36.765 257.705 36.825 ;
        RECT 257.960 36.965 258.250 37.010 ;
        RECT 261.540 36.965 261.830 37.010 ;
        RECT 263.375 36.965 263.665 37.010 ;
        RECT 269.665 36.965 269.805 37.505 ;
        RECT 272.105 37.305 272.425 37.365 ;
        RECT 275.875 37.350 276.015 37.505 ;
        RECT 282.240 37.460 282.530 37.505 ;
        RECT 284.525 37.645 284.845 37.705 ;
        RECT 285.000 37.645 285.290 37.690 ;
        RECT 284.525 37.505 285.290 37.645 ;
        RECT 284.525 37.445 284.845 37.505 ;
        RECT 285.000 37.460 285.290 37.505 ;
        RECT 275.340 37.305 275.630 37.350 ;
        RECT 272.105 37.165 275.630 37.305 ;
        RECT 272.105 37.105 272.425 37.165 ;
        RECT 275.340 37.120 275.630 37.165 ;
        RECT 275.800 37.120 276.090 37.350 ;
        RECT 284.615 37.305 284.755 37.445 ;
        RECT 276.335 37.165 284.755 37.305 ;
        RECT 257.960 36.825 263.665 36.965 ;
        RECT 257.960 36.780 258.250 36.825 ;
        RECT 261.540 36.780 261.830 36.825 ;
        RECT 263.375 36.780 263.665 36.825 ;
        RECT 263.915 36.825 269.805 36.965 ;
        RECT 270.265 36.965 270.585 37.025 ;
        RECT 274.880 36.965 275.170 37.010 ;
        RECT 270.265 36.825 275.170 36.965 ;
        RECT 275.415 36.965 275.555 37.120 ;
        RECT 276.335 36.965 276.475 37.165 ;
        RECT 306.605 37.105 306.925 37.365 ;
        RECT 275.415 36.825 276.475 36.965 ;
        RECT 247.800 36.625 248.390 36.670 ;
        RECT 244.500 36.485 248.390 36.625 ;
        RECT 244.500 36.440 245.285 36.485 ;
        RECT 248.100 36.440 248.390 36.485 ;
        RECT 256.580 36.625 257.170 36.670 ;
        RECT 259.820 36.625 260.470 36.670 ;
        RECT 256.580 36.485 260.470 36.625 ;
        RECT 256.580 36.440 256.870 36.485 ;
        RECT 259.820 36.440 260.470 36.485 ;
        RECT 244.965 36.425 245.285 36.440 ;
        RECT 193.445 36.285 193.765 36.345 ;
        RECT 192.615 36.145 193.765 36.285 ;
        RECT 193.445 36.085 193.765 36.145 ;
        RECT 193.905 36.285 194.225 36.345 ;
        RECT 198.060 36.285 198.350 36.330 ;
        RECT 193.905 36.145 198.350 36.285 ;
        RECT 193.905 36.085 194.225 36.145 ;
        RECT 198.060 36.100 198.350 36.145 ;
        RECT 205.865 36.085 206.185 36.345 ;
        RECT 215.985 36.085 216.305 36.345 ;
        RECT 226.105 36.085 226.425 36.345 ;
        RECT 228.405 36.285 228.725 36.345 ;
        RECT 236.685 36.285 237.005 36.345 ;
        RECT 263.915 36.285 264.055 36.825 ;
        RECT 270.265 36.765 270.585 36.825 ;
        RECT 274.880 36.780 275.170 36.825 ;
        RECT 277.625 36.765 277.945 37.025 ;
        RECT 281.765 36.765 282.085 37.025 ;
        RECT 304.765 36.765 305.085 37.025 ;
        RECT 264.745 36.625 265.065 36.685 ;
        RECT 267.045 36.625 267.365 36.685 ;
        RECT 267.820 36.625 268.110 36.670 ;
        RECT 264.745 36.485 265.895 36.625 ;
        RECT 264.745 36.425 265.065 36.485 ;
        RECT 228.405 36.145 264.055 36.285 ;
        RECT 228.405 36.085 228.725 36.145 ;
        RECT 236.685 36.085 237.005 36.145 ;
        RECT 265.205 36.085 265.525 36.345 ;
        RECT 265.755 36.285 265.895 36.485 ;
        RECT 267.045 36.485 268.110 36.625 ;
        RECT 267.045 36.425 267.365 36.485 ;
        RECT 267.820 36.440 268.110 36.485 ;
        RECT 268.885 36.425 269.205 36.685 ;
        RECT 277.715 36.625 277.855 36.765 ;
        RECT 283.160 36.625 283.450 36.670 ;
        RECT 277.715 36.485 283.450 36.625 ;
        RECT 283.160 36.440 283.450 36.485 ;
        RECT 306.605 36.285 306.925 36.345 ;
        RECT 265.755 36.145 306.925 36.285 ;
        RECT 306.605 36.085 306.925 36.145 ;
        RECT 307.065 36.285 307.385 36.345 ;
        RECT 309.380 36.285 309.670 36.330 ;
        RECT 307.065 36.145 309.670 36.285 ;
        RECT 307.065 36.085 307.385 36.145 ;
        RECT 309.380 36.100 309.670 36.145 ;
        RECT 162.095 35.465 311.135 35.945 ;
        RECT 165.860 35.265 166.150 35.310 ;
        RECT 171.365 35.265 171.685 35.325 ;
        RECT 165.860 35.125 171.685 35.265 ;
        RECT 165.860 35.080 166.150 35.125 ;
        RECT 171.365 35.065 171.685 35.125 ;
        RECT 172.285 35.065 172.605 35.325 ;
        RECT 176.885 35.265 177.205 35.325 ;
        RECT 177.360 35.265 177.650 35.310 ;
        RECT 176.885 35.125 177.650 35.265 ;
        RECT 176.885 35.065 177.205 35.125 ;
        RECT 177.360 35.080 177.650 35.125 ;
        RECT 185.625 35.065 185.945 35.325 ;
        RECT 187.465 35.265 187.785 35.325 ;
        RECT 188.400 35.265 188.690 35.310 ;
        RECT 197.585 35.265 197.905 35.325 ;
        RECT 187.465 35.125 188.690 35.265 ;
        RECT 187.465 35.065 187.785 35.125 ;
        RECT 188.400 35.080 188.690 35.125 ;
        RECT 188.935 35.125 197.905 35.265 ;
        RECT 167.340 34.925 167.630 34.970 ;
        RECT 170.580 34.925 171.230 34.970 ;
        RECT 172.375 34.925 172.515 35.065 ;
        RECT 167.340 34.785 172.515 34.925 ;
        RECT 180.105 34.925 180.425 34.985 ;
        RECT 181.040 34.925 181.330 34.970 ;
        RECT 180.105 34.785 181.330 34.925 ;
        RECT 167.340 34.740 167.930 34.785 ;
        RECT 170.580 34.740 171.230 34.785 ;
        RECT 167.640 34.425 167.930 34.740 ;
        RECT 180.105 34.725 180.425 34.785 ;
        RECT 181.040 34.740 181.330 34.785 ;
        RECT 181.500 34.925 181.790 34.970 ;
        RECT 187.005 34.925 187.325 34.985 ;
        RECT 181.500 34.785 187.325 34.925 ;
        RECT 181.500 34.740 181.790 34.785 ;
        RECT 187.005 34.725 187.325 34.785 ;
        RECT 168.720 34.585 169.010 34.630 ;
        RECT 172.300 34.585 172.590 34.630 ;
        RECT 174.135 34.585 174.425 34.630 ;
        RECT 168.720 34.445 174.425 34.585 ;
        RECT 168.720 34.400 169.010 34.445 ;
        RECT 172.300 34.400 172.590 34.445 ;
        RECT 174.135 34.400 174.425 34.445 ;
        RECT 174.600 34.585 174.890 34.630 ;
        RECT 175.505 34.585 175.825 34.645 ;
        RECT 174.600 34.445 175.825 34.585 ;
        RECT 174.600 34.400 174.890 34.445 ;
        RECT 175.505 34.385 175.825 34.445 ;
        RECT 176.885 34.385 177.205 34.645 ;
        RECT 178.725 34.585 179.045 34.645 ;
        RECT 188.935 34.585 189.075 35.125 ;
        RECT 197.585 35.065 197.905 35.125 ;
        RECT 205.865 35.265 206.185 35.325 ;
        RECT 205.865 35.125 208.855 35.265 ;
        RECT 205.865 35.065 206.185 35.125 ;
        RECT 193.445 34.970 193.765 34.985 ;
        RECT 189.880 34.925 190.170 34.970 ;
        RECT 193.120 34.925 193.770 34.970 ;
        RECT 189.880 34.785 193.770 34.925 ;
        RECT 189.880 34.740 190.470 34.785 ;
        RECT 193.120 34.740 193.770 34.785 ;
        RECT 201.740 34.925 202.030 34.970 ;
        RECT 202.185 34.925 202.505 34.985 ;
        RECT 201.740 34.785 202.505 34.925 ;
        RECT 201.740 34.740 202.030 34.785 ;
        RECT 178.725 34.445 180.795 34.585 ;
        RECT 178.725 34.385 179.045 34.445 ;
        RECT 173.220 34.245 173.510 34.290 ;
        RECT 178.280 34.245 178.570 34.290 ;
        RECT 179.645 34.245 179.965 34.305 ;
        RECT 180.655 34.290 180.795 34.445 ;
        RECT 184.795 34.445 189.075 34.585 ;
        RECT 184.795 34.290 184.935 34.445 ;
        RECT 190.180 34.425 190.470 34.740 ;
        RECT 193.445 34.725 193.765 34.740 ;
        RECT 202.185 34.725 202.505 34.785 ;
        RECT 204.020 34.925 204.670 34.970 ;
        RECT 207.620 34.925 207.910 34.970 ;
        RECT 208.165 34.925 208.485 34.985 ;
        RECT 204.020 34.785 208.485 34.925 ;
        RECT 208.715 34.925 208.855 35.125 ;
        RECT 209.085 35.065 209.405 35.325 ;
        RECT 215.985 35.265 216.305 35.325 ;
        RECT 218.300 35.265 218.590 35.310 ;
        RECT 225.645 35.265 225.965 35.325 ;
        RECT 234.385 35.265 234.705 35.325 ;
        RECT 215.985 35.125 218.590 35.265 ;
        RECT 215.985 35.065 216.305 35.125 ;
        RECT 218.300 35.080 218.590 35.125 ;
        RECT 221.365 35.125 224.035 35.265 ;
        RECT 216.460 34.925 216.750 34.970 ;
        RECT 208.715 34.785 216.750 34.925 ;
        RECT 204.020 34.740 204.670 34.785 ;
        RECT 207.320 34.740 207.910 34.785 ;
        RECT 191.260 34.585 191.550 34.630 ;
        RECT 194.840 34.585 195.130 34.630 ;
        RECT 196.675 34.585 196.965 34.630 ;
        RECT 191.260 34.445 196.965 34.585 ;
        RECT 191.260 34.400 191.550 34.445 ;
        RECT 194.840 34.400 195.130 34.445 ;
        RECT 196.675 34.400 196.965 34.445 ;
        RECT 200.825 34.585 201.115 34.630 ;
        RECT 202.660 34.585 202.950 34.630 ;
        RECT 206.240 34.585 206.530 34.630 ;
        RECT 200.825 34.445 206.530 34.585 ;
        RECT 200.825 34.400 201.115 34.445 ;
        RECT 202.660 34.400 202.950 34.445 ;
        RECT 206.240 34.400 206.530 34.445 ;
        RECT 207.320 34.425 207.610 34.740 ;
        RECT 208.165 34.725 208.485 34.785 ;
        RECT 216.460 34.740 216.750 34.785 ;
        RECT 216.905 34.925 217.225 34.985 ;
        RECT 219.780 34.925 220.070 34.970 ;
        RECT 221.365 34.925 221.505 35.125 ;
        RECT 223.020 34.925 223.670 34.970 ;
        RECT 223.895 34.925 224.035 35.125 ;
        RECT 225.645 35.125 234.705 35.265 ;
        RECT 225.645 35.065 225.965 35.125 ;
        RECT 234.385 35.065 234.705 35.125 ;
        RECT 234.845 35.265 235.165 35.325 ;
        RECT 238.080 35.265 238.370 35.310 ;
        RECT 234.845 35.125 238.370 35.265 ;
        RECT 234.845 35.065 235.165 35.125 ;
        RECT 238.080 35.080 238.370 35.125 ;
        RECT 249.120 35.265 249.410 35.310 ;
        RECT 253.245 35.265 253.565 35.325 ;
        RECT 263.825 35.265 264.145 35.325 ;
        RECT 249.120 35.125 253.565 35.265 ;
        RECT 249.120 35.080 249.410 35.125 ;
        RECT 253.245 35.065 253.565 35.125 ;
        RECT 255.635 35.125 264.145 35.265 ;
        RECT 228.865 34.925 229.185 34.985 ;
        RECT 216.905 34.785 229.185 34.925 ;
        RECT 216.905 34.725 217.225 34.785 ;
        RECT 219.780 34.740 220.370 34.785 ;
        RECT 223.020 34.740 223.670 34.785 ;
        RECT 216.000 34.585 216.290 34.630 ;
        RECT 216.000 34.445 219.895 34.585 ;
        RECT 216.000 34.400 216.290 34.445 ;
        RECT 173.220 34.105 175.275 34.245 ;
        RECT 173.220 34.060 173.510 34.105 ;
        RECT 175.135 33.950 175.275 34.105 ;
        RECT 178.280 34.105 179.965 34.245 ;
        RECT 178.280 34.060 178.570 34.105 ;
        RECT 179.645 34.045 179.965 34.105 ;
        RECT 180.580 34.245 180.870 34.290 ;
        RECT 184.720 34.245 185.010 34.290 ;
        RECT 180.580 34.105 185.010 34.245 ;
        RECT 180.580 34.060 180.870 34.105 ;
        RECT 184.720 34.060 185.010 34.105 ;
        RECT 185.180 34.060 185.470 34.290 ;
        RECT 195.760 34.245 196.050 34.290 ;
        RECT 187.555 34.105 196.050 34.245 ;
        RECT 168.720 33.905 169.010 33.950 ;
        RECT 171.840 33.905 172.130 33.950 ;
        RECT 173.730 33.905 174.020 33.950 ;
        RECT 168.720 33.765 174.020 33.905 ;
        RECT 168.720 33.720 169.010 33.765 ;
        RECT 171.840 33.720 172.130 33.765 ;
        RECT 173.730 33.720 174.020 33.765 ;
        RECT 175.060 33.720 175.350 33.950 ;
        RECT 183.325 33.365 183.645 33.625 ;
        RECT 185.255 33.565 185.395 34.060 ;
        RECT 187.555 33.950 187.695 34.105 ;
        RECT 195.760 34.060 196.050 34.105 ;
        RECT 197.125 34.245 197.445 34.305 ;
        RECT 199.885 34.245 200.205 34.305 ;
        RECT 200.360 34.245 200.650 34.290 ;
        RECT 197.125 34.105 200.650 34.245 ;
        RECT 197.125 34.045 197.445 34.105 ;
        RECT 199.885 34.045 200.205 34.105 ;
        RECT 200.360 34.060 200.650 34.105 ;
        RECT 210.480 34.060 210.770 34.290 ;
        RECT 210.925 34.245 211.245 34.305 ;
        RECT 217.380 34.245 217.670 34.290 ;
        RECT 210.925 34.105 217.670 34.245 ;
        RECT 219.755 34.245 219.895 34.445 ;
        RECT 220.080 34.425 220.370 34.740 ;
        RECT 228.865 34.725 229.185 34.785 ;
        RECT 230.720 34.925 231.010 34.970 ;
        RECT 232.085 34.925 232.405 34.985 ;
        RECT 230.720 34.785 232.405 34.925 ;
        RECT 230.720 34.740 231.010 34.785 ;
        RECT 232.085 34.725 232.405 34.785 ;
        RECT 233.000 34.925 233.650 34.970 ;
        RECT 236.600 34.925 236.890 34.970 ;
        RECT 237.605 34.925 237.925 34.985 ;
        RECT 233.000 34.785 237.925 34.925 ;
        RECT 233.000 34.740 233.650 34.785 ;
        RECT 236.300 34.740 236.890 34.785 ;
        RECT 221.160 34.585 221.450 34.630 ;
        RECT 224.740 34.585 225.030 34.630 ;
        RECT 226.575 34.585 226.865 34.630 ;
        RECT 221.160 34.445 226.865 34.585 ;
        RECT 221.160 34.400 221.450 34.445 ;
        RECT 224.740 34.400 225.030 34.445 ;
        RECT 226.575 34.400 226.865 34.445 ;
        RECT 229.805 34.585 230.095 34.630 ;
        RECT 231.640 34.585 231.930 34.630 ;
        RECT 235.220 34.585 235.510 34.630 ;
        RECT 229.805 34.445 235.510 34.585 ;
        RECT 229.805 34.400 230.095 34.445 ;
        RECT 231.640 34.400 231.930 34.445 ;
        RECT 235.220 34.400 235.510 34.445 ;
        RECT 236.300 34.425 236.590 34.740 ;
        RECT 237.605 34.725 237.925 34.785 ;
        RECT 241.760 34.925 242.050 34.970 ;
        RECT 243.125 34.925 243.445 34.985 ;
        RECT 241.760 34.785 243.445 34.925 ;
        RECT 241.760 34.740 242.050 34.785 ;
        RECT 243.125 34.725 243.445 34.785 ;
        RECT 244.040 34.925 244.690 34.970 ;
        RECT 244.965 34.925 245.285 34.985 ;
        RECT 247.640 34.925 247.930 34.970 ;
        RECT 244.040 34.785 247.930 34.925 ;
        RECT 244.040 34.740 244.690 34.785 ;
        RECT 244.965 34.725 245.285 34.785 ;
        RECT 247.340 34.740 247.930 34.785 ;
        RECT 240.365 34.385 240.685 34.645 ;
        RECT 240.845 34.585 241.135 34.630 ;
        RECT 242.680 34.585 242.970 34.630 ;
        RECT 246.260 34.585 246.550 34.630 ;
        RECT 240.845 34.445 246.550 34.585 ;
        RECT 240.845 34.400 241.135 34.445 ;
        RECT 242.680 34.400 242.970 34.445 ;
        RECT 246.260 34.400 246.550 34.445 ;
        RECT 247.340 34.425 247.630 34.740 ;
        RECT 220.585 34.245 220.905 34.305 ;
        RECT 219.755 34.105 220.905 34.245 ;
        RECT 187.480 33.720 187.770 33.950 ;
        RECT 191.260 33.905 191.550 33.950 ;
        RECT 194.380 33.905 194.670 33.950 ;
        RECT 196.270 33.905 196.560 33.950 ;
        RECT 191.260 33.765 196.560 33.905 ;
        RECT 191.260 33.720 191.550 33.765 ;
        RECT 194.380 33.720 194.670 33.765 ;
        RECT 196.270 33.720 196.560 33.765 ;
        RECT 201.230 33.905 201.520 33.950 ;
        RECT 203.120 33.905 203.410 33.950 ;
        RECT 206.240 33.905 206.530 33.950 ;
        RECT 201.230 33.765 206.530 33.905 ;
        RECT 210.555 33.905 210.695 34.060 ;
        RECT 210.925 34.045 211.245 34.105 ;
        RECT 217.380 34.060 217.670 34.105 ;
        RECT 214.160 33.905 214.450 33.950 ;
        RECT 210.555 33.765 214.450 33.905 ;
        RECT 201.230 33.720 201.520 33.765 ;
        RECT 203.120 33.720 203.410 33.765 ;
        RECT 206.240 33.720 206.530 33.765 ;
        RECT 214.160 33.720 214.450 33.765 ;
        RECT 193.905 33.565 194.225 33.625 ;
        RECT 185.255 33.425 194.225 33.565 ;
        RECT 193.905 33.365 194.225 33.425 ;
        RECT 213.225 33.365 213.545 33.625 ;
        RECT 217.455 33.565 217.595 34.060 ;
        RECT 220.585 34.045 220.905 34.105 ;
        RECT 225.645 34.045 225.965 34.305 ;
        RECT 227.025 34.245 227.345 34.305 ;
        RECT 229.340 34.245 229.630 34.290 ;
        RECT 227.025 34.105 229.630 34.245 ;
        RECT 240.455 34.245 240.595 34.385 ;
        RECT 255.635 34.290 255.775 35.125 ;
        RECT 263.825 35.065 264.145 35.125 ;
        RECT 281.765 35.265 282.085 35.325 ;
        RECT 299.720 35.265 300.010 35.310 ;
        RECT 281.765 35.125 300.010 35.265 ;
        RECT 281.765 35.065 282.085 35.125 ;
        RECT 299.720 35.080 300.010 35.125 ;
        RECT 256.925 34.725 257.245 34.985 ;
        RECT 257.385 34.925 257.705 34.985 ;
        RECT 259.220 34.925 259.870 34.970 ;
        RECT 262.820 34.925 263.110 34.970 ;
        RECT 257.385 34.785 263.110 34.925 ;
        RECT 257.385 34.725 257.705 34.785 ;
        RECT 259.220 34.740 259.870 34.785 ;
        RECT 262.520 34.740 263.110 34.785 ;
        RECT 301.200 34.925 301.490 34.970 ;
        RECT 303.385 34.925 303.705 34.985 ;
        RECT 304.440 34.925 305.090 34.970 ;
        RECT 301.200 34.785 305.090 34.925 ;
        RECT 301.200 34.740 301.790 34.785 ;
        RECT 256.025 34.585 256.315 34.630 ;
        RECT 257.860 34.585 258.150 34.630 ;
        RECT 261.440 34.585 261.730 34.630 ;
        RECT 256.025 34.445 261.730 34.585 ;
        RECT 256.025 34.400 256.315 34.445 ;
        RECT 257.860 34.400 258.150 34.445 ;
        RECT 261.440 34.400 261.730 34.445 ;
        RECT 262.520 34.425 262.810 34.740 ;
        RECT 265.205 34.585 265.525 34.645 ;
        RECT 263.915 34.445 265.525 34.585 ;
        RECT 255.560 34.245 255.850 34.290 ;
        RECT 240.455 34.105 255.850 34.245 ;
        RECT 227.025 34.045 227.345 34.105 ;
        RECT 229.340 34.060 229.630 34.105 ;
        RECT 255.560 34.060 255.850 34.105 ;
        RECT 257.385 34.245 257.705 34.305 ;
        RECT 263.915 34.245 264.055 34.445 ;
        RECT 265.205 34.385 265.525 34.445 ;
        RECT 266.600 34.585 266.890 34.630 ;
        RECT 268.425 34.585 268.745 34.645 ;
        RECT 266.600 34.445 268.745 34.585 ;
        RECT 266.600 34.400 266.890 34.445 ;
        RECT 268.425 34.385 268.745 34.445 ;
        RECT 301.500 34.425 301.790 34.740 ;
        RECT 303.385 34.725 303.705 34.785 ;
        RECT 304.440 34.740 305.090 34.785 ;
        RECT 305.685 34.925 306.005 34.985 ;
        RECT 305.685 34.785 308.675 34.925 ;
        RECT 305.685 34.725 306.005 34.785 ;
        RECT 308.535 34.630 308.675 34.785 ;
        RECT 302.580 34.585 302.870 34.630 ;
        RECT 306.160 34.585 306.450 34.630 ;
        RECT 307.995 34.585 308.285 34.630 ;
        RECT 302.580 34.445 308.285 34.585 ;
        RECT 302.580 34.400 302.870 34.445 ;
        RECT 306.160 34.400 306.450 34.445 ;
        RECT 307.995 34.400 308.285 34.445 ;
        RECT 308.460 34.400 308.750 34.630 ;
        RECT 257.385 34.105 264.055 34.245 ;
        RECT 264.300 34.245 264.590 34.290 ;
        RECT 267.505 34.245 267.825 34.305 ;
        RECT 264.300 34.105 267.825 34.245 ;
        RECT 257.385 34.045 257.705 34.105 ;
        RECT 264.300 34.060 264.590 34.105 ;
        RECT 267.505 34.045 267.825 34.105 ;
        RECT 307.065 34.045 307.385 34.305 ;
        RECT 221.160 33.905 221.450 33.950 ;
        RECT 224.280 33.905 224.570 33.950 ;
        RECT 226.170 33.905 226.460 33.950 ;
        RECT 221.160 33.765 226.460 33.905 ;
        RECT 221.160 33.720 221.450 33.765 ;
        RECT 224.280 33.720 224.570 33.765 ;
        RECT 226.170 33.720 226.460 33.765 ;
        RECT 230.210 33.905 230.500 33.950 ;
        RECT 232.100 33.905 232.390 33.950 ;
        RECT 235.220 33.905 235.510 33.950 ;
        RECT 230.210 33.765 235.510 33.905 ;
        RECT 230.210 33.720 230.500 33.765 ;
        RECT 232.100 33.720 232.390 33.765 ;
        RECT 235.220 33.720 235.510 33.765 ;
        RECT 241.250 33.905 241.540 33.950 ;
        RECT 243.140 33.905 243.430 33.950 ;
        RECT 246.260 33.905 246.550 33.950 ;
        RECT 241.250 33.765 246.550 33.905 ;
        RECT 241.250 33.720 241.540 33.765 ;
        RECT 243.140 33.720 243.430 33.765 ;
        RECT 246.260 33.720 246.550 33.765 ;
        RECT 256.430 33.905 256.720 33.950 ;
        RECT 258.320 33.905 258.610 33.950 ;
        RECT 261.440 33.905 261.730 33.950 ;
        RECT 256.430 33.765 261.730 33.905 ;
        RECT 256.430 33.720 256.720 33.765 ;
        RECT 258.320 33.720 258.610 33.765 ;
        RECT 261.440 33.720 261.730 33.765 ;
        RECT 302.580 33.905 302.870 33.950 ;
        RECT 305.700 33.905 305.990 33.950 ;
        RECT 307.590 33.905 307.880 33.950 ;
        RECT 302.580 33.765 307.880 33.905 ;
        RECT 302.580 33.720 302.870 33.765 ;
        RECT 305.700 33.720 305.990 33.765 ;
        RECT 307.590 33.720 307.880 33.765 ;
        RECT 228.405 33.565 228.725 33.625 ;
        RECT 217.455 33.425 228.725 33.565 ;
        RECT 228.405 33.365 228.725 33.425 ;
        RECT 259.685 33.565 260.005 33.625 ;
        RECT 260.605 33.565 260.925 33.625 ;
        RECT 265.680 33.565 265.970 33.610 ;
        RECT 259.685 33.425 265.970 33.565 ;
        RECT 259.685 33.365 260.005 33.425 ;
        RECT 260.605 33.365 260.925 33.425 ;
        RECT 265.680 33.380 265.970 33.425 ;
        RECT 162.095 32.745 311.135 33.225 ;
        RECT 167.175 32.545 167.465 32.590 ;
        RECT 175.520 32.545 175.810 32.590 ;
        RECT 167.175 32.405 175.810 32.545 ;
        RECT 167.175 32.360 167.465 32.405 ;
        RECT 175.520 32.360 175.810 32.405 ;
        RECT 181.960 32.545 182.250 32.590 ;
        RECT 182.865 32.545 183.185 32.605 ;
        RECT 205.865 32.545 206.185 32.605 ;
        RECT 206.340 32.545 206.630 32.590 ;
        RECT 210.925 32.545 211.245 32.605 ;
        RECT 181.960 32.405 183.185 32.545 ;
        RECT 181.960 32.360 182.250 32.405 ;
        RECT 182.865 32.345 183.185 32.405 ;
        RECT 183.415 32.405 194.595 32.545 ;
        RECT 166.730 32.205 167.020 32.250 ;
        RECT 168.620 32.205 168.910 32.250 ;
        RECT 171.740 32.205 172.030 32.250 ;
        RECT 166.730 32.065 172.030 32.205 ;
        RECT 166.730 32.020 167.020 32.065 ;
        RECT 168.620 32.020 168.910 32.065 ;
        RECT 171.740 32.020 172.030 32.065 ;
        RECT 174.600 32.205 174.890 32.250 ;
        RECT 175.045 32.205 175.365 32.265 ;
        RECT 179.645 32.205 179.965 32.265 ;
        RECT 183.415 32.205 183.555 32.405 ;
        RECT 174.600 32.065 175.365 32.205 ;
        RECT 174.600 32.020 174.890 32.065 ;
        RECT 175.045 32.005 175.365 32.065 ;
        RECT 178.815 32.065 183.555 32.205 ;
        RECT 184.820 32.205 185.110 32.250 ;
        RECT 187.940 32.205 188.230 32.250 ;
        RECT 189.830 32.205 190.120 32.250 ;
        RECT 184.820 32.065 190.120 32.205 ;
        RECT 165.845 31.665 166.165 31.925 ;
        RECT 176.885 31.865 177.205 31.925 ;
        RECT 178.815 31.910 178.955 32.065 ;
        RECT 179.645 32.005 179.965 32.065 ;
        RECT 184.820 32.020 185.110 32.065 ;
        RECT 187.940 32.020 188.230 32.065 ;
        RECT 189.830 32.020 190.120 32.065 ;
        RECT 194.455 32.205 194.595 32.405 ;
        RECT 205.865 32.405 206.630 32.545 ;
        RECT 205.865 32.345 206.185 32.405 ;
        RECT 206.340 32.360 206.630 32.405 ;
        RECT 206.875 32.405 211.245 32.545 ;
        RECT 206.875 32.205 207.015 32.405 ;
        RECT 210.925 32.345 211.245 32.405 ;
        RECT 213.225 32.545 213.545 32.605 ;
        RECT 213.760 32.545 214.050 32.590 ;
        RECT 213.225 32.405 214.050 32.545 ;
        RECT 213.225 32.345 213.545 32.405 ;
        RECT 213.760 32.360 214.050 32.405 ;
        RECT 220.585 32.545 220.905 32.605 ;
        RECT 222.440 32.545 222.730 32.590 ;
        RECT 225.645 32.545 225.965 32.605 ;
        RECT 220.585 32.405 221.505 32.545 ;
        RECT 220.585 32.345 220.905 32.405 ;
        RECT 194.455 32.065 207.015 32.205 ;
        RECT 209.200 32.205 209.490 32.250 ;
        RECT 212.320 32.205 212.610 32.250 ;
        RECT 214.210 32.205 214.500 32.250 ;
        RECT 209.200 32.065 214.500 32.205 ;
        RECT 194.455 31.910 194.595 32.065 ;
        RECT 204.575 31.910 204.715 32.065 ;
        RECT 209.200 32.020 209.490 32.065 ;
        RECT 212.320 32.020 212.610 32.065 ;
        RECT 214.210 32.020 214.500 32.065 ;
        RECT 177.820 31.865 178.110 31.910 ;
        RECT 176.885 31.725 178.110 31.865 ;
        RECT 176.885 31.665 177.205 31.725 ;
        RECT 177.820 31.680 178.110 31.725 ;
        RECT 178.740 31.680 179.030 31.910 ;
        RECT 193.460 31.865 193.750 31.910 ;
        RECT 182.955 31.725 193.750 31.865 ;
        RECT 166.325 31.525 166.615 31.570 ;
        RECT 168.160 31.525 168.450 31.570 ;
        RECT 171.740 31.525 172.030 31.570 ;
        RECT 166.325 31.385 172.030 31.525 ;
        RECT 166.325 31.340 166.615 31.385 ;
        RECT 168.160 31.340 168.450 31.385 ;
        RECT 171.740 31.340 172.030 31.385 ;
        RECT 172.820 31.230 173.110 31.545 ;
        RECT 177.360 31.525 177.650 31.570 ;
        RECT 179.645 31.525 179.965 31.585 ;
        RECT 182.955 31.525 183.095 31.725 ;
        RECT 193.460 31.680 193.750 31.725 ;
        RECT 194.380 31.680 194.670 31.910 ;
        RECT 204.500 31.680 204.790 31.910 ;
        RECT 215.080 31.865 215.370 31.910 ;
        RECT 221.365 31.865 221.505 32.405 ;
        RECT 222.440 32.405 225.965 32.545 ;
        RECT 222.440 32.360 222.730 32.405 ;
        RECT 225.645 32.345 225.965 32.405 ;
        RECT 226.105 32.545 226.425 32.605 ;
        RECT 228.325 32.545 228.615 32.590 ;
        RECT 226.105 32.405 228.615 32.545 ;
        RECT 226.105 32.345 226.425 32.405 ;
        RECT 228.325 32.360 228.615 32.405 ;
        RECT 234.385 32.545 234.705 32.605 ;
        RECT 243.140 32.545 243.430 32.590 ;
        RECT 249.105 32.545 249.425 32.605 ;
        RECT 234.385 32.405 249.425 32.545 ;
        RECT 234.385 32.345 234.705 32.405 ;
        RECT 243.140 32.360 243.430 32.405 ;
        RECT 249.105 32.345 249.425 32.405 ;
        RECT 260.145 32.545 260.465 32.605 ;
        RECT 260.620 32.545 260.910 32.590 ;
        RECT 260.145 32.405 260.910 32.545 ;
        RECT 260.145 32.345 260.465 32.405 ;
        RECT 260.620 32.360 260.910 32.405 ;
        RECT 227.910 32.205 228.200 32.250 ;
        RECT 229.800 32.205 230.090 32.250 ;
        RECT 232.920 32.205 233.210 32.250 ;
        RECT 264.745 32.205 265.065 32.265 ;
        RECT 227.910 32.065 233.210 32.205 ;
        RECT 227.910 32.020 228.200 32.065 ;
        RECT 229.800 32.020 230.090 32.065 ;
        RECT 232.920 32.020 233.210 32.065 ;
        RECT 255.635 32.065 265.065 32.205 ;
        RECT 224.740 31.865 225.030 31.910 ;
        RECT 215.080 31.725 218.515 31.865 ;
        RECT 221.365 31.725 225.030 31.865 ;
        RECT 215.080 31.680 215.370 31.725 ;
        RECT 177.360 31.385 183.095 31.525 ;
        RECT 177.360 31.340 177.650 31.385 ;
        RECT 179.645 31.325 179.965 31.385 ;
        RECT 183.740 31.230 184.030 31.545 ;
        RECT 184.820 31.525 185.110 31.570 ;
        RECT 188.400 31.525 188.690 31.570 ;
        RECT 190.235 31.525 190.525 31.570 ;
        RECT 184.820 31.385 190.525 31.525 ;
        RECT 184.820 31.340 185.110 31.385 ;
        RECT 188.400 31.340 188.690 31.385 ;
        RECT 190.235 31.340 190.525 31.385 ;
        RECT 190.700 31.525 190.990 31.570 ;
        RECT 197.125 31.525 197.445 31.585 ;
        RECT 203.580 31.525 203.870 31.570 ;
        RECT 208.165 31.545 208.485 31.585 ;
        RECT 190.700 31.385 197.445 31.525 ;
        RECT 190.700 31.340 190.990 31.385 ;
        RECT 197.125 31.325 197.445 31.385 ;
        RECT 197.675 31.385 203.870 31.525 ;
        RECT 169.520 31.185 170.170 31.230 ;
        RECT 172.820 31.185 173.410 31.230 ;
        RECT 183.440 31.185 184.030 31.230 ;
        RECT 186.545 31.230 186.865 31.245 ;
        RECT 186.545 31.185 187.330 31.230 ;
        RECT 169.520 31.045 183.095 31.185 ;
        RECT 169.520 31.000 170.170 31.045 ;
        RECT 173.120 31.000 173.410 31.045 ;
        RECT 182.955 30.845 183.095 31.045 ;
        RECT 183.440 31.045 187.330 31.185 ;
        RECT 183.440 31.000 183.730 31.045 ;
        RECT 186.545 31.000 187.330 31.045 ;
        RECT 187.925 31.185 188.245 31.245 ;
        RECT 189.320 31.185 189.610 31.230 ;
        RECT 187.925 31.045 189.610 31.185 ;
        RECT 186.545 30.985 186.865 31.000 ;
        RECT 187.925 30.985 188.245 31.045 ;
        RECT 189.320 31.000 189.610 31.045 ;
        RECT 193.000 31.185 193.290 31.230 ;
        RECT 193.905 31.185 194.225 31.245 ;
        RECT 197.675 31.185 197.815 31.385 ;
        RECT 203.580 31.340 203.870 31.385 ;
        RECT 208.120 31.325 208.485 31.545 ;
        RECT 209.200 31.525 209.490 31.570 ;
        RECT 212.780 31.525 213.070 31.570 ;
        RECT 214.615 31.525 214.905 31.570 ;
        RECT 209.200 31.385 214.905 31.525 ;
        RECT 209.200 31.340 209.490 31.385 ;
        RECT 212.780 31.340 213.070 31.385 ;
        RECT 214.615 31.340 214.905 31.385 ;
        RECT 215.985 31.525 216.305 31.585 ;
        RECT 217.380 31.525 217.670 31.570 ;
        RECT 215.985 31.385 217.670 31.525 ;
        RECT 218.375 31.525 218.515 31.725 ;
        RECT 224.740 31.680 225.030 31.725 ;
        RECT 225.660 31.865 225.950 31.910 ;
        RECT 228.405 31.865 228.725 31.925 ;
        RECT 225.660 31.725 228.725 31.865 ;
        RECT 225.660 31.680 225.950 31.725 ;
        RECT 228.405 31.665 228.725 31.725 ;
        RECT 228.865 31.865 229.185 31.925 ;
        RECT 235.780 31.865 236.070 31.910 ;
        RECT 239.000 31.865 239.290 31.910 ;
        RECT 255.635 31.865 255.775 32.065 ;
        RECT 264.745 32.005 265.065 32.065 ;
        RECT 228.865 31.725 234.615 31.865 ;
        RECT 228.865 31.665 229.185 31.725 ;
        RECT 227.025 31.525 227.345 31.585 ;
        RECT 218.375 31.385 227.345 31.525 ;
        RECT 215.985 31.325 216.305 31.385 ;
        RECT 217.380 31.340 217.670 31.385 ;
        RECT 227.025 31.325 227.345 31.385 ;
        RECT 227.505 31.525 227.795 31.570 ;
        RECT 229.340 31.525 229.630 31.570 ;
        RECT 232.920 31.525 233.210 31.570 ;
        RECT 227.505 31.385 233.210 31.525 ;
        RECT 227.505 31.340 227.795 31.385 ;
        RECT 229.340 31.340 229.630 31.385 ;
        RECT 232.920 31.340 233.210 31.385 ;
        RECT 193.000 31.045 197.815 31.185 ;
        RECT 198.505 31.185 198.825 31.245 ;
        RECT 199.900 31.185 200.190 31.230 ;
        RECT 198.505 31.045 200.190 31.185 ;
        RECT 193.000 31.000 193.290 31.045 ;
        RECT 193.905 30.985 194.225 31.045 ;
        RECT 198.505 30.985 198.825 31.045 ;
        RECT 199.900 31.000 200.190 31.045 ;
        RECT 203.120 31.185 203.410 31.230 ;
        RECT 204.945 31.185 205.265 31.245 ;
        RECT 208.120 31.230 208.410 31.325 ;
        RECT 234.000 31.230 234.290 31.545 ;
        RECT 234.475 31.230 234.615 31.725 ;
        RECT 235.780 31.725 239.290 31.865 ;
        RECT 235.780 31.680 236.070 31.725 ;
        RECT 239.000 31.680 239.290 31.725 ;
        RECT 245.515 31.725 255.775 31.865 ;
        RECT 256.005 31.865 256.325 31.925 ;
        RECT 256.005 31.725 261.295 31.865 ;
        RECT 245.515 31.585 245.655 31.725 ;
        RECT 256.005 31.665 256.325 31.725 ;
        RECT 235.305 31.525 235.625 31.585 ;
        RECT 236.240 31.525 236.530 31.570 ;
        RECT 235.305 31.385 236.530 31.525 ;
        RECT 235.305 31.325 235.625 31.385 ;
        RECT 236.240 31.340 236.530 31.385 ;
        RECT 243.600 31.525 243.890 31.570 ;
        RECT 245.425 31.525 245.745 31.585 ;
        RECT 243.600 31.385 245.745 31.525 ;
        RECT 243.600 31.340 243.890 31.385 ;
        RECT 245.425 31.325 245.745 31.385 ;
        RECT 260.160 31.525 260.450 31.570 ;
        RECT 260.605 31.525 260.925 31.585 ;
        RECT 261.155 31.570 261.295 31.725 ;
        RECT 260.160 31.385 260.925 31.525 ;
        RECT 260.160 31.340 260.450 31.385 ;
        RECT 260.605 31.325 260.925 31.385 ;
        RECT 261.080 31.340 261.370 31.570 ;
        RECT 203.120 31.045 205.265 31.185 ;
        RECT 203.120 31.000 203.410 31.045 ;
        RECT 204.945 30.985 205.265 31.045 ;
        RECT 207.820 31.185 208.410 31.230 ;
        RECT 211.060 31.185 211.710 31.230 ;
        RECT 207.820 31.045 211.710 31.185 ;
        RECT 207.820 31.000 208.110 31.045 ;
        RECT 211.060 31.000 211.710 31.045 ;
        RECT 230.700 31.185 231.350 31.230 ;
        RECT 234.000 31.185 234.615 31.230 ;
        RECT 237.605 31.185 237.925 31.245 ;
        RECT 239.920 31.185 240.210 31.230 ;
        RECT 230.700 31.045 240.210 31.185 ;
        RECT 230.700 31.000 231.350 31.045 ;
        RECT 234.300 31.000 234.590 31.045 ;
        RECT 237.605 30.985 237.925 31.045 ;
        RECT 239.920 31.000 240.210 31.045 ;
        RECT 241.745 31.185 242.065 31.245 ;
        RECT 254.625 31.185 254.945 31.245 ;
        RECT 241.745 31.045 254.945 31.185 ;
        RECT 241.745 30.985 242.065 31.045 ;
        RECT 254.625 30.985 254.945 31.045 ;
        RECT 184.245 30.845 184.565 30.905 ;
        RECT 182.955 30.705 184.565 30.845 ;
        RECT 184.245 30.645 184.565 30.705 ;
        RECT 186.085 30.845 186.405 30.905 ;
        RECT 191.160 30.845 191.450 30.890 ;
        RECT 186.085 30.705 191.450 30.845 ;
        RECT 186.085 30.645 186.405 30.705 ;
        RECT 191.160 30.660 191.450 30.705 ;
        RECT 193.445 30.845 193.765 30.905 ;
        RECT 199.425 30.845 199.745 30.905 ;
        RECT 193.445 30.705 199.745 30.845 ;
        RECT 193.445 30.645 193.765 30.705 ;
        RECT 199.425 30.645 199.745 30.705 ;
        RECT 201.280 30.845 201.570 30.890 ;
        RECT 202.645 30.845 202.965 30.905 ;
        RECT 201.280 30.705 202.965 30.845 ;
        RECT 201.280 30.660 201.570 30.705 ;
        RECT 202.645 30.645 202.965 30.705 ;
        RECT 224.280 30.845 224.570 30.890 ;
        RECT 235.765 30.845 236.085 30.905 ;
        RECT 224.280 30.705 236.085 30.845 ;
        RECT 224.280 30.660 224.570 30.705 ;
        RECT 235.765 30.645 236.085 30.705 ;
        RECT 162.095 30.025 311.135 30.505 ;
        RECT 176.885 29.825 177.205 29.885 ;
        RECT 178.280 29.825 178.570 29.870 ;
        RECT 176.885 29.685 178.570 29.825 ;
        RECT 176.885 29.625 177.205 29.685 ;
        RECT 178.280 29.640 178.570 29.685 ;
        RECT 184.245 29.825 184.565 29.885 ;
        RECT 186.545 29.825 186.865 29.885 ;
        RECT 193.445 29.825 193.765 29.885 ;
        RECT 184.245 29.685 193.765 29.825 ;
        RECT 184.245 29.625 184.565 29.685 ;
        RECT 186.545 29.625 186.865 29.685 ;
        RECT 193.445 29.625 193.765 29.685 ;
        RECT 195.285 29.825 195.605 29.885 ;
        RECT 195.760 29.825 196.050 29.870 ;
        RECT 195.285 29.685 196.050 29.825 ;
        RECT 195.285 29.625 195.605 29.685 ;
        RECT 195.760 29.640 196.050 29.685 ;
        RECT 199.885 29.825 200.205 29.885 ;
        RECT 199.885 29.685 204.715 29.825 ;
        RECT 199.885 29.625 200.205 29.685 ;
        RECT 180.220 29.485 180.510 29.530 ;
        RECT 183.460 29.485 184.110 29.530 ;
        RECT 184.335 29.485 184.475 29.625 ;
        RECT 180.220 29.345 184.475 29.485 ;
        RECT 180.220 29.300 180.810 29.345 ;
        RECT 183.460 29.300 184.110 29.345 ;
        RECT 164.940 29.145 165.230 29.190 ;
        RECT 170.905 29.145 171.225 29.205 ;
        RECT 164.940 29.005 171.225 29.145 ;
        RECT 164.940 28.960 165.230 29.005 ;
        RECT 170.905 28.945 171.225 29.005 ;
        RECT 175.045 28.945 175.365 29.205 ;
        RECT 180.520 28.985 180.810 29.300 ;
        RECT 186.085 29.285 186.405 29.545 ;
        RECT 197.240 29.485 197.530 29.530 ;
        RECT 199.425 29.485 199.745 29.545 ;
        RECT 200.480 29.485 201.130 29.530 ;
        RECT 197.240 29.345 201.130 29.485 ;
        RECT 197.240 29.300 197.830 29.345 ;
        RECT 181.600 29.145 181.890 29.190 ;
        RECT 185.180 29.145 185.470 29.190 ;
        RECT 187.015 29.145 187.305 29.190 ;
        RECT 181.600 29.005 187.305 29.145 ;
        RECT 181.600 28.960 181.890 29.005 ;
        RECT 185.180 28.960 185.470 29.005 ;
        RECT 187.015 28.960 187.305 29.005 ;
        RECT 187.480 29.145 187.770 29.190 ;
        RECT 189.305 29.145 189.625 29.205 ;
        RECT 187.480 29.005 189.625 29.145 ;
        RECT 187.480 28.960 187.770 29.005 ;
        RECT 189.305 28.945 189.625 29.005 ;
        RECT 197.540 28.985 197.830 29.300 ;
        RECT 199.425 29.285 199.745 29.345 ;
        RECT 200.480 29.300 201.130 29.345 ;
        RECT 202.645 29.485 202.965 29.545 ;
        RECT 203.120 29.485 203.410 29.530 ;
        RECT 202.645 29.345 203.410 29.485 ;
        RECT 202.645 29.285 202.965 29.345 ;
        RECT 203.120 29.300 203.410 29.345 ;
        RECT 204.575 29.190 204.715 29.685 ;
        RECT 204.945 29.625 205.265 29.885 ;
        RECT 231.640 29.825 231.930 29.870 ;
        RECT 235.765 29.825 236.085 29.885 ;
        RECT 231.640 29.685 236.085 29.825 ;
        RECT 231.640 29.640 231.930 29.685 ;
        RECT 235.765 29.625 236.085 29.685 ;
        RECT 198.620 29.145 198.910 29.190 ;
        RECT 202.200 29.145 202.490 29.190 ;
        RECT 204.035 29.145 204.325 29.190 ;
        RECT 198.620 29.005 204.325 29.145 ;
        RECT 198.620 28.960 198.910 29.005 ;
        RECT 202.200 28.960 202.490 29.005 ;
        RECT 204.035 28.960 204.325 29.005 ;
        RECT 204.500 28.960 204.790 29.190 ;
        RECT 205.865 29.145 206.185 29.205 ;
        RECT 207.720 29.145 208.010 29.190 ;
        RECT 205.865 29.005 208.010 29.145 ;
        RECT 205.865 28.945 206.185 29.005 ;
        RECT 207.720 28.960 208.010 29.005 ;
        RECT 234.845 28.945 235.165 29.205 ;
        RECT 178.740 28.805 179.030 28.850 ;
        RECT 180.105 28.805 180.425 28.865 ;
        RECT 178.740 28.665 180.425 28.805 ;
        RECT 178.740 28.620 179.030 28.665 ;
        RECT 180.105 28.605 180.425 28.665 ;
        RECT 181.600 28.465 181.890 28.510 ;
        RECT 184.720 28.465 185.010 28.510 ;
        RECT 186.610 28.465 186.900 28.510 ;
        RECT 181.600 28.325 186.900 28.465 ;
        RECT 181.600 28.280 181.890 28.325 ;
        RECT 184.720 28.280 185.010 28.325 ;
        RECT 186.610 28.280 186.900 28.325 ;
        RECT 198.620 28.465 198.910 28.510 ;
        RECT 201.740 28.465 202.030 28.510 ;
        RECT 203.630 28.465 203.920 28.510 ;
        RECT 198.620 28.325 203.920 28.465 ;
        RECT 198.620 28.280 198.910 28.325 ;
        RECT 201.740 28.280 202.030 28.325 ;
        RECT 203.630 28.280 203.920 28.325 ;
        RECT 164.005 27.925 164.325 28.185 ;
        RECT 162.095 27.305 311.135 27.785 ;
        RECT 178.280 27.105 178.570 27.150 ;
        RECT 179.645 27.105 179.965 27.165 ;
        RECT 178.280 26.965 179.965 27.105 ;
        RECT 178.280 26.920 178.570 26.965 ;
        RECT 179.645 26.905 179.965 26.965 ;
        RECT 186.560 27.105 186.850 27.150 ;
        RECT 187.925 27.105 188.245 27.165 ;
        RECT 186.560 26.965 188.245 27.105 ;
        RECT 186.560 26.920 186.850 26.965 ;
        RECT 187.925 26.905 188.245 26.965 ;
        RECT 180.105 26.425 180.425 26.485 ;
        RECT 181.040 26.425 181.330 26.470 ;
        RECT 180.105 26.285 181.330 26.425 ;
        RECT 180.105 26.225 180.425 26.285 ;
        RECT 181.040 26.240 181.330 26.285 ;
        RECT 183.325 26.225 183.645 26.485 ;
        RECT 162.095 24.585 311.135 25.065 ;
        RECT 162.095 21.865 311.135 22.345 ;
        RECT 162.095 19.145 311.135 19.625 ;
        RECT 135.120 14.050 138.400 18.845 ;
        RECT 146.290 14.050 155.900 18.845 ;
        RECT 162.095 16.425 311.135 16.905 ;
        RECT 135.120 4.900 155.900 14.050 ;
        RECT 162.095 13.705 311.135 14.185 ;
        RECT 4.100 4.100 155.900 4.900 ;
      LAYER met2 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.410 213.985 225.710 ;
        RECT 64.710 225.310 65.510 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 67.470 224.810 204.325 225.110 ;
        RECT 67.470 224.710 68.270 224.810 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.210 194.665 224.510 ;
        RECT 70.230 224.110 71.030 224.210 ;
        RECT 72.990 223.610 185.005 223.910 ;
        RECT 72.990 223.510 73.790 223.610 ;
        RECT 75.700 223.010 175.345 223.310 ;
        RECT 75.700 222.910 76.500 223.010 ;
        RECT 78.545 222.410 165.685 222.710 ;
        RECT 78.545 222.310 79.345 222.410 ;
        RECT 83.980 221.810 164.500 222.110 ;
        RECT 83.980 221.710 84.780 221.810 ;
        RECT 86.740 221.210 163.500 221.510 ;
        RECT 164.100 221.310 164.500 221.810 ;
        RECT 86.740 221.110 87.540 221.210 ;
        RECT 92.260 220.610 162.500 220.910 ;
        RECT 163.100 220.710 163.500 221.210 ;
        RECT 92.260 220.510 93.060 220.610 ;
        RECT 162.100 220.110 162.500 220.610 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.495 208.765 51.905 210.765 ;
        RECT 9.495 205.765 45.165 207.765 ;
        RECT 51.315 207.460 51.905 208.765 ;
        RECT 9.495 202.765 48.270 204.765 ;
        RECT 9.495 198.745 48.270 200.745 ;
        RECT 9.495 195.745 45.165 197.745 ;
        RECT 9.495 192.745 46.670 194.745 ;
        RECT 9.495 187.420 15.245 188.980 ;
        RECT 16.515 188.295 45.165 190.295 ;
        RECT 52.860 188.465 54.245 190.570 ;
        RECT 16.515 184.775 56.920 186.775 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.495 182.570 15.245 184.130 ;
        RECT 16.515 181.255 46.670 183.255 ;
        RECT 5.910 176.050 7.510 179.250 ;
        RECT 57.020 178.865 57.820 178.990 ;
        RECT 9.500 177.365 58.420 178.865 ;
        RECT 53.870 176.720 54.670 176.890 ;
        RECT 9.500 175.220 54.670 176.720 ;
        RECT 9.500 172.820 54.670 174.320 ;
        RECT 53.870 172.640 54.670 172.820 ;
        RECT 52.220 171.920 53.020 172.040 ;
        RECT 9.500 170.420 53.020 171.920 ;
        RECT 63.470 170.855 65.220 217.105 ;
        RECT 66.220 170.855 67.970 217.105 ;
        RECT 68.970 170.855 70.720 217.105 ;
        RECT 71.720 170.855 73.470 217.105 ;
        RECT 74.470 170.855 76.220 217.105 ;
        RECT 77.220 170.855 78.970 217.105 ;
        RECT 79.970 170.115 81.970 217.845 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 109.240 219.705 111.675 220.105 ;
        RECT 113.270 219.705 115.705 220.105 ;
        RECT 117.300 219.705 119.735 220.105 ;
        RECT 121.330 219.705 123.765 220.105 ;
        RECT 125.360 219.705 127.795 220.105 ;
        RECT 129.390 219.705 131.825 220.105 ;
        RECT 133.420 219.705 135.855 220.105 ;
        RECT 137.450 219.705 139.885 220.105 ;
        RECT 141.480 219.705 143.915 220.105 ;
        RECT 145.510 219.705 147.945 220.105 ;
        RECT 149.540 219.705 151.975 220.105 ;
        RECT 109.240 217.705 109.640 219.705 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 111.820 217.295 112.220 219.305 ;
        RECT 113.270 217.705 113.670 219.705 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 115.850 217.295 116.250 219.305 ;
        RECT 117.300 217.705 117.700 219.705 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 119.880 217.295 120.280 219.305 ;
        RECT 121.330 217.705 121.730 219.705 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 123.910 217.295 124.310 219.305 ;
        RECT 125.360 217.705 125.760 219.705 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 127.940 217.295 128.340 219.305 ;
        RECT 129.390 217.705 129.790 219.705 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 131.970 217.295 132.370 219.305 ;
        RECT 133.420 217.705 133.820 219.705 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 136.000 217.295 136.400 219.305 ;
        RECT 137.450 217.705 137.850 219.705 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 140.030 217.295 140.430 219.305 ;
        RECT 141.480 217.705 141.880 219.705 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 144.060 217.295 144.460 219.305 ;
        RECT 145.510 217.705 145.910 219.705 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 148.090 217.295 148.490 219.305 ;
        RECT 149.540 217.705 149.940 219.705 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 152.120 217.295 152.520 219.305 ;
        RECT 82.970 170.855 84.720 217.105 ;
        RECT 85.720 170.855 87.470 217.105 ;
        RECT 88.470 170.855 90.220 217.105 ;
        RECT 91.220 170.855 92.970 217.105 ;
        RECT 93.970 170.855 95.720 217.105 ;
        RECT 96.720 170.855 98.470 217.105 ;
        RECT 109.785 216.895 112.220 217.295 ;
        RECT 113.815 216.895 116.250 217.295 ;
        RECT 117.845 216.895 120.280 217.295 ;
        RECT 121.875 216.895 124.310 217.295 ;
        RECT 125.905 216.895 128.340 217.295 ;
        RECT 129.935 216.895 132.370 217.295 ;
        RECT 133.965 216.895 136.400 217.295 ;
        RECT 137.995 216.895 140.430 217.295 ;
        RECT 142.025 216.895 144.460 217.295 ;
        RECT 146.055 216.895 148.490 217.295 ;
        RECT 150.085 216.895 152.520 217.295 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 111.820 205.955 112.220 206.755 ;
        RECT 115.850 205.955 116.250 206.755 ;
        RECT 119.880 205.955 120.280 206.755 ;
        RECT 123.910 205.955 124.310 206.755 ;
        RECT 127.940 205.955 128.340 206.755 ;
        RECT 131.970 205.955 132.370 206.755 ;
        RECT 136.000 205.955 136.400 206.755 ;
        RECT 140.030 205.955 140.430 206.755 ;
        RECT 144.060 205.955 144.460 206.755 ;
        RECT 148.090 205.955 148.490 206.755 ;
        RECT 152.120 205.955 152.520 206.755 ;
        RECT 109.240 204.745 111.675 205.545 ;
        RECT 113.270 204.745 115.705 205.545 ;
        RECT 117.300 204.745 119.735 205.545 ;
        RECT 121.330 204.745 123.765 205.545 ;
        RECT 125.360 204.745 127.795 205.545 ;
        RECT 129.390 204.745 131.825 205.545 ;
        RECT 133.420 204.745 135.855 205.545 ;
        RECT 137.450 204.745 139.885 205.545 ;
        RECT 141.480 204.745 143.915 205.545 ;
        RECT 145.510 204.745 147.945 205.545 ;
        RECT 149.540 204.745 151.975 205.545 ;
        RECT 108.540 202.425 108.940 202.625 ;
        RECT 109.785 202.425 110.385 204.345 ;
        RECT 108.540 202.025 110.385 202.425 ;
        RECT 108.540 201.825 108.940 202.025 ;
        RECT 109.785 199.970 110.385 202.025 ;
        RECT 111.075 199.970 111.675 204.745 ;
        RECT 112.570 202.425 112.970 202.625 ;
        RECT 113.815 202.425 114.415 204.345 ;
        RECT 112.570 202.025 114.415 202.425 ;
        RECT 112.570 201.825 112.970 202.025 ;
        RECT 113.815 199.970 114.415 202.025 ;
        RECT 115.105 199.970 115.705 204.745 ;
        RECT 116.600 202.425 117.000 202.625 ;
        RECT 117.845 202.425 118.445 204.345 ;
        RECT 116.600 202.025 118.445 202.425 ;
        RECT 116.600 201.825 117.000 202.025 ;
        RECT 117.845 199.970 118.445 202.025 ;
        RECT 119.135 199.970 119.735 204.745 ;
        RECT 120.630 202.425 121.030 202.625 ;
        RECT 121.875 202.425 122.475 204.345 ;
        RECT 120.630 202.025 122.475 202.425 ;
        RECT 120.630 201.825 121.030 202.025 ;
        RECT 121.875 199.970 122.475 202.025 ;
        RECT 123.165 199.970 123.765 204.745 ;
        RECT 124.660 202.425 125.060 202.625 ;
        RECT 125.905 202.425 126.505 204.345 ;
        RECT 124.660 202.025 126.505 202.425 ;
        RECT 124.660 201.825 125.060 202.025 ;
        RECT 125.905 199.970 126.505 202.025 ;
        RECT 127.195 199.970 127.795 204.745 ;
        RECT 128.690 202.425 129.090 202.625 ;
        RECT 129.935 202.425 130.535 204.345 ;
        RECT 128.690 202.025 130.535 202.425 ;
        RECT 128.690 201.825 129.090 202.025 ;
        RECT 129.935 199.970 130.535 202.025 ;
        RECT 131.225 199.970 131.825 204.745 ;
        RECT 132.720 202.425 133.120 202.625 ;
        RECT 133.965 202.425 134.565 204.345 ;
        RECT 132.720 202.025 134.565 202.425 ;
        RECT 132.720 201.825 133.120 202.025 ;
        RECT 133.965 199.970 134.565 202.025 ;
        RECT 135.255 199.970 135.855 204.745 ;
        RECT 136.750 202.425 137.150 202.625 ;
        RECT 137.995 202.425 138.595 204.345 ;
        RECT 136.750 202.025 138.595 202.425 ;
        RECT 136.750 201.825 137.150 202.025 ;
        RECT 137.995 199.970 138.595 202.025 ;
        RECT 139.285 199.970 139.885 204.745 ;
        RECT 140.780 202.425 141.180 202.625 ;
        RECT 142.025 202.425 142.625 204.345 ;
        RECT 140.780 202.025 142.625 202.425 ;
        RECT 140.780 201.825 141.180 202.025 ;
        RECT 142.025 199.970 142.625 202.025 ;
        RECT 143.315 199.970 143.915 204.745 ;
        RECT 144.810 202.425 145.210 202.625 ;
        RECT 146.055 202.425 146.655 204.345 ;
        RECT 144.810 202.025 146.655 202.425 ;
        RECT 144.810 201.825 145.210 202.025 ;
        RECT 146.055 199.970 146.655 202.025 ;
        RECT 147.345 199.970 147.945 204.745 ;
        RECT 148.840 202.425 149.240 202.625 ;
        RECT 150.085 202.425 150.685 204.345 ;
        RECT 148.840 202.025 150.685 202.425 ;
        RECT 148.840 201.825 149.240 202.025 ;
        RECT 150.085 199.970 150.685 202.025 ;
        RECT 151.375 199.970 151.975 204.745 ;
        RECT 165.405 202.290 165.685 222.410 ;
        RECT 175.065 202.290 175.345 223.010 ;
        RECT 184.725 202.290 185.005 223.610 ;
        RECT 194.385 202.290 194.665 224.210 ;
        RECT 204.045 202.290 204.325 224.810 ;
        RECT 213.705 202.290 213.985 225.410 ;
        RECT 246.615 225.060 247.015 225.660 ;
        RECT 223.365 224.460 223.645 224.510 ;
        RECT 232.965 224.460 233.365 225.060 ;
        RECT 223.305 223.860 223.705 224.460 ;
        RECT 223.365 202.290 223.645 223.860 ;
        RECT 233.025 202.290 233.305 224.460 ;
        RECT 246.665 218.450 246.965 225.060 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 165.475 201.140 165.615 202.290 ;
        RECT 175.135 201.140 175.275 202.290 ;
        RECT 177.645 201.305 179.185 201.675 ;
        RECT 184.795 201.140 184.935 202.290 ;
        RECT 194.455 201.140 194.595 202.290 ;
        RECT 204.115 201.140 204.255 202.290 ;
        RECT 213.775 201.140 213.915 202.290 ;
        RECT 217.645 201.305 219.185 201.675 ;
        RECT 223.435 201.140 223.575 202.290 ;
        RECT 233.095 201.140 233.235 202.290 ;
        RECT 165.415 200.820 165.675 201.140 ;
        RECT 175.075 200.820 175.335 201.140 ;
        RECT 184.735 200.820 184.995 201.140 ;
        RECT 194.395 200.820 194.655 201.140 ;
        RECT 204.055 200.820 204.315 201.140 ;
        RECT 213.715 200.820 213.975 201.140 ;
        RECT 223.375 200.820 223.635 201.140 ;
        RECT 233.035 200.820 233.295 201.140 ;
        RECT 167.255 199.800 167.515 200.120 ;
        RECT 175.535 199.800 175.795 200.120 ;
        RECT 185.195 199.800 185.455 200.120 ;
        RECT 194.855 199.800 195.115 200.120 ;
        RECT 204.515 199.800 204.775 200.120 ;
        RECT 214.175 199.800 214.435 200.120 ;
        RECT 223.835 199.800 224.095 200.120 ;
        RECT 233.035 199.800 233.295 200.120 ;
        RECT 109.240 194.440 109.640 199.685 ;
        RECT 109.240 194.040 110.255 194.440 ;
        RECT 109.240 191.285 109.640 192.885 ;
        RECT 110.530 187.540 110.930 198.905 ;
        RECT 111.820 194.440 112.220 199.685 ;
        RECT 111.205 194.040 112.220 194.440 ;
        RECT 113.270 194.440 113.670 199.685 ;
        RECT 113.270 194.040 114.285 194.440 ;
        RECT 111.820 191.285 112.220 192.885 ;
        RECT 113.270 191.285 113.670 192.885 ;
        RECT 114.560 187.540 114.960 198.905 ;
        RECT 115.850 194.440 116.250 199.685 ;
        RECT 115.235 194.040 116.250 194.440 ;
        RECT 117.300 194.440 117.700 199.685 ;
        RECT 117.300 194.040 118.315 194.440 ;
        RECT 115.850 191.285 116.250 192.885 ;
        RECT 117.300 191.285 117.700 192.885 ;
        RECT 118.590 187.540 118.990 198.905 ;
        RECT 119.880 194.440 120.280 199.685 ;
        RECT 119.265 194.040 120.280 194.440 ;
        RECT 121.330 194.440 121.730 199.685 ;
        RECT 121.330 194.040 122.345 194.440 ;
        RECT 119.880 191.285 120.280 192.885 ;
        RECT 121.330 191.285 121.730 192.885 ;
        RECT 122.620 187.540 123.020 198.905 ;
        RECT 123.910 194.440 124.310 199.685 ;
        RECT 123.295 194.040 124.310 194.440 ;
        RECT 125.360 194.440 125.760 199.685 ;
        RECT 125.360 194.040 126.375 194.440 ;
        RECT 123.910 191.285 124.310 192.885 ;
        RECT 125.360 191.285 125.760 192.885 ;
        RECT 126.650 187.540 127.050 198.905 ;
        RECT 127.940 194.440 128.340 199.685 ;
        RECT 127.325 194.040 128.340 194.440 ;
        RECT 129.390 194.440 129.790 199.685 ;
        RECT 129.390 194.040 130.405 194.440 ;
        RECT 127.940 191.285 128.340 192.885 ;
        RECT 129.390 191.285 129.790 192.885 ;
        RECT 130.680 187.540 131.080 198.905 ;
        RECT 131.970 194.440 132.370 199.685 ;
        RECT 131.355 194.040 132.370 194.440 ;
        RECT 133.420 194.440 133.820 199.685 ;
        RECT 133.420 194.040 134.435 194.440 ;
        RECT 131.970 191.285 132.370 192.885 ;
        RECT 133.420 191.285 133.820 192.885 ;
        RECT 134.710 187.540 135.110 198.905 ;
        RECT 136.000 194.440 136.400 199.685 ;
        RECT 135.385 194.040 136.400 194.440 ;
        RECT 137.450 194.440 137.850 199.685 ;
        RECT 137.450 194.040 138.465 194.440 ;
        RECT 136.000 191.285 136.400 192.885 ;
        RECT 137.450 191.285 137.850 192.885 ;
        RECT 138.740 187.540 139.140 198.905 ;
        RECT 140.030 194.440 140.430 199.685 ;
        RECT 139.415 194.040 140.430 194.440 ;
        RECT 141.480 194.440 141.880 199.685 ;
        RECT 141.480 194.040 142.495 194.440 ;
        RECT 140.030 191.285 140.430 192.885 ;
        RECT 141.480 191.285 141.880 192.885 ;
        RECT 142.770 187.540 143.170 198.905 ;
        RECT 144.060 194.440 144.460 199.685 ;
        RECT 143.445 194.040 144.460 194.440 ;
        RECT 145.510 194.440 145.910 199.685 ;
        RECT 145.510 194.040 146.525 194.440 ;
        RECT 144.060 191.285 144.460 192.885 ;
        RECT 145.510 191.285 145.910 192.885 ;
        RECT 146.800 187.540 147.200 198.905 ;
        RECT 148.090 194.440 148.490 199.685 ;
        RECT 147.475 194.040 148.490 194.440 ;
        RECT 149.540 194.440 149.940 199.685 ;
        RECT 149.540 194.040 150.555 194.440 ;
        RECT 148.090 191.285 148.490 192.885 ;
        RECT 149.540 191.285 149.940 192.885 ;
        RECT 150.830 187.540 151.230 198.905 ;
        RECT 152.120 194.440 152.520 199.685 ;
        RECT 164.035 199.460 164.295 199.780 ;
        RECT 164.095 197.935 164.235 199.460 ;
        RECT 164.025 197.565 164.305 197.935 ;
        RECT 151.505 194.040 152.520 194.440 ;
        RECT 152.120 191.285 152.520 192.885 ;
        RECT 166.335 190.960 166.595 191.280 ;
        RECT 163.575 188.920 163.835 189.240 ;
        RECT 164.035 188.920 164.295 189.240 ;
        RECT 163.635 188.415 163.775 188.920 ;
        RECT 163.565 188.045 163.845 188.415 ;
        RECT 109.240 184.370 109.640 184.770 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 163.115 186.540 163.375 186.860 ;
        RECT 109.240 183.970 154.345 184.370 ;
        RECT 153.945 183.570 154.345 183.970 ;
        RECT 115.265 175.815 117.965 176.215 ;
        RECT 119.885 175.815 122.585 176.215 ;
        RECT 124.505 175.815 127.205 176.215 ;
        RECT 129.125 175.815 131.825 176.215 ;
        RECT 133.745 175.815 136.445 176.215 ;
        RECT 138.365 175.815 141.065 176.215 ;
        RECT 142.985 175.815 145.685 176.215 ;
        RECT 147.605 175.815 150.305 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 163.175 176.660 163.315 186.540 ;
        RECT 163.565 178.525 163.845 178.895 ;
        RECT 163.635 178.360 163.775 178.525 ;
        RECT 163.575 178.040 163.835 178.360 ;
        RECT 164.095 177.535 164.235 188.920 ;
        RECT 165.415 186.540 165.675 186.860 ;
        RECT 164.495 183.480 164.755 183.800 ;
        RECT 164.555 180.400 164.695 183.480 ;
        RECT 164.955 182.800 165.215 183.120 ;
        RECT 165.015 181.615 165.155 182.800 ;
        RECT 164.945 181.245 165.225 181.615 ;
        RECT 164.495 180.080 164.755 180.400 ;
        RECT 165.475 178.215 165.615 186.540 ;
        RECT 166.395 181.760 166.535 190.960 ;
        RECT 167.315 187.540 167.455 199.800 ;
        RECT 175.075 199.460 175.335 199.780 ;
        RECT 175.135 195.020 175.275 199.460 ;
        RECT 175.075 194.700 175.335 195.020 ;
        RECT 173.235 193.680 173.495 194.000 ;
        RECT 168.175 191.980 168.435 192.300 ;
        RECT 167.255 187.220 167.515 187.540 ;
        RECT 166.795 186.540 167.055 186.860 ;
        RECT 166.855 184.820 166.995 186.540 ;
        RECT 168.235 186.260 168.375 191.980 ;
        RECT 171.395 191.300 171.655 191.620 ;
        RECT 170.015 189.150 170.275 189.240 ;
        RECT 170.015 189.010 170.675 189.150 ;
        RECT 170.015 188.920 170.275 189.010 ;
        RECT 169.095 188.240 169.355 188.560 ;
        RECT 168.235 186.120 168.835 186.260 ;
        RECT 168.175 185.520 168.435 185.840 ;
        RECT 166.795 184.500 167.055 184.820 ;
        RECT 167.255 184.160 167.515 184.480 ;
        RECT 166.795 183.480 167.055 183.800 ;
        RECT 166.335 181.440 166.595 181.760 ;
        RECT 166.855 180.740 166.995 183.480 ;
        RECT 166.795 180.420 167.055 180.740 ;
        RECT 167.315 179.380 167.455 184.160 ;
        RECT 168.235 184.140 168.375 185.520 ;
        RECT 168.175 183.820 168.435 184.140 ;
        RECT 167.715 183.480 167.975 183.800 ;
        RECT 167.775 182.100 167.915 183.480 ;
        RECT 168.175 183.140 168.435 183.460 ;
        RECT 167.715 181.780 167.975 182.100 ;
        RECT 167.715 180.080 167.975 180.400 ;
        RECT 167.255 179.060 167.515 179.380 ;
        RECT 165.405 177.845 165.685 178.215 ;
        RECT 165.875 178.040 166.135 178.360 ;
        RECT 164.025 177.165 164.305 177.535 ;
        RECT 163.115 176.340 163.375 176.660 ;
        RECT 165.935 175.640 166.075 178.040 ;
        RECT 165.875 175.320 166.135 175.640 ;
        RECT 167.775 175.300 167.915 180.080 ;
        RECT 168.235 179.380 168.375 183.140 ;
        RECT 168.695 181.500 168.835 186.120 ;
        RECT 169.155 182.295 169.295 188.240 ;
        RECT 170.005 188.045 170.285 188.415 ;
        RECT 169.545 187.365 169.825 187.735 ;
        RECT 169.615 187.200 169.755 187.365 ;
        RECT 169.555 186.880 169.815 187.200 ;
        RECT 169.555 186.200 169.815 186.520 ;
        RECT 169.615 184.820 169.755 186.200 ;
        RECT 169.555 184.500 169.815 184.820 ;
        RECT 170.075 184.480 170.215 188.045 ;
        RECT 170.015 184.160 170.275 184.480 ;
        RECT 170.075 183.800 170.215 184.160 ;
        RECT 169.555 183.480 169.815 183.800 ;
        RECT 170.015 183.480 170.275 183.800 ;
        RECT 169.085 181.925 169.365 182.295 ;
        RECT 169.615 181.760 169.755 183.480 ;
        RECT 170.005 181.925 170.285 182.295 ;
        RECT 168.695 181.360 169.295 181.500 ;
        RECT 169.555 181.440 169.815 181.760 ;
        RECT 170.075 181.420 170.215 181.925 ;
        RECT 168.635 180.760 168.895 181.080 ;
        RECT 169.155 180.820 169.295 181.360 ;
        RECT 170.015 181.100 170.275 181.420 ;
        RECT 168.175 179.060 168.435 179.380 ;
        RECT 168.695 178.895 168.835 180.760 ;
        RECT 169.155 180.680 170.215 180.820 ;
        RECT 169.095 180.080 169.355 180.400 ;
        RECT 168.625 178.525 168.905 178.895 ;
        RECT 168.695 178.360 168.835 178.525 ;
        RECT 169.155 178.360 169.295 180.080 ;
        RECT 168.635 178.040 168.895 178.360 ;
        RECT 169.095 178.040 169.355 178.360 ;
        RECT 169.555 178.040 169.815 178.360 ;
        RECT 169.615 176.855 169.755 178.040 ;
        RECT 169.545 176.485 169.825 176.855 ;
        RECT 170.075 176.290 170.215 180.680 ;
        RECT 170.535 178.950 170.675 189.010 ;
        RECT 170.935 188.580 171.195 188.900 ;
        RECT 170.995 187.735 171.135 188.580 ;
        RECT 171.455 188.560 171.595 191.300 ;
        RECT 171.855 190.960 172.115 191.280 ;
        RECT 171.915 189.240 172.055 190.960 ;
        RECT 171.855 188.920 172.115 189.240 ;
        RECT 172.775 188.920 173.035 189.240 ;
        RECT 171.395 188.240 171.655 188.560 ;
        RECT 170.925 187.365 171.205 187.735 ;
        RECT 170.935 187.110 171.195 187.200 ;
        RECT 171.915 187.110 172.055 188.920 ;
        RECT 170.935 186.970 172.055 187.110 ;
        RECT 170.935 186.880 171.195 186.970 ;
        RECT 171.455 184.335 171.595 186.970 ;
        RECT 172.835 186.860 172.975 188.920 ;
        RECT 173.295 187.540 173.435 193.680 ;
        RECT 175.135 192.300 175.275 194.700 ;
        RECT 175.075 191.980 175.335 192.300 ;
        RECT 174.615 189.095 174.875 189.240 ;
        RECT 174.605 188.725 174.885 189.095 ;
        RECT 175.595 187.540 175.735 199.800 ;
        RECT 180.945 198.585 182.485 198.955 ;
        RECT 177.645 195.865 179.185 196.235 ;
        RECT 176.915 194.360 177.175 194.680 ;
        RECT 175.995 191.980 176.255 192.300 ;
        RECT 176.055 190.260 176.195 191.980 ;
        RECT 176.455 191.640 176.715 191.960 ;
        RECT 175.995 189.940 176.255 190.260 ;
        RECT 175.995 188.920 176.255 189.240 ;
        RECT 173.235 187.220 173.495 187.540 ;
        RECT 175.535 187.220 175.795 187.540 ;
        RECT 172.775 186.770 173.035 186.860 ;
        RECT 172.375 186.630 173.035 186.770 ;
        RECT 171.855 185.520 172.115 185.840 ;
        RECT 171.385 183.965 171.665 184.335 ;
        RECT 170.935 183.140 171.195 183.460 ;
        RECT 170.995 182.295 171.135 183.140 ;
        RECT 170.925 181.925 171.205 182.295 ;
        RECT 171.455 181.080 171.595 183.965 ;
        RECT 171.395 180.760 171.655 181.080 ;
        RECT 171.915 180.935 172.055 185.520 ;
        RECT 172.375 183.460 172.515 186.630 ;
        RECT 172.775 186.540 173.035 186.630 ;
        RECT 174.615 186.540 174.875 186.860 ;
        RECT 174.155 186.200 174.415 186.520 ;
        RECT 172.775 183.480 173.035 183.800 ;
        RECT 173.235 183.480 173.495 183.800 ;
        RECT 173.695 183.480 173.955 183.800 ;
        RECT 172.315 183.140 172.575 183.460 ;
        RECT 172.375 181.760 172.515 183.140 ;
        RECT 172.835 182.975 172.975 183.480 ;
        RECT 172.765 182.605 173.045 182.975 ;
        RECT 172.315 181.440 172.575 181.760 ;
        RECT 172.765 181.245 173.045 181.615 ;
        RECT 172.775 181.100 173.035 181.245 ;
        RECT 171.845 180.565 172.125 180.935 ;
        RECT 173.295 179.290 173.435 183.480 ;
        RECT 173.755 182.100 173.895 183.480 ;
        RECT 173.695 181.780 173.955 182.100 ;
        RECT 173.695 179.290 173.955 179.380 ;
        RECT 173.295 179.150 173.955 179.290 ;
        RECT 173.695 179.060 173.955 179.150 ;
        RECT 170.535 178.810 172.055 178.950 ;
        RECT 171.395 178.040 171.655 178.360 ;
        RECT 171.915 178.270 172.055 178.810 ;
        RECT 172.775 178.780 173.035 179.040 ;
        RECT 174.215 178.780 174.355 186.200 ;
        RECT 174.675 184.820 174.815 186.540 ;
        RECT 176.055 185.840 176.195 188.920 ;
        RECT 175.995 185.520 176.255 185.840 ;
        RECT 174.615 184.500 174.875 184.820 ;
        RECT 175.075 184.160 175.335 184.480 ;
        RECT 175.525 184.220 175.805 184.335 ;
        RECT 176.055 184.220 176.195 185.520 ;
        RECT 175.135 179.460 175.275 184.160 ;
        RECT 175.525 184.080 176.195 184.220 ;
        RECT 175.525 183.965 175.805 184.080 ;
        RECT 175.595 183.800 175.735 183.965 ;
        RECT 175.535 183.480 175.795 183.800 ;
        RECT 176.515 183.540 176.655 191.640 ;
        RECT 176.975 188.415 177.115 194.360 ;
        RECT 178.755 194.020 179.015 194.340 ;
        RECT 178.815 192.980 178.955 194.020 ;
        RECT 180.945 193.145 182.485 193.515 ;
        RECT 185.255 192.980 185.395 199.800 ;
        RECT 187.035 193.680 187.295 194.000 ;
        RECT 178.755 192.660 179.015 192.980 ;
        RECT 185.195 192.660 185.455 192.980 ;
        RECT 187.095 192.300 187.235 193.680 ;
        RECT 194.915 192.980 195.055 199.800 ;
        RECT 199.455 194.700 199.715 195.020 ;
        RECT 194.855 192.660 195.115 192.980 ;
        RECT 189.795 192.320 190.055 192.640 ;
        RECT 182.895 191.980 183.155 192.300 ;
        RECT 187.035 191.980 187.295 192.300 ;
        RECT 189.335 191.980 189.595 192.300 ;
        RECT 179.675 190.960 179.935 191.280 ;
        RECT 177.645 190.425 179.185 190.795 ;
        RECT 177.365 189.405 177.645 189.775 ;
        RECT 177.435 188.560 177.575 189.405 ;
        RECT 179.215 188.920 179.475 189.240 ;
        RECT 176.905 188.045 177.185 188.415 ;
        RECT 177.375 188.240 177.635 188.560 ;
        RECT 179.275 188.415 179.415 188.920 ;
        RECT 176.915 186.540 177.175 186.860 ;
        RECT 176.975 186.375 177.115 186.540 ;
        RECT 176.905 186.005 177.185 186.375 ;
        RECT 177.435 185.750 177.575 188.240 ;
        RECT 179.205 188.045 179.485 188.415 ;
        RECT 177.835 186.540 178.095 186.860 ;
        RECT 177.895 186.180 178.035 186.540 ;
        RECT 177.835 185.860 178.095 186.180 ;
        RECT 176.055 183.400 176.655 183.540 ;
        RECT 176.975 185.610 177.575 185.750 ;
        RECT 175.525 181.925 175.805 182.295 ;
        RECT 175.535 181.780 175.795 181.925 ;
        RECT 175.535 180.420 175.795 180.740 ;
        RECT 172.775 178.720 174.355 178.780 ;
        RECT 172.835 178.640 174.355 178.720 ;
        RECT 174.675 179.320 175.275 179.460 ;
        RECT 171.915 178.130 172.975 178.270 ;
        RECT 170.925 177.165 171.205 177.535 ;
        RECT 170.995 176.290 171.135 177.165 ;
        RECT 171.455 176.320 171.595 178.040 ;
        RECT 172.315 177.535 172.575 177.680 ;
        RECT 172.305 177.165 172.585 177.535 ;
        RECT 172.315 176.570 172.575 176.660 ;
        RECT 171.915 176.430 172.575 176.570 ;
        RECT 167.715 174.980 167.975 175.300 ;
        RECT 114.835 172.120 118.395 174.820 ;
        RECT 119.155 172.120 123.015 174.820 ;
        RECT 123.775 172.120 127.635 174.820 ;
        RECT 128.395 172.120 132.255 174.820 ;
        RECT 133.015 172.120 136.875 174.820 ;
        RECT 137.635 172.120 141.495 174.820 ;
        RECT 142.255 172.120 146.115 174.820 ;
        RECT 146.875 172.120 150.735 174.820 ;
        RECT 57.020 169.775 57.820 169.890 ;
        RECT 9.500 168.275 58.420 169.775 ;
        RECT 9.500 165.715 56.920 166.715 ;
        RECT 103.350 164.990 103.750 170.890 ;
        RECT 105.930 168.490 106.330 170.890 ;
        RECT 9.500 163.915 55.070 164.915 ;
        RECT 102.625 164.590 103.750 164.990 ;
        RECT 104.640 164.790 105.040 167.190 ;
        RECT 107.380 164.990 107.780 170.890 ;
        RECT 109.960 168.490 110.360 170.890 ;
        RECT 115.625 169.795 117.605 170.845 ;
        RECT 119.155 169.795 119.755 172.120 ;
        RECT 115.625 169.195 119.755 169.795 ;
        RECT 120.245 169.795 122.225 170.845 ;
        RECT 123.775 169.795 124.375 172.120 ;
        RECT 120.245 169.195 124.375 169.795 ;
        RECT 124.865 169.795 126.845 170.845 ;
        RECT 128.395 169.795 128.995 172.120 ;
        RECT 124.865 169.195 128.995 169.795 ;
        RECT 129.485 169.795 131.465 170.845 ;
        RECT 133.015 169.795 133.615 172.120 ;
        RECT 129.485 169.195 133.615 169.795 ;
        RECT 134.105 169.795 136.085 170.845 ;
        RECT 137.635 169.795 138.235 172.120 ;
        RECT 134.105 169.195 138.235 169.795 ;
        RECT 138.725 169.795 140.705 170.845 ;
        RECT 142.255 169.795 142.855 172.120 ;
        RECT 138.725 169.195 142.855 169.795 ;
        RECT 143.345 169.795 145.325 170.845 ;
        RECT 146.875 169.795 147.475 172.120 ;
        RECT 143.345 169.195 147.475 169.795 ;
        RECT 115.625 168.145 117.605 169.195 ;
        RECT 120.245 168.145 122.225 169.195 ;
        RECT 124.865 168.145 126.845 169.195 ;
        RECT 129.485 168.145 131.465 169.195 ;
        RECT 134.105 168.145 136.085 169.195 ;
        RECT 138.725 168.145 140.705 169.195 ;
        RECT 143.345 168.145 145.325 169.195 ;
        RECT 147.965 168.145 150.345 170.845 ;
        RECT 106.655 164.590 107.780 164.990 ;
        RECT 108.670 164.790 109.070 167.190 ;
        RECT 9.500 162.115 51.610 163.115 ;
        RECT 9.500 159.815 53.170 161.315 ;
        RECT 2.705 157.015 51.610 159.015 ;
        RECT 2.705 1.285 3.505 157.015 ;
        RECT 9.500 154.715 53.170 156.215 ;
        RECT 9.500 152.915 51.610 153.915 ;
        RECT 9.500 151.115 55.070 152.115 ;
        RECT 74.940 151.875 86.100 155.595 ;
        RECT 9.500 149.315 56.520 150.315 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 148.155 78.660 151.875 ;
        RECT 80.100 149.595 80.930 150.425 ;
        RECT 82.380 148.155 86.100 151.875 ;
        RECT 102.625 149.850 103.025 164.590 ;
        RECT 103.350 162.940 104.365 163.340 ;
        RECT 105.315 162.940 106.330 163.340 ;
        RECT 103.350 159.695 103.750 162.940 ;
        RECT 105.930 160.395 106.330 162.940 ;
        RECT 104.190 159.795 106.330 160.395 ;
        RECT 104.190 159.410 104.495 159.795 ;
        RECT 105.930 159.695 106.330 159.795 ;
        RECT 103.895 154.535 104.495 159.410 ;
        RECT 105.185 155.035 105.785 159.410 ;
        RECT 103.895 153.935 106.330 154.535 ;
        RECT 103.350 150.640 103.750 153.565 ;
        RECT 105.930 152.190 106.330 153.935 ;
        RECT 103.895 151.790 106.330 152.190 ;
        RECT 103.895 151.015 104.495 151.790 ;
        RECT 105.185 150.640 105.785 151.415 ;
        RECT 103.350 150.240 105.785 150.640 ;
        RECT 106.655 149.850 107.055 164.590 ;
        RECT 107.380 162.940 108.395 163.340 ;
        RECT 109.345 162.940 110.360 163.340 ;
        RECT 107.380 159.695 107.780 162.940 ;
        RECT 109.960 160.395 110.360 162.940 ;
        RECT 108.220 159.795 110.360 160.395 ;
        RECT 108.220 159.410 108.525 159.795 ;
        RECT 109.960 159.695 110.360 159.795 ;
        RECT 107.925 154.535 108.525 159.410 ;
        RECT 109.215 155.035 109.815 159.410 ;
        RECT 107.925 153.935 110.360 154.535 ;
        RECT 107.380 150.640 107.780 153.565 ;
        RECT 109.960 152.190 110.360 153.935 ;
        RECT 107.925 151.790 110.360 152.190 ;
        RECT 107.925 151.015 108.525 151.790 ;
        RECT 109.215 150.640 109.815 151.415 ;
        RECT 107.380 150.240 109.815 150.640 ;
        RECT 102.625 149.450 103.750 149.850 ;
        RECT 74.940 144.435 86.100 148.155 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 11.195 139.800 23.015 140.200 ;
        RECT 11.195 137.185 11.795 139.800 ;
        RECT 14.860 138.370 21.050 138.770 ;
        RECT 14.860 137.585 15.260 138.370 ;
        RECT 20.650 137.970 21.050 138.370 ;
        RECT 14.130 137.185 16.020 137.585 ;
        RECT 16.805 137.185 18.955 137.585 ;
        RECT 16.805 136.875 17.205 137.185 ;
        RECT 11.940 136.275 15.275 136.875 ;
        RECT 16.165 136.275 17.205 136.875 ;
        RECT 5.910 132.225 7.510 135.425 ;
        RECT 13.485 133.130 14.085 135.875 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 16.805 129.110 17.205 136.275 ;
        RECT 19.100 136.125 20.750 136.725 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 19.100 128.925 19.500 136.125 ;
        RECT 22.615 134.120 23.015 139.800 ;
        RECT 24.255 135.155 25.755 143.745 ;
        RECT 27.765 135.155 29.265 143.745 ;
        RECT 36.055 135.155 37.555 143.745 ;
        RECT 44.345 135.155 45.845 143.745 ;
        RECT 52.635 135.155 54.135 143.745 ;
        RECT 56.145 135.155 57.645 143.745 ;
        RECT 103.350 143.435 103.750 149.450 ;
        RECT 104.640 147.135 105.040 149.535 ;
        RECT 106.655 149.450 107.780 149.850 ;
        RECT 105.930 143.435 106.330 145.835 ;
        RECT 107.380 143.435 107.780 149.450 ;
        RECT 108.670 147.135 109.070 149.535 ;
        RECT 109.960 143.435 110.360 145.835 ;
        RECT 116.310 143.410 116.910 168.145 ;
        RECT 120.930 147.550 121.530 168.145 ;
        RECT 125.550 159.440 126.150 168.145 ;
        RECT 125.550 158.840 128.940 159.440 ;
        RECT 120.930 146.950 126.935 147.550 ;
        RECT 122.645 144.030 124.245 144.830 ;
        RECT 128.340 144.540 128.940 158.840 ;
        RECT 130.170 148.610 130.770 168.145 ;
        RECT 134.795 164.330 135.395 168.145 ;
        RECT 133.685 163.140 134.485 163.740 ;
        RECT 133.785 155.610 134.385 163.140 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 139.410 157.075 140.010 168.145 ;
        RECT 144.035 163.040 144.635 168.145 ;
        RECT 146.855 164.430 147.655 165.030 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 141.615 158.550 142.415 159.150 ;
        RECT 138.070 156.475 140.010 157.075 ;
        RECT 133.285 155.010 134.885 155.610 ;
        RECT 133.275 151.400 134.875 152.200 ;
        RECT 133.275 150.230 134.875 151.030 ;
        RECT 138.070 149.760 138.670 156.475 ;
        RECT 141.715 152.110 142.315 158.550 ;
        RECT 141.215 151.905 142.815 152.110 ;
        RECT 140.950 151.505 143.050 151.905 ;
        RECT 133.285 149.160 138.670 149.760 ;
        RECT 130.170 148.010 134.430 148.610 ;
        RECT 130.615 146.830 132.215 147.630 ;
        RECT 133.285 147.410 134.885 148.010 ;
        RECT 138.525 147.310 140.125 148.110 ;
        RECT 128.340 143.940 134.885 144.540 ;
        RECT 138.525 143.820 140.125 144.620 ;
        RECT 116.310 142.810 132.215 143.410 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 141.990 142.815 142.790 ;
        RECT 146.955 142.730 147.555 164.430 ;
        RECT 148.655 158.450 149.255 168.145 ;
        RECT 146.455 142.640 148.055 142.730 ;
        RECT 146.195 142.240 148.295 142.640 ;
        RECT 146.455 142.130 148.055 142.240 ;
        RECT 104.640 139.365 152.360 140.165 ;
        RECT 97.200 137.420 147.750 138.220 ;
        RECT 107.380 135.525 132.465 136.325 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 56.145 133.555 77.110 135.155 ;
        RECT 80.120 133.320 137.265 134.120 ;
        RECT 137.945 133.410 144.375 133.810 ;
        RECT 21.615 131.745 135.665 132.545 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 142.980 131.990 143.630 132.590 ;
        RECT 27.065 129.995 134.065 130.795 ;
        RECT 19.100 128.125 101.315 128.925 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 142.980 126.815 143.230 131.990 ;
        RECT 144.025 131.050 144.375 133.410 ;
        RECT 143.725 129.545 144.425 131.050 ;
        RECT 153.945 129.545 154.345 129.945 ;
        RECT 143.725 129.145 154.345 129.545 ;
        RECT 143.725 127.640 144.425 129.145 ;
        RECT 142.980 126.215 143.630 126.815 ;
        RECT 10.025 122.800 70.175 123.810 ;
        RECT 71.775 122.750 114.165 123.850 ;
        RECT 10.025 120.300 70.175 122.300 ;
        RECT 71.775 121.250 114.165 122.350 ;
        RECT 115.905 121.575 128.935 123.145 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 10.025 117.800 70.175 119.800 ;
        RECT 71.775 119.750 114.165 120.850 ;
        RECT 71.775 118.250 114.165 119.350 ;
        RECT 10.025 115.300 70.175 117.300 ;
        RECT 71.775 116.750 114.165 117.850 ;
        RECT 115.905 117.075 128.935 118.645 ;
        RECT 141.900 116.370 150.745 117.170 ;
        RECT 71.775 115.250 114.165 116.350 ;
        RECT 10.025 112.780 70.175 114.800 ;
        RECT 71.775 112.730 114.165 114.850 ;
        RECT 136.465 114.770 144.870 115.570 ;
        RECT 170.005 115.285 170.285 176.290 ;
        RECT 115.905 112.615 128.935 114.185 ;
        RECT 10.025 110.280 70.175 112.280 ;
        RECT 71.775 111.230 114.165 112.330 ;
        RECT 133.265 111.795 141.675 112.595 ;
        RECT 10.025 107.780 70.175 109.780 ;
        RECT 71.775 109.730 114.165 110.830 ;
        RECT 140.875 110.315 141.675 111.795 ;
        RECT 144.070 110.315 144.870 114.770 ;
        RECT 164.025 115.005 170.285 115.285 ;
        RECT 71.775 108.230 114.165 109.330 ;
        RECT 115.905 108.115 128.935 109.685 ;
        RECT 139.560 109.515 142.995 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 10.025 105.280 70.175 107.280 ;
        RECT 71.775 106.730 114.165 107.830 ;
        RECT 71.775 105.230 114.165 106.330 ;
        RECT 10.025 103.770 70.175 104.780 ;
        RECT 71.775 103.730 114.165 104.830 ;
        RECT 115.905 103.655 128.935 105.225 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 10.025 91.525 128.935 92.775 ;
        RECT 10.025 89.640 128.935 91.140 ;
        RECT 10.025 85.640 128.935 88.640 ;
        RECT 136.295 86.115 138.400 90.215 ;
        RECT 10.025 83.140 128.935 84.640 ;
        RECT 10.025 81.505 128.935 82.755 ;
        RECT 10.025 79.620 128.935 81.120 ;
        RECT 136.295 80.265 138.400 85.535 ;
        RECT 139.560 82.025 140.860 109.515 ;
        RECT 141.695 91.385 142.995 109.515 ;
        RECT 141.290 90.795 143.395 91.385 ;
        RECT 139.155 81.435 141.260 82.025 ;
        RECT 10.025 75.620 128.935 78.620 ;
        RECT 136.295 75.585 138.400 79.685 ;
        RECT 10.025 73.120 128.935 74.620 ;
        RECT 10.025 71.485 128.935 72.735 ;
        RECT 10.025 69.600 128.935 71.100 ;
        RECT 136.295 70.905 138.400 75.005 ;
        RECT 10.025 65.600 128.935 68.600 ;
        RECT 136.295 66.225 138.400 70.325 ;
        RECT 10.025 63.100 128.935 64.600 ;
        RECT 10.025 61.465 128.935 62.715 ;
        RECT 10.025 59.580 128.935 61.080 ;
        RECT 136.295 60.375 138.400 65.645 ;
        RECT 10.025 55.580 128.935 58.580 ;
        RECT 136.295 55.695 138.400 59.795 ;
        RECT 10.025 53.080 128.935 54.580 ;
        RECT 10.025 51.445 128.935 52.695 ;
        RECT 136.295 51.015 138.400 55.115 ;
        RECT 12.915 45.565 14.515 47.165 ;
        RECT 90.715 45.565 92.315 47.165 ;
        RECT 136.295 46.335 138.400 50.435 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 136.295 40.485 138.400 45.755 ;
        RECT 143.835 42.245 145.135 110.315 ;
        RECT 164.025 109.225 164.305 115.005 ;
        RECT 170.925 114.705 171.205 176.290 ;
        RECT 171.395 176.000 171.655 176.320 ;
        RECT 171.915 176.290 172.055 176.430 ;
        RECT 172.315 176.340 172.575 176.430 ;
        RECT 172.835 176.290 172.975 178.130 ;
        RECT 173.235 178.040 173.495 178.360 ;
        RECT 166.325 114.425 171.205 114.705 ;
        RECT 166.325 109.225 166.605 114.425 ;
        RECT 171.845 114.125 172.125 176.290 ;
        RECT 168.625 113.845 172.125 114.125 ;
        RECT 168.625 109.225 168.905 113.845 ;
        RECT 172.765 113.545 173.045 176.290 ;
        RECT 173.295 174.620 173.435 178.040 ;
        RECT 173.685 177.845 173.965 178.215 ;
        RECT 173.755 176.290 173.895 177.845 ;
        RECT 174.155 177.700 174.415 178.020 ;
        RECT 173.235 174.300 173.495 174.620 ;
        RECT 170.925 113.265 173.045 113.545 ;
        RECT 170.925 109.225 171.205 113.265 ;
        RECT 173.685 112.965 173.965 176.290 ;
        RECT 174.215 175.980 174.355 177.700 ;
        RECT 174.675 176.290 174.815 179.320 ;
        RECT 175.595 177.590 175.735 180.420 ;
        RECT 176.055 179.290 176.195 183.400 ;
        RECT 176.455 182.800 176.715 183.120 ;
        RECT 176.515 181.420 176.655 182.800 ;
        RECT 176.975 181.420 177.115 185.610 ;
        RECT 177.645 184.985 179.185 185.355 ;
        RECT 178.295 184.500 178.555 184.820 ;
        RECT 177.365 182.605 177.645 182.975 ;
        RECT 177.835 182.800 178.095 183.120 ;
        RECT 176.455 181.100 176.715 181.420 ;
        RECT 176.915 181.100 177.175 181.420 ;
        RECT 177.435 180.310 177.575 182.605 ;
        RECT 177.895 180.740 178.035 182.800 ;
        RECT 178.355 181.760 178.495 184.500 ;
        RECT 179.735 184.220 179.875 190.960 ;
        RECT 182.955 189.920 183.095 191.980 ;
        RECT 186.575 190.960 186.835 191.280 ;
        RECT 180.655 189.520 181.715 189.660 ;
        RECT 182.895 189.600 183.155 189.920 ;
        RECT 186.635 189.775 186.775 190.960 ;
        RECT 189.395 190.260 189.535 191.980 ;
        RECT 189.855 190.260 189.995 192.320 ;
        RECT 198.535 191.980 198.795 192.300 ;
        RECT 196.235 190.960 196.495 191.280 ;
        RECT 189.335 189.940 189.595 190.260 ;
        RECT 189.795 189.940 190.055 190.260 ;
        RECT 185.185 189.660 185.465 189.775 ;
        RECT 180.655 187.540 180.795 189.520 ;
        RECT 181.575 189.240 181.715 189.520 ;
        RECT 185.185 189.520 186.315 189.660 ;
        RECT 185.185 189.405 185.465 189.520 ;
        RECT 181.055 188.920 181.315 189.240 ;
        RECT 181.515 188.920 181.775 189.240 ;
        RECT 182.895 188.920 183.155 189.240 ;
        RECT 183.355 188.920 183.615 189.240 ;
        RECT 184.735 188.920 184.995 189.240 ;
        RECT 186.175 189.150 186.315 189.520 ;
        RECT 186.565 189.405 186.845 189.775 ;
        RECT 188.415 189.600 188.675 189.920 ;
        RECT 187.035 189.260 187.295 189.580 ;
        RECT 186.575 189.150 186.835 189.240 ;
        RECT 186.175 189.010 186.835 189.150 ;
        RECT 186.575 188.920 186.835 189.010 ;
        RECT 181.115 188.560 181.255 188.920 ;
        RECT 181.055 188.240 181.315 188.560 ;
        RECT 180.945 187.705 182.485 188.075 ;
        RECT 180.595 187.220 180.855 187.540 ;
        RECT 182.955 187.450 183.095 188.920 ;
        RECT 183.415 187.540 183.555 188.920 ;
        RECT 183.815 188.240 184.075 188.560 ;
        RECT 182.035 187.310 183.095 187.450 ;
        RECT 180.135 186.540 180.395 186.860 ;
        RECT 181.045 186.685 181.325 187.055 ;
        RECT 182.035 186.860 182.175 187.310 ;
        RECT 183.355 187.220 183.615 187.540 ;
        RECT 179.275 184.080 179.875 184.220 ;
        RECT 178.295 181.440 178.555 181.760 ;
        RECT 177.835 180.420 178.095 180.740 ;
        RECT 179.275 180.400 179.415 184.080 ;
        RECT 179.675 183.480 179.935 183.800 ;
        RECT 179.735 181.420 179.875 183.480 ;
        RECT 179.675 181.100 179.935 181.420 ;
        RECT 179.675 180.420 179.935 180.740 ;
        RECT 176.975 180.170 177.575 180.310 ;
        RECT 176.055 179.150 176.655 179.290 ;
        RECT 175.985 178.525 176.265 178.895 ;
        RECT 176.055 178.360 176.195 178.525 ;
        RECT 175.995 178.040 176.255 178.360 ;
        RECT 176.515 178.270 176.655 179.150 ;
        RECT 176.975 178.610 177.115 180.170 ;
        RECT 179.215 180.080 179.475 180.400 ;
        RECT 177.645 179.545 179.185 179.915 ;
        RECT 179.735 179.380 179.875 180.420 ;
        RECT 179.675 179.060 179.935 179.380 ;
        RECT 176.975 178.470 178.035 178.610 ;
        RECT 176.515 178.130 177.575 178.270 ;
        RECT 175.595 177.450 176.655 177.590 ;
        RECT 175.135 176.430 175.735 176.570 ;
        RECT 174.155 175.660 174.415 175.980 ;
        RECT 173.225 112.685 173.965 112.965 ;
        RECT 174.605 112.965 174.885 176.290 ;
        RECT 175.135 175.300 175.275 176.430 ;
        RECT 175.595 176.290 175.735 176.430 ;
        RECT 176.515 176.290 176.655 177.450 ;
        RECT 177.435 176.290 177.575 178.130 ;
        RECT 177.895 177.680 178.035 178.470 ;
        RECT 178.755 178.040 179.015 178.360 ;
        RECT 179.675 178.040 179.935 178.360 ;
        RECT 177.835 177.360 178.095 177.680 ;
        RECT 177.895 176.430 178.495 176.570 ;
        RECT 175.075 174.980 175.335 175.300 ;
        RECT 175.525 113.690 175.805 176.290 ;
        RECT 176.445 114.500 176.725 176.290 ;
        RECT 177.365 115.080 177.645 176.290 ;
        RECT 177.895 175.640 178.035 176.430 ;
        RECT 178.355 176.290 178.495 176.430 ;
        RECT 177.835 175.320 178.095 175.640 ;
        RECT 178.285 115.660 178.565 176.290 ;
        RECT 178.815 175.300 178.955 178.040 ;
        RECT 179.205 176.485 179.485 176.855 ;
        RECT 179.275 176.290 179.415 176.485 ;
        RECT 178.755 174.980 179.015 175.300 ;
        RECT 179.205 116.240 179.485 176.290 ;
        RECT 179.735 175.640 179.875 178.040 ;
        RECT 180.195 176.290 180.335 186.540 ;
        RECT 181.115 184.140 181.255 186.685 ;
        RECT 181.975 186.540 182.235 186.860 ;
        RECT 182.895 186.540 183.155 186.860 ;
        RECT 181.515 186.200 181.775 186.520 ;
        RECT 181.575 184.820 181.715 186.200 ;
        RECT 181.515 184.500 181.775 184.820 ;
        RECT 182.435 184.500 182.695 184.820 ;
        RECT 181.055 183.820 181.315 184.140 ;
        RECT 182.495 183.800 182.635 184.500 ;
        RECT 181.505 183.285 181.785 183.655 ;
        RECT 182.435 183.480 182.695 183.800 ;
        RECT 181.515 183.140 181.775 183.285 ;
        RECT 181.055 183.030 181.315 183.120 ;
        RECT 180.655 182.890 181.315 183.030 ;
        RECT 180.655 182.100 180.795 182.890 ;
        RECT 181.055 182.800 181.315 182.890 ;
        RECT 180.945 182.265 182.485 182.635 ;
        RECT 180.595 181.780 180.855 182.100 ;
        RECT 181.975 181.615 182.235 181.760 ;
        RECT 181.965 181.245 182.245 181.615 ;
        RECT 181.055 180.760 181.315 181.080 ;
        RECT 182.435 180.760 182.695 181.080 ;
        RECT 181.115 179.380 181.255 180.760 ;
        RECT 181.975 180.080 182.235 180.400 ;
        RECT 182.035 179.380 182.175 180.080 ;
        RECT 181.055 179.060 181.315 179.380 ;
        RECT 181.975 179.060 182.235 179.380 ;
        RECT 182.495 178.700 182.635 180.760 ;
        RECT 182.435 178.380 182.695 178.700 ;
        RECT 182.955 177.420 183.095 186.540 ;
        RECT 183.355 185.520 183.615 185.840 ;
        RECT 183.415 184.140 183.555 185.520 ;
        RECT 183.355 183.820 183.615 184.140 ;
        RECT 183.355 182.800 183.615 183.120 ;
        RECT 183.415 182.100 183.555 182.800 ;
        RECT 183.355 181.780 183.615 182.100 ;
        RECT 183.355 181.100 183.615 181.420 ;
        RECT 183.415 179.290 183.555 181.100 ;
        RECT 183.875 180.740 184.015 188.240 ;
        RECT 184.795 185.840 184.935 188.920 ;
        RECT 186.105 187.365 186.385 187.735 ;
        RECT 186.635 187.540 186.775 188.920 ;
        RECT 186.175 186.860 186.315 187.365 ;
        RECT 186.575 187.220 186.835 187.540 ;
        RECT 186.115 186.540 186.375 186.860 ;
        RECT 184.735 185.520 184.995 185.840 ;
        RECT 186.575 185.750 186.835 185.840 ;
        RECT 187.095 185.750 187.235 189.260 ;
        RECT 187.495 188.580 187.755 188.900 ;
        RECT 186.575 185.610 187.235 185.750 ;
        RECT 186.575 185.520 186.835 185.610 ;
        RECT 185.655 184.500 185.915 184.820 ;
        RECT 185.195 183.480 185.455 183.800 ;
        RECT 184.275 183.140 184.535 183.460 ;
        RECT 183.815 180.420 184.075 180.740 ;
        RECT 184.335 179.290 184.475 183.140 ;
        RECT 184.735 182.800 184.995 183.120 ;
        RECT 184.795 181.760 184.935 182.800 ;
        RECT 184.735 181.440 184.995 181.760 ;
        RECT 185.255 181.420 185.395 183.480 ;
        RECT 185.195 181.100 185.455 181.420 ;
        RECT 183.415 179.150 184.015 179.290 ;
        RECT 184.335 179.150 184.935 179.290 ;
        RECT 182.955 177.280 183.555 177.420 ;
        RECT 180.945 176.825 182.485 177.195 ;
        RECT 180.595 176.570 180.855 176.660 ;
        RECT 180.595 176.430 181.255 176.570 ;
        RECT 180.595 176.340 180.855 176.430 ;
        RECT 181.115 176.290 181.255 176.430 ;
        RECT 182.035 176.430 182.635 176.570 ;
        RECT 182.885 176.485 183.165 176.855 ;
        RECT 182.035 176.290 182.175 176.430 ;
        RECT 179.675 175.320 179.935 175.640 ;
        RECT 180.125 116.820 180.405 176.290 ;
        RECT 181.045 117.400 181.325 176.290 ;
        RECT 181.965 117.980 182.245 176.290 ;
        RECT 182.495 176.175 182.635 176.430 ;
        RECT 182.955 176.290 183.095 176.485 ;
        RECT 182.425 175.805 182.705 176.175 ;
        RECT 182.885 118.560 183.165 176.290 ;
        RECT 183.415 176.175 183.555 177.280 ;
        RECT 183.875 176.290 184.015 179.150 ;
        RECT 184.265 176.485 184.545 176.855 ;
        RECT 183.345 175.805 183.625 176.175 ;
        RECT 183.805 119.140 184.085 176.290 ;
        RECT 184.335 175.980 184.475 176.485 ;
        RECT 184.795 176.290 184.935 179.150 ;
        RECT 185.195 179.060 185.455 179.380 ;
        RECT 185.255 178.360 185.395 179.060 ;
        RECT 185.195 178.040 185.455 178.360 ;
        RECT 185.715 177.590 185.855 184.500 ;
        RECT 186.635 183.710 186.775 185.520 ;
        RECT 187.035 183.710 187.295 183.800 ;
        RECT 186.635 183.570 187.295 183.710 ;
        RECT 186.115 181.780 186.375 182.100 ;
        RECT 186.175 180.400 186.315 181.780 ;
        RECT 186.635 181.080 186.775 183.570 ;
        RECT 187.035 183.480 187.295 183.570 ;
        RECT 187.035 182.800 187.295 183.120 ;
        RECT 186.575 180.760 186.835 181.080 ;
        RECT 186.115 180.080 186.375 180.400 ;
        RECT 186.635 179.460 186.775 180.760 ;
        RECT 186.175 179.320 186.775 179.460 ;
        RECT 186.175 178.700 186.315 179.320 ;
        RECT 187.095 179.290 187.235 182.800 ;
        RECT 187.555 182.100 187.695 188.580 ;
        RECT 188.475 187.450 188.615 189.600 ;
        RECT 188.875 189.095 189.135 189.240 ;
        RECT 188.865 188.725 189.145 189.095 ;
        RECT 189.855 188.810 189.995 189.940 ;
        RECT 189.395 188.670 189.995 188.810 ;
        RECT 191.235 189.580 191.835 189.660 ;
        RECT 191.235 189.520 191.895 189.580 ;
        RECT 189.395 187.735 189.535 188.670 ;
        RECT 188.475 187.310 189.075 187.450 ;
        RECT 189.325 187.365 189.605 187.735 ;
        RECT 190.715 187.450 190.975 187.540 ;
        RECT 191.235 187.450 191.375 189.520 ;
        RECT 191.635 189.260 191.895 189.520 ;
        RECT 191.635 188.580 191.895 188.900 ;
        RECT 188.415 186.540 188.675 186.860 ;
        RECT 187.955 184.160 188.215 184.480 ;
        RECT 187.495 181.780 187.755 182.100 ;
        RECT 187.095 179.150 187.695 179.290 ;
        RECT 186.575 178.895 186.835 179.040 ;
        RECT 186.115 178.380 186.375 178.700 ;
        RECT 186.565 178.525 186.845 178.895 ;
        RECT 187.035 178.040 187.295 178.360 ;
        RECT 185.715 177.450 186.775 177.590 ;
        RECT 185.255 176.430 185.855 176.570 ;
        RECT 184.275 175.660 184.535 175.980 ;
        RECT 184.725 119.720 185.005 176.290 ;
        RECT 185.255 174.620 185.395 176.430 ;
        RECT 185.715 176.290 185.855 176.430 ;
        RECT 186.635 176.290 186.775 177.450 ;
        RECT 187.095 176.660 187.235 178.040 ;
        RECT 187.035 176.340 187.295 176.660 ;
        RECT 187.555 176.290 187.695 179.150 ;
        RECT 188.015 178.360 188.155 184.160 ;
        RECT 187.955 178.040 188.215 178.360 ;
        RECT 188.475 176.290 188.615 186.540 ;
        RECT 188.935 186.180 189.075 187.310 ;
        RECT 190.715 187.310 191.375 187.450 ;
        RECT 190.715 187.220 190.975 187.310 ;
        RECT 189.335 186.880 189.595 187.200 ;
        RECT 188.875 185.860 189.135 186.180 ;
        RECT 188.935 184.335 189.075 185.860 ;
        RECT 188.865 183.965 189.145 184.335 ;
        RECT 188.935 183.800 189.075 183.965 ;
        RECT 189.395 183.800 189.535 186.880 ;
        RECT 189.795 186.540 190.055 186.860 ;
        RECT 188.875 183.480 189.135 183.800 ;
        RECT 189.335 183.480 189.595 183.800 ;
        RECT 189.335 181.100 189.595 181.420 ;
        RECT 189.395 176.290 189.535 181.100 ;
        RECT 189.855 180.650 189.995 186.540 ;
        RECT 191.695 186.260 191.835 188.580 ;
        RECT 193.075 187.480 195.055 187.620 ;
        RECT 192.095 186.540 192.355 186.860 ;
        RECT 192.545 186.685 192.825 187.055 ;
        RECT 192.555 186.540 192.815 186.685 ;
        RECT 191.235 186.120 191.835 186.260 ;
        RECT 190.255 183.140 190.515 183.460 ;
        RECT 190.715 183.140 190.975 183.460 ;
        RECT 190.315 182.100 190.455 183.140 ;
        RECT 190.255 181.780 190.515 182.100 ;
        RECT 189.855 180.510 190.455 180.650 ;
        RECT 189.785 179.885 190.065 180.255 ;
        RECT 189.855 179.040 189.995 179.885 ;
        RECT 189.795 178.720 190.055 179.040 ;
        RECT 190.315 176.290 190.455 180.510 ;
        RECT 190.775 180.255 190.915 183.140 ;
        RECT 190.705 179.885 190.985 180.255 ;
        RECT 190.715 178.040 190.975 178.360 ;
        RECT 191.235 178.215 191.375 186.120 ;
        RECT 191.635 185.520 191.895 185.840 ;
        RECT 191.695 184.480 191.835 185.520 ;
        RECT 191.635 184.160 191.895 184.480 ;
        RECT 191.635 183.480 191.895 183.800 ;
        RECT 191.695 181.615 191.835 183.480 ;
        RECT 191.625 181.245 191.905 181.615 ;
        RECT 192.155 179.380 192.295 186.540 ;
        RECT 192.545 183.965 192.825 184.335 ;
        RECT 192.615 183.800 192.755 183.965 ;
        RECT 192.555 183.480 192.815 183.800 ;
        RECT 192.555 182.975 192.815 183.120 ;
        RECT 192.545 182.605 192.825 182.975 ;
        RECT 192.555 180.760 192.815 181.080 ;
        RECT 192.095 179.060 192.355 179.380 ;
        RECT 191.625 178.525 191.905 178.895 ;
        RECT 192.615 178.700 192.755 180.760 ;
        RECT 190.775 177.590 190.915 178.040 ;
        RECT 191.165 177.845 191.445 178.215 ;
        RECT 191.695 177.590 191.835 178.525 ;
        RECT 192.555 178.380 192.815 178.700 ;
        RECT 190.775 177.450 191.835 177.590 ;
        RECT 190.775 176.430 191.375 176.570 ;
        RECT 185.195 174.300 185.455 174.620 ;
        RECT 185.645 120.300 185.925 176.290 ;
        RECT 186.565 120.880 186.845 176.290 ;
        RECT 187.485 121.460 187.765 176.290 ;
        RECT 188.405 122.040 188.685 176.290 ;
        RECT 189.325 122.620 189.605 176.290 ;
        RECT 190.245 123.200 190.525 176.290 ;
        RECT 190.775 175.300 190.915 176.430 ;
        RECT 191.235 176.290 191.375 176.430 ;
        RECT 191.695 176.430 192.295 176.570 ;
        RECT 190.715 174.980 190.975 175.300 ;
        RECT 191.165 123.780 191.445 176.290 ;
        RECT 191.695 175.640 191.835 176.430 ;
        RECT 192.155 176.290 192.295 176.430 ;
        RECT 193.075 176.290 193.215 187.480 ;
        RECT 193.475 186.880 193.735 187.200 ;
        RECT 193.535 179.380 193.675 186.880 ;
        RECT 194.915 186.860 195.055 187.480 ;
        RECT 194.855 186.540 195.115 186.860 ;
        RECT 195.315 186.540 195.575 186.860 ;
        RECT 194.395 186.200 194.655 186.520 ;
        RECT 193.475 179.060 193.735 179.380 ;
        RECT 194.455 179.040 194.595 186.200 ;
        RECT 194.855 184.160 195.115 184.480 ;
        RECT 195.375 184.335 195.515 186.540 ;
        RECT 195.775 185.860 196.035 186.180 ;
        RECT 195.835 184.480 195.975 185.860 ;
        RECT 194.395 178.720 194.655 179.040 ;
        RECT 194.915 178.360 195.055 184.160 ;
        RECT 195.305 183.965 195.585 184.335 ;
        RECT 195.775 184.160 196.035 184.480 ;
        RECT 195.315 183.655 195.575 183.800 ;
        RECT 195.305 183.285 195.585 183.655 ;
        RECT 196.295 183.540 196.435 190.960 ;
        RECT 197.615 189.600 197.875 189.920 ;
        RECT 197.155 188.580 197.415 188.900 ;
        RECT 196.695 188.240 196.955 188.560 ;
        RECT 196.755 187.200 196.895 188.240 ;
        RECT 197.215 187.200 197.355 188.580 ;
        RECT 196.695 186.880 196.955 187.200 ;
        RECT 197.155 186.880 197.415 187.200 ;
        RECT 197.675 186.860 197.815 189.600 ;
        RECT 198.075 188.240 198.335 188.560 ;
        RECT 197.615 186.540 197.875 186.860 ;
        RECT 196.695 186.200 196.955 186.520 ;
        RECT 195.835 183.400 196.435 183.540 ;
        RECT 195.315 182.800 195.575 183.120 ;
        RECT 194.855 178.040 195.115 178.360 ;
        RECT 193.935 177.360 194.195 177.680 ;
        RECT 195.375 177.590 195.515 182.800 ;
        RECT 195.835 179.380 195.975 183.400 ;
        RECT 196.235 182.800 196.495 183.120 ;
        RECT 195.775 179.060 196.035 179.380 ;
        RECT 196.295 178.360 196.435 182.800 ;
        RECT 196.235 178.040 196.495 178.360 ;
        RECT 195.775 177.700 196.035 178.020 ;
        RECT 194.915 177.450 195.515 177.590 ;
        RECT 193.995 176.290 194.135 177.360 ;
        RECT 194.915 176.290 195.055 177.450 ;
        RECT 195.835 176.290 195.975 177.700 ;
        RECT 196.755 176.290 196.895 186.200 ;
        RECT 197.615 185.520 197.875 185.840 ;
        RECT 197.675 184.820 197.815 185.520 ;
        RECT 197.615 184.500 197.875 184.820 ;
        RECT 197.155 184.160 197.415 184.480 ;
        RECT 197.215 183.460 197.355 184.160 ;
        RECT 197.155 183.140 197.415 183.460 ;
        RECT 197.615 183.140 197.875 183.460 ;
        RECT 197.675 176.290 197.815 183.140 ;
        RECT 198.135 176.660 198.275 188.240 ;
        RECT 198.595 187.540 198.735 191.980 ;
        RECT 198.535 187.220 198.795 187.540 ;
        RECT 198.535 185.520 198.795 185.840 ;
        RECT 198.595 184.140 198.735 185.520 ;
        RECT 199.515 184.140 199.655 194.700 ;
        RECT 204.575 192.980 204.715 199.800 ;
        RECT 205.435 194.020 205.695 194.340 ;
        RECT 204.515 192.660 204.775 192.980 ;
        RECT 202.675 190.960 202.935 191.280 ;
        RECT 202.735 189.775 202.875 190.960 ;
        RECT 202.665 189.405 202.945 189.775 ;
        RECT 204.975 185.860 205.235 186.180 ;
        RECT 204.055 185.520 204.315 185.840 ;
        RECT 198.535 183.820 198.795 184.140 ;
        RECT 199.455 183.820 199.715 184.140 ;
        RECT 201.755 183.030 202.015 183.120 ;
        RECT 200.895 182.890 202.015 183.030 ;
        RECT 200.895 181.760 201.035 182.890 ;
        RECT 201.755 182.800 202.015 182.890 ;
        RECT 201.815 182.040 203.335 182.180 ;
        RECT 201.815 181.760 201.955 182.040 ;
        RECT 200.835 181.440 201.095 181.760 ;
        RECT 201.755 181.440 202.015 181.760 ;
        RECT 198.535 181.100 198.795 181.420 ;
        RECT 202.215 181.100 202.475 181.420 ;
        RECT 198.075 176.340 198.335 176.660 ;
        RECT 198.595 176.290 198.735 181.100 ;
        RECT 201.755 180.760 202.015 181.080 ;
        RECT 200.835 180.420 201.095 180.740 ;
        RECT 200.895 179.380 201.035 180.420 ;
        RECT 200.835 179.060 201.095 179.380 ;
        RECT 198.995 178.270 199.255 178.360 ;
        RECT 198.995 178.130 199.655 178.270 ;
        RECT 198.995 178.040 199.255 178.130 ;
        RECT 199.515 176.290 199.655 178.130 ;
        RECT 200.375 178.040 200.635 178.360 ;
        RECT 201.295 178.040 201.555 178.360 ;
        RECT 200.435 176.290 200.575 178.040 ;
        RECT 201.355 176.290 201.495 178.040 ;
        RECT 201.815 177.680 201.955 180.760 ;
        RECT 201.755 177.360 202.015 177.680 ;
        RECT 202.275 176.290 202.415 181.100 ;
        RECT 202.675 177.360 202.935 177.680 ;
        RECT 202.735 176.660 202.875 177.360 ;
        RECT 202.675 176.340 202.935 176.660 ;
        RECT 203.195 176.290 203.335 182.040 ;
        RECT 204.115 181.420 204.255 185.520 ;
        RECT 204.515 183.480 204.775 183.800 ;
        RECT 204.055 181.100 204.315 181.420 ;
        RECT 204.055 180.420 204.315 180.740 ;
        RECT 204.115 176.290 204.255 180.420 ;
        RECT 204.575 179.040 204.715 183.480 ;
        RECT 205.035 181.760 205.175 185.860 ;
        RECT 204.975 181.440 205.235 181.760 ;
        RECT 204.515 178.720 204.775 179.040 ;
        RECT 205.495 178.700 205.635 194.020 ;
        RECT 211.415 191.640 211.675 191.960 ;
        RECT 211.475 189.580 211.615 191.640 ;
        RECT 214.235 190.260 214.375 199.800 ;
        RECT 220.945 198.585 222.485 198.955 ;
        RECT 217.645 195.865 219.185 196.235 ;
        RECT 220.945 193.145 222.485 193.515 ;
        RECT 217.645 190.425 219.185 190.795 ;
        RECT 223.895 190.260 224.035 199.800 ;
        RECT 214.175 189.940 214.435 190.260 ;
        RECT 223.835 189.940 224.095 190.260 ;
        RECT 229.355 189.940 229.615 190.260 ;
        RECT 226.595 189.600 226.855 189.920 ;
        RECT 228.435 189.600 228.695 189.920 ;
        RECT 207.735 189.260 207.995 189.580 ;
        RECT 211.415 189.260 211.675 189.580 ;
        RECT 207.795 186.940 207.935 189.260 ;
        RECT 220.155 188.920 220.415 189.240 ;
        RECT 225.675 188.920 225.935 189.240 ;
        RECT 208.195 188.580 208.455 188.900 ;
        RECT 208.255 187.540 208.395 188.580 ;
        RECT 208.195 187.220 208.455 187.540 ;
        RECT 209.115 187.220 209.375 187.540 ;
        RECT 206.815 186.540 207.075 186.860 ;
        RECT 207.335 186.800 207.935 186.940 ;
        RECT 206.355 184.160 206.615 184.480 ;
        RECT 206.415 180.740 206.555 184.160 ;
        RECT 206.355 180.420 206.615 180.740 ;
        RECT 205.435 178.380 205.695 178.700 ;
        RECT 204.975 177.360 205.235 177.680 ;
        RECT 205.035 176.290 205.175 177.360 ;
        RECT 205.955 176.600 206.555 176.740 ;
        RECT 205.955 176.290 206.095 176.600 ;
        RECT 206.415 176.320 206.555 176.600 ;
        RECT 191.635 175.320 191.895 175.640 ;
        RECT 192.085 124.360 192.365 176.290 ;
        RECT 193.005 124.940 193.285 176.290 ;
        RECT 193.925 125.520 194.205 176.290 ;
        RECT 194.845 126.100 195.125 176.290 ;
        RECT 195.765 126.680 196.045 176.290 ;
        RECT 196.685 127.260 196.965 176.290 ;
        RECT 197.605 127.840 197.885 176.290 ;
        RECT 198.525 128.420 198.805 176.290 ;
        RECT 199.445 129.000 199.725 176.290 ;
        RECT 200.365 129.580 200.645 176.290 ;
        RECT 201.285 130.160 201.565 176.290 ;
        RECT 202.205 130.740 202.485 176.290 ;
        RECT 203.125 131.320 203.405 176.290 ;
        RECT 204.045 131.900 204.325 176.290 ;
        RECT 204.965 132.480 205.245 176.290 ;
        RECT 205.885 133.060 206.165 176.290 ;
        RECT 206.355 176.000 206.615 176.320 ;
        RECT 206.875 176.290 207.015 186.540 ;
        RECT 207.335 184.480 207.475 186.800 ;
        RECT 208.185 186.685 208.465 187.055 ;
        RECT 208.255 186.260 208.395 186.685 ;
        RECT 208.655 186.540 208.915 186.860 ;
        RECT 207.795 186.180 208.395 186.260 ;
        RECT 207.735 186.120 208.395 186.180 ;
        RECT 207.735 185.860 207.995 186.120 ;
        RECT 208.195 185.520 208.455 185.840 ;
        RECT 207.725 184.645 208.005 185.015 ;
        RECT 207.275 184.160 207.535 184.480 ;
        RECT 207.275 182.975 207.535 183.120 ;
        RECT 207.265 182.605 207.545 182.975 ;
        RECT 207.275 178.380 207.535 178.700 ;
        RECT 206.805 133.640 207.085 176.290 ;
        RECT 207.335 174.620 207.475 178.380 ;
        RECT 207.795 176.290 207.935 184.645 ;
        RECT 208.255 184.140 208.395 185.520 ;
        RECT 208.715 185.015 208.855 186.540 ;
        RECT 208.645 184.645 208.925 185.015 ;
        RECT 208.195 183.820 208.455 184.140 ;
        RECT 209.175 183.655 209.315 187.220 ;
        RECT 210.955 186.770 211.215 186.860 ;
        RECT 209.635 186.630 211.215 186.770 ;
        RECT 208.185 183.285 208.465 183.655 ;
        RECT 209.105 183.285 209.385 183.655 ;
        RECT 208.255 178.700 208.395 183.285 ;
        RECT 209.115 182.800 209.375 183.120 ;
        RECT 208.655 181.100 208.915 181.420 ;
        RECT 209.175 181.340 209.315 182.800 ;
        RECT 208.715 180.650 208.855 181.100 ;
        RECT 209.115 181.020 209.375 181.340 ;
        RECT 208.715 180.510 209.315 180.650 ;
        RECT 208.645 179.885 208.925 180.255 ;
        RECT 208.195 178.380 208.455 178.700 ;
        RECT 208.715 176.290 208.855 179.885 ;
        RECT 209.175 178.895 209.315 180.510 ;
        RECT 209.105 178.525 209.385 178.895 ;
        RECT 209.635 176.290 209.775 186.630 ;
        RECT 210.955 186.540 211.215 186.630 ;
        RECT 211.875 186.540 212.135 186.860 ;
        RECT 216.475 186.540 216.735 186.860 ;
        RECT 219.695 186.540 219.955 186.860 ;
        RECT 210.495 185.860 210.755 186.180 ;
        RECT 210.555 185.695 210.695 185.860 ;
        RECT 210.485 185.325 210.765 185.695 ;
        RECT 210.495 183.655 210.755 183.800 ;
        RECT 210.485 183.285 210.765 183.655 ;
        RECT 211.415 183.480 211.675 183.800 ;
        RECT 211.475 182.860 211.615 183.480 ;
        RECT 211.015 182.720 211.615 182.860 ;
        RECT 210.035 181.330 210.295 181.420 ;
        RECT 211.015 181.330 211.155 182.720 ;
        RECT 211.935 182.010 212.075 186.540 ;
        RECT 212.795 186.200 213.055 186.520 ;
        RECT 210.035 181.190 211.155 181.330 ;
        RECT 210.035 181.100 210.295 181.190 ;
        RECT 210.035 180.080 210.295 180.400 ;
        RECT 210.095 179.040 210.235 180.080 ;
        RECT 210.485 179.205 210.765 179.575 ;
        RECT 210.035 178.720 210.295 179.040 ;
        RECT 210.555 176.290 210.695 179.205 ;
        RECT 211.015 177.535 211.155 181.190 ;
        RECT 211.475 181.870 212.075 182.010 ;
        RECT 210.945 177.165 211.225 177.535 ;
        RECT 207.275 174.300 207.535 174.620 ;
        RECT 207.725 134.220 208.005 176.290 ;
        RECT 208.645 134.800 208.925 176.290 ;
        RECT 209.565 135.380 209.845 176.290 ;
        RECT 210.485 135.960 210.765 176.290 ;
        RECT 211.015 174.620 211.155 177.165 ;
        RECT 211.475 176.290 211.615 181.870 ;
        RECT 212.335 181.780 212.595 182.100 ;
        RECT 211.865 181.245 212.145 181.615 ;
        RECT 211.935 178.700 212.075 181.245 ;
        RECT 212.395 178.700 212.535 181.780 ;
        RECT 211.875 178.380 212.135 178.700 ;
        RECT 212.335 178.380 212.595 178.700 ;
        RECT 212.855 178.100 212.995 186.200 ;
        RECT 214.175 185.860 214.435 186.180 ;
        RECT 214.625 186.005 214.905 186.375 ;
        RECT 213.255 185.520 213.515 185.840 ;
        RECT 213.315 178.700 213.455 185.520 ;
        RECT 213.705 181.925 213.985 182.295 ;
        RECT 213.715 181.780 213.975 181.925 ;
        RECT 214.235 181.420 214.375 185.860 ;
        RECT 214.695 184.820 214.835 186.005 ;
        RECT 215.095 185.520 215.355 185.840 ;
        RECT 215.555 185.520 215.815 185.840 ;
        RECT 214.635 184.500 214.895 184.820 ;
        RECT 214.635 183.480 214.895 183.800 ;
        RECT 214.175 181.100 214.435 181.420 ;
        RECT 213.715 180.760 213.975 181.080 ;
        RECT 213.255 178.380 213.515 178.700 ;
        RECT 212.395 177.960 212.995 178.100 ;
        RECT 212.395 176.290 212.535 177.960 ;
        RECT 213.775 177.590 213.915 180.760 ;
        RECT 214.695 179.575 214.835 183.480 ;
        RECT 214.625 179.205 214.905 179.575 ;
        RECT 215.155 178.700 215.295 185.520 ;
        RECT 215.615 183.120 215.755 185.520 ;
        RECT 216.535 184.820 216.675 186.540 ;
        RECT 216.935 186.200 217.195 186.520 ;
        RECT 216.475 184.500 216.735 184.820 ;
        RECT 216.015 183.820 216.275 184.140 ;
        RECT 216.475 183.820 216.735 184.140 ;
        RECT 215.555 182.800 215.815 183.120 ;
        RECT 216.075 182.100 216.215 183.820 ;
        RECT 216.015 181.780 216.275 182.100 ;
        RECT 216.005 180.565 216.285 180.935 ;
        RECT 215.555 180.080 215.815 180.400 ;
        RECT 215.095 178.380 215.355 178.700 ;
        RECT 214.165 177.845 214.445 178.215 ;
        RECT 214.635 178.040 214.895 178.360 ;
        RECT 212.855 177.450 213.915 177.590 ;
        RECT 212.855 176.660 212.995 177.450 ;
        RECT 212.795 176.340 213.055 176.660 ;
        RECT 213.315 176.430 213.915 176.570 ;
        RECT 213.315 176.290 213.455 176.430 ;
        RECT 210.955 174.300 211.215 174.620 ;
        RECT 211.405 136.540 211.685 176.290 ;
        RECT 212.325 137.120 212.605 176.290 ;
        RECT 213.245 137.700 213.525 176.290 ;
        RECT 213.775 175.300 213.915 176.430 ;
        RECT 214.235 176.290 214.375 177.845 ;
        RECT 214.695 176.320 214.835 178.040 ;
        RECT 215.615 177.680 215.755 180.080 ;
        RECT 216.075 178.215 216.215 180.565 ;
        RECT 216.535 179.380 216.675 183.820 ;
        RECT 216.475 179.060 216.735 179.380 ;
        RECT 216.005 177.845 216.285 178.215 ;
        RECT 215.555 177.360 215.815 177.680 ;
        RECT 215.155 176.430 215.755 176.570 ;
        RECT 213.715 174.980 213.975 175.300 ;
        RECT 214.165 138.280 214.445 176.290 ;
        RECT 214.635 176.000 214.895 176.320 ;
        RECT 215.155 176.290 215.295 176.430 ;
        RECT 215.085 138.860 215.365 176.290 ;
        RECT 215.615 175.640 215.755 176.430 ;
        RECT 216.075 176.430 216.675 176.570 ;
        RECT 216.075 176.290 216.215 176.430 ;
        RECT 215.555 175.320 215.815 175.640 ;
        RECT 216.005 139.440 216.285 176.290 ;
        RECT 216.535 175.980 216.675 176.430 ;
        RECT 216.995 176.290 217.135 186.200 ;
        RECT 217.645 184.985 219.185 185.355 ;
        RECT 219.755 184.820 219.895 186.540 ;
        RECT 220.215 184.820 220.355 188.920 ;
        RECT 222.915 188.240 223.175 188.560 ;
        RECT 220.945 187.705 222.485 188.075 ;
        RECT 221.995 187.220 222.255 187.540 ;
        RECT 221.075 185.860 221.335 186.180 ;
        RECT 217.395 184.500 217.655 184.820 ;
        RECT 217.855 184.500 218.115 184.820 ;
        RECT 219.695 184.500 219.955 184.820 ;
        RECT 220.155 184.500 220.415 184.820 ;
        RECT 217.455 180.935 217.595 184.500 ;
        RECT 217.385 180.565 217.665 180.935 ;
        RECT 217.395 180.310 217.655 180.400 ;
        RECT 217.915 180.310 218.055 184.500 ;
        RECT 221.135 184.220 221.275 185.860 ;
        RECT 222.055 184.390 222.195 187.220 ;
        RECT 220.215 184.140 221.275 184.220 ;
        RECT 219.695 183.820 219.955 184.140 ;
        RECT 220.155 184.080 221.275 184.140 ;
        RECT 221.595 184.250 222.195 184.390 ;
        RECT 220.155 183.820 220.415 184.080 ;
        RECT 219.755 181.500 219.895 183.820 ;
        RECT 220.215 182.975 220.355 183.820 ;
        RECT 221.595 183.800 221.735 184.250 ;
        RECT 222.975 184.220 223.115 188.240 ;
        RECT 225.735 188.160 225.875 188.920 ;
        RECT 226.135 188.580 226.395 188.900 ;
        RECT 225.275 188.020 225.875 188.160 ;
        RECT 224.745 186.685 225.025 187.055 ;
        RECT 222.515 184.080 223.115 184.220 ;
        RECT 221.535 183.480 221.795 183.800 ;
        RECT 222.515 183.030 222.655 184.080 ;
        RECT 222.915 183.710 223.175 183.800 ;
        RECT 222.915 183.570 224.035 183.710 ;
        RECT 222.915 183.480 223.175 183.570 ;
        RECT 220.145 182.605 220.425 182.975 ;
        RECT 222.515 182.890 223.115 183.030 ;
        RECT 220.215 182.180 220.355 182.605 ;
        RECT 220.945 182.265 222.485 182.635 ;
        RECT 220.215 182.040 220.815 182.180 ;
        RECT 219.755 181.360 220.355 181.500 ;
        RECT 218.775 180.935 219.035 181.080 ;
        RECT 218.765 180.565 219.045 180.935 ;
        RECT 219.695 180.760 219.955 181.080 ;
        RECT 217.395 180.170 218.055 180.310 ;
        RECT 217.395 180.080 217.655 180.170 ;
        RECT 217.645 179.545 219.185 179.915 ;
        RECT 219.755 179.380 219.895 180.760 ;
        RECT 220.215 180.255 220.355 181.360 ;
        RECT 220.145 179.885 220.425 180.255 ;
        RECT 219.695 179.060 219.955 179.380 ;
        RECT 220.675 179.040 220.815 182.040 ;
        RECT 222.975 182.010 223.115 182.890 ;
        RECT 223.375 182.800 223.635 183.120 ;
        RECT 223.895 183.030 224.035 183.570 ;
        RECT 224.295 183.030 224.555 183.120 ;
        RECT 223.895 182.890 224.555 183.030 ;
        RECT 221.595 181.870 223.115 182.010 ;
        RECT 221.075 180.760 221.335 181.080 ;
        RECT 220.615 178.720 220.875 179.040 ;
        RECT 221.135 178.270 221.275 180.760 ;
        RECT 221.595 178.700 221.735 181.870 ;
        RECT 223.435 181.420 223.575 182.800 ;
        RECT 223.375 181.100 223.635 181.420 ;
        RECT 223.895 180.990 224.035 182.890 ;
        RECT 224.295 182.800 224.555 182.890 ;
        RECT 224.815 181.080 224.955 186.685 ;
        RECT 224.295 180.990 224.555 181.080 ;
        RECT 223.895 180.850 224.555 180.990 ;
        RECT 224.295 180.760 224.555 180.850 ;
        RECT 224.755 180.760 225.015 181.080 ;
        RECT 222.905 179.885 223.185 180.255 ;
        RECT 223.375 180.080 223.635 180.400 ;
        RECT 223.835 180.080 224.095 180.400 ;
        RECT 222.975 178.780 223.115 179.885 ;
        RECT 223.435 179.575 223.575 180.080 ;
        RECT 223.365 179.205 223.645 179.575 ;
        RECT 221.535 178.380 221.795 178.700 ;
        RECT 222.975 178.640 223.575 178.780 ;
        RECT 219.685 177.845 219.965 178.215 ;
        RECT 220.675 178.130 221.275 178.270 ;
        RECT 217.915 177.280 219.435 177.420 ;
        RECT 217.915 176.290 218.055 177.280 ;
        RECT 218.375 176.600 218.975 176.740 ;
        RECT 219.295 176.660 219.435 177.280 ;
        RECT 218.375 176.320 218.515 176.600 ;
        RECT 216.475 175.660 216.735 175.980 ;
        RECT 216.925 140.020 217.205 176.290 ;
        RECT 217.845 140.600 218.125 176.290 ;
        RECT 218.315 176.000 218.575 176.320 ;
        RECT 218.835 176.290 218.975 176.600 ;
        RECT 219.235 176.340 219.495 176.660 ;
        RECT 219.755 176.290 219.895 177.845 ;
        RECT 220.145 177.420 220.425 177.535 ;
        RECT 220.675 177.420 220.815 178.130 ;
        RECT 221.135 178.100 221.275 178.130 ;
        RECT 222.915 178.100 223.175 178.360 ;
        RECT 221.135 178.040 223.175 178.100 ;
        RECT 221.135 177.960 223.115 178.040 ;
        RECT 223.435 177.680 223.575 178.640 ;
        RECT 220.145 177.280 220.815 177.420 ;
        RECT 223.375 177.360 223.635 177.680 ;
        RECT 220.145 177.165 220.425 177.280 ;
        RECT 220.945 176.825 222.485 177.195 ;
        RECT 222.905 176.570 223.185 176.855 ;
        RECT 223.895 176.570 224.035 180.080 ;
        RECT 224.285 179.205 224.565 179.575 ;
        RECT 220.675 176.430 221.275 176.570 ;
        RECT 220.675 176.290 220.815 176.430 ;
        RECT 218.765 141.180 219.045 176.290 ;
        RECT 219.685 141.760 219.965 176.290 ;
        RECT 220.605 142.340 220.885 176.290 ;
        RECT 221.135 174.960 221.275 176.430 ;
        RECT 221.595 176.430 222.195 176.570 ;
        RECT 221.595 176.290 221.735 176.430 ;
        RECT 221.075 174.640 221.335 174.960 ;
        RECT 221.525 142.920 221.805 176.290 ;
        RECT 222.055 176.175 222.195 176.430 ;
        RECT 222.515 176.485 223.185 176.570 ;
        RECT 222.515 176.430 223.115 176.485 ;
        RECT 223.435 176.430 224.035 176.570 ;
        RECT 222.515 176.290 222.655 176.430 ;
        RECT 223.435 176.290 223.575 176.430 ;
        RECT 224.355 176.290 224.495 179.205 ;
        RECT 225.275 176.290 225.415 188.020 ;
        RECT 225.675 186.200 225.935 186.520 ;
        RECT 225.735 184.820 225.875 186.200 ;
        RECT 225.675 184.500 225.935 184.820 ;
        RECT 225.675 183.140 225.935 183.460 ;
        RECT 225.735 180.400 225.875 183.140 ;
        RECT 225.675 180.080 225.935 180.400 ;
        RECT 226.195 176.290 226.335 188.580 ;
        RECT 226.655 179.380 226.795 189.600 ;
        RECT 227.055 186.200 227.315 186.520 ;
        RECT 227.975 186.200 228.235 186.520 ;
        RECT 227.115 183.120 227.255 186.200 ;
        RECT 228.035 184.220 228.175 186.200 ;
        RECT 227.575 184.080 228.175 184.220 ;
        RECT 227.055 182.800 227.315 183.120 ;
        RECT 227.045 179.885 227.325 180.255 ;
        RECT 226.595 179.060 226.855 179.380 ;
        RECT 226.595 178.040 226.855 178.360 ;
        RECT 221.985 175.805 222.265 176.175 ;
        RECT 222.445 143.500 222.725 176.290 ;
        RECT 223.365 144.080 223.645 176.290 ;
        RECT 224.285 144.660 224.565 176.290 ;
        RECT 225.205 145.240 225.485 176.290 ;
        RECT 226.125 145.820 226.405 176.290 ;
        RECT 226.655 175.300 226.795 178.040 ;
        RECT 227.115 176.290 227.255 179.885 ;
        RECT 227.575 177.590 227.715 184.080 ;
        RECT 227.975 183.480 228.235 183.800 ;
        RECT 228.035 178.215 228.175 183.480 ;
        RECT 228.495 181.340 228.635 189.600 ;
        RECT 228.895 188.240 229.155 188.560 ;
        RECT 228.955 185.840 229.095 188.240 ;
        RECT 229.415 187.540 229.555 189.940 ;
        RECT 229.815 189.260 230.075 189.580 ;
        RECT 229.355 187.220 229.615 187.540 ;
        RECT 229.875 186.860 230.015 189.260 ;
        RECT 230.735 188.920 230.995 189.240 ;
        RECT 229.815 186.540 230.075 186.860 ;
        RECT 228.895 185.520 229.155 185.840 ;
        RECT 230.275 185.520 230.535 185.840 ;
        RECT 230.335 184.820 230.475 185.520 ;
        RECT 230.275 184.500 230.535 184.820 ;
        RECT 228.885 183.285 229.165 183.655 ;
        RECT 230.275 183.480 230.535 183.800 ;
        RECT 228.435 181.020 228.695 181.340 ;
        RECT 228.955 179.380 229.095 183.285 ;
        RECT 229.815 182.800 230.075 183.120 ;
        RECT 229.355 180.760 229.615 181.080 ;
        RECT 229.415 179.380 229.555 180.760 ;
        RECT 228.895 179.060 229.155 179.380 ;
        RECT 229.355 179.060 229.615 179.380 ;
        RECT 229.875 178.895 230.015 182.800 ;
        RECT 229.805 178.525 230.085 178.895 ;
        RECT 227.965 177.845 228.245 178.215 ;
        RECT 229.355 178.040 229.615 178.360 ;
        RECT 227.575 177.450 228.175 177.590 ;
        RECT 228.035 176.290 228.175 177.450 ;
        RECT 226.595 174.980 226.855 175.300 ;
        RECT 227.045 146.400 227.325 176.290 ;
        RECT 227.965 146.980 228.245 176.290 ;
        RECT 229.415 175.640 229.555 178.040 ;
        RECT 230.335 176.175 230.475 183.480 ;
        RECT 230.795 180.255 230.935 188.920 ;
        RECT 233.095 187.540 233.235 199.800 ;
        RECT 233.035 187.220 233.295 187.540 ;
        RECT 231.195 186.540 231.455 186.860 ;
        RECT 231.255 184.335 231.395 186.540 ;
        RECT 231.185 183.965 231.465 184.335 ;
        RECT 231.655 183.820 231.915 184.140 ;
        RECT 231.195 182.800 231.455 183.120 ;
        RECT 231.255 180.935 231.395 182.800 ;
        RECT 231.185 180.565 231.465 180.935 ;
        RECT 230.725 179.885 231.005 180.255 ;
        RECT 230.735 178.040 230.995 178.360 ;
        RECT 230.265 175.805 230.545 176.175 ;
        RECT 230.795 175.980 230.935 178.040 ;
        RECT 230.735 175.660 230.995 175.980 ;
        RECT 229.355 175.320 229.615 175.640 ;
        RECT 231.715 174.960 231.855 183.820 ;
        RECT 233.495 183.480 233.755 183.800 ;
        RECT 232.575 182.800 232.835 183.120 ;
        RECT 232.635 181.615 232.775 182.800 ;
        RECT 232.565 181.245 232.845 181.615 ;
        RECT 233.035 180.080 233.295 180.400 ;
        RECT 232.115 178.040 232.375 178.360 ;
        RECT 232.175 176.660 232.315 178.040 ;
        RECT 232.115 176.340 232.375 176.660 ;
        RECT 231.655 174.640 231.915 174.960 ;
        RECT 233.095 174.815 233.235 180.080 ;
        RECT 233.555 179.575 233.695 183.480 ;
        RECT 234.415 181.100 234.675 181.420 ;
        RECT 233.485 179.205 233.765 179.575 ;
        RECT 233.495 178.040 233.755 178.360 ;
        RECT 233.555 176.320 233.695 178.040 ;
        RECT 234.475 176.855 234.615 181.100 ;
        RECT 234.405 176.485 234.685 176.855 ;
        RECT 233.495 176.000 233.755 176.320 ;
        RECT 233.025 174.445 233.305 174.815 ;
        RECT 227.965 146.700 309.205 146.980 ;
        RECT 227.045 146.120 306.905 146.400 ;
        RECT 226.125 145.540 304.605 145.820 ;
        RECT 225.205 144.960 302.305 145.240 ;
        RECT 224.285 144.380 300.005 144.660 ;
        RECT 223.365 143.800 297.705 144.080 ;
        RECT 222.445 143.220 295.405 143.500 ;
        RECT 221.525 142.640 293.105 142.920 ;
        RECT 220.605 142.060 290.805 142.340 ;
        RECT 219.685 141.480 288.505 141.760 ;
        RECT 218.765 140.900 286.205 141.180 ;
        RECT 217.845 140.320 283.905 140.600 ;
        RECT 216.925 139.740 281.605 140.020 ;
        RECT 216.005 139.160 279.305 139.440 ;
        RECT 215.085 138.580 277.005 138.860 ;
        RECT 214.165 138.000 274.705 138.280 ;
        RECT 213.245 137.420 272.405 137.700 ;
        RECT 212.325 136.840 270.105 137.120 ;
        RECT 211.405 136.260 267.805 136.540 ;
        RECT 210.485 135.680 265.505 135.960 ;
        RECT 209.565 135.100 263.205 135.380 ;
        RECT 208.645 134.520 260.905 134.800 ;
        RECT 207.725 133.940 258.605 134.220 ;
        RECT 206.805 133.360 256.305 133.640 ;
        RECT 205.885 132.780 254.005 133.060 ;
        RECT 204.965 132.200 251.705 132.480 ;
        RECT 204.045 131.620 249.405 131.900 ;
        RECT 203.125 131.040 247.105 131.320 ;
        RECT 202.205 130.460 244.805 130.740 ;
        RECT 201.285 129.880 242.505 130.160 ;
        RECT 200.365 129.300 240.205 129.580 ;
        RECT 199.445 128.720 237.905 129.000 ;
        RECT 198.525 128.140 235.605 128.420 ;
        RECT 197.605 127.560 233.305 127.840 ;
        RECT 196.685 126.980 231.005 127.260 ;
        RECT 195.765 126.400 228.705 126.680 ;
        RECT 194.845 125.820 226.405 126.100 ;
        RECT 193.925 125.240 224.105 125.520 ;
        RECT 193.005 124.660 221.805 124.940 ;
        RECT 192.085 124.080 219.505 124.360 ;
        RECT 191.165 123.500 217.205 123.780 ;
        RECT 190.245 122.920 214.905 123.200 ;
        RECT 189.325 122.340 212.605 122.620 ;
        RECT 188.405 121.760 210.305 122.040 ;
        RECT 187.485 121.180 208.005 121.460 ;
        RECT 186.565 120.600 205.705 120.880 ;
        RECT 185.645 120.020 203.405 120.300 ;
        RECT 184.725 119.440 201.105 119.720 ;
        RECT 183.805 118.860 198.805 119.140 ;
        RECT 182.885 118.280 196.505 118.560 ;
        RECT 181.965 117.700 194.205 117.980 ;
        RECT 181.045 117.120 191.905 117.400 ;
        RECT 180.125 116.540 189.605 116.820 ;
        RECT 179.205 115.960 187.305 116.240 ;
        RECT 178.285 115.380 185.005 115.660 ;
        RECT 177.365 114.800 182.705 115.080 ;
        RECT 176.445 114.220 180.405 114.500 ;
        RECT 175.525 113.410 178.105 113.690 ;
        RECT 174.605 112.685 175.805 112.965 ;
        RECT 173.225 109.225 173.505 112.685 ;
        RECT 175.525 109.225 175.805 112.685 ;
        RECT 177.825 109.225 178.105 113.410 ;
        RECT 180.125 109.225 180.405 114.220 ;
        RECT 182.425 109.225 182.705 114.800 ;
        RECT 184.725 109.225 185.005 115.380 ;
        RECT 187.025 109.225 187.305 115.960 ;
        RECT 189.325 109.225 189.605 116.540 ;
        RECT 191.625 109.225 191.905 117.120 ;
        RECT 193.925 109.225 194.205 117.700 ;
        RECT 196.225 109.225 196.505 118.280 ;
        RECT 198.525 109.225 198.805 118.860 ;
        RECT 200.825 109.225 201.105 119.440 ;
        RECT 203.125 109.225 203.405 120.020 ;
        RECT 205.425 109.225 205.705 120.600 ;
        RECT 207.725 109.225 208.005 121.180 ;
        RECT 210.025 109.225 210.305 121.760 ;
        RECT 212.325 109.225 212.605 122.340 ;
        RECT 214.625 109.225 214.905 122.920 ;
        RECT 216.925 109.225 217.205 123.500 ;
        RECT 219.225 109.225 219.505 124.080 ;
        RECT 221.525 109.225 221.805 124.660 ;
        RECT 223.825 109.225 224.105 125.240 ;
        RECT 226.125 109.225 226.405 125.820 ;
        RECT 228.425 109.225 228.705 126.400 ;
        RECT 230.725 109.225 231.005 126.980 ;
        RECT 233.025 109.225 233.305 127.560 ;
        RECT 235.325 109.225 235.605 128.140 ;
        RECT 235.795 109.495 236.055 109.815 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 164.095 100.635 164.235 109.225 ;
        RECT 164.495 105.075 164.755 105.395 ;
        RECT 164.035 100.315 164.295 100.635 ;
        RECT 164.035 93.350 164.295 93.495 ;
        RECT 164.025 92.980 164.305 93.350 ;
        RECT 146.290 88.455 148.395 92.555 ;
        RECT 146.290 83.775 148.395 87.875 ;
        RECT 146.290 77.925 148.395 83.195 ;
        RECT 146.290 73.245 148.395 77.345 ;
        RECT 146.290 68.565 148.395 72.665 ;
        RECT 164.555 69.355 164.695 105.075 ;
        RECT 165.415 102.015 165.675 102.335 ;
        RECT 165.475 100.715 165.615 102.015 ;
        RECT 165.475 100.575 166.075 100.715 ;
        RECT 166.395 100.635 166.535 109.225 ;
        RECT 167.255 105.075 167.515 105.395 ;
        RECT 166.795 101.675 167.055 101.995 ;
        RECT 164.955 99.635 165.215 99.955 ;
        RECT 165.415 99.635 165.675 99.955 ;
        RECT 165.015 81.595 165.155 99.635 ;
        RECT 165.475 91.795 165.615 99.635 ;
        RECT 165.415 91.475 165.675 91.795 ;
        RECT 165.475 87.035 165.615 91.475 ;
        RECT 165.935 91.115 166.075 100.575 ;
        RECT 166.335 100.315 166.595 100.635 ;
        RECT 166.855 99.955 166.995 101.675 ;
        RECT 166.795 99.635 167.055 99.955 ;
        RECT 166.855 95.195 166.995 99.635 ;
        RECT 166.795 94.875 167.055 95.195 ;
        RECT 165.875 90.795 166.135 91.115 ;
        RECT 165.935 89.755 166.075 90.795 ;
        RECT 165.875 89.435 166.135 89.755 ;
        RECT 165.415 86.715 165.675 87.035 ;
        RECT 164.955 81.275 165.215 81.595 ;
        RECT 164.495 69.035 164.755 69.355 ;
        RECT 146.290 63.885 148.395 67.985 ;
        RECT 164.555 65.275 164.695 69.035 ;
        RECT 167.315 67.995 167.455 105.075 ;
        RECT 168.695 101.655 168.835 109.225 ;
        RECT 169.555 107.455 169.815 107.775 ;
        RECT 169.095 105.075 169.355 105.395 ;
        RECT 168.635 101.335 168.895 101.655 ;
        RECT 168.635 96.235 168.895 96.555 ;
        RECT 168.695 87.115 168.835 96.235 ;
        RECT 168.235 87.035 168.835 87.115 ;
        RECT 168.175 86.975 168.835 87.035 ;
        RECT 168.175 86.715 168.435 86.975 ;
        RECT 168.695 84.315 168.835 86.975 ;
        RECT 168.635 83.995 168.895 84.315 ;
        RECT 167.255 67.675 167.515 67.995 ;
        RECT 164.495 64.955 164.755 65.275 ;
        RECT 169.155 65.185 169.295 105.075 ;
        RECT 169.615 104.375 169.755 107.455 ;
        RECT 169.555 104.055 169.815 104.375 ;
        RECT 170.015 104.055 170.275 104.375 ;
        RECT 170.075 100.295 170.215 104.055 ;
        RECT 170.015 99.975 170.275 100.295 ;
        RECT 170.995 96.215 171.135 109.225 ;
        RECT 173.295 106.075 173.435 109.225 ;
        RECT 173.235 105.755 173.495 106.075 ;
        RECT 173.695 105.075 173.955 105.395 ;
        RECT 173.235 104.735 173.495 105.055 ;
        RECT 170.935 95.895 171.195 96.215 ;
        RECT 173.295 90.775 173.435 104.735 ;
        RECT 173.755 99.470 173.895 105.075 ;
        RECT 175.595 105.055 175.735 109.225 ;
        RECT 177.895 105.735 178.035 109.225 ;
        RECT 178.295 107.115 178.555 107.435 ;
        RECT 177.835 105.415 178.095 105.735 ;
        RECT 175.535 104.735 175.795 105.055 ;
        RECT 177.835 104.795 178.095 105.055 ;
        RECT 178.355 104.795 178.495 107.115 ;
        RECT 176.975 104.655 178.495 104.795 ;
        RECT 175.535 104.055 175.795 104.375 ;
        RECT 175.995 104.055 176.255 104.375 ;
        RECT 175.595 103.355 175.735 104.055 ;
        RECT 175.535 103.035 175.795 103.355 ;
        RECT 176.055 103.015 176.195 104.055 ;
        RECT 175.995 102.695 176.255 103.015 ;
        RECT 174.155 101.675 174.415 101.995 ;
        RECT 174.215 99.955 174.355 101.675 ;
        RECT 174.155 99.635 174.415 99.955 ;
        RECT 173.685 99.100 173.965 99.470 ;
        RECT 174.215 96.555 174.355 99.635 ;
        RECT 175.995 99.470 176.255 99.615 ;
        RECT 175.985 99.100 176.265 99.470 ;
        RECT 176.455 98.615 176.715 98.935 ;
        RECT 176.515 97.915 176.655 98.615 ;
        RECT 176.455 97.595 176.715 97.915 ;
        RECT 174.615 97.255 174.875 97.575 ;
        RECT 174.155 96.235 174.415 96.555 ;
        RECT 174.215 93.495 174.355 96.235 ;
        RECT 173.695 93.175 173.955 93.495 ;
        RECT 174.155 93.175 174.415 93.495 ;
        RECT 173.235 90.455 173.495 90.775 ;
        RECT 173.235 87.735 173.495 88.055 ;
        RECT 173.295 86.355 173.435 87.735 ;
        RECT 173.235 86.035 173.495 86.355 ;
        RECT 173.755 85.755 173.895 93.175 ;
        RECT 174.215 89.415 174.355 93.175 ;
        RECT 174.155 89.095 174.415 89.415 ;
        RECT 171.855 85.355 172.115 85.675 ;
        RECT 173.295 85.615 173.895 85.755 ;
        RECT 171.915 84.315 172.055 85.355 ;
        RECT 171.855 83.995 172.115 84.315 ;
        RECT 172.775 79.915 173.035 80.235 ;
        RECT 172.835 73.630 172.975 79.915 ;
        RECT 172.765 73.260 173.045 73.630 ;
        RECT 172.835 73.095 172.975 73.260 ;
        RECT 172.775 72.775 173.035 73.095 ;
        RECT 172.315 68.695 172.575 69.015 ;
        RECT 172.375 67.995 172.515 68.695 ;
        RECT 172.315 67.675 172.575 67.995 ;
        RECT 172.375 67.510 172.515 67.675 ;
        RECT 172.835 67.655 172.975 72.775 ;
        RECT 173.295 70.715 173.435 85.615 ;
        RECT 174.215 84.315 174.355 89.095 ;
        RECT 174.675 86.355 174.815 97.255 ;
        RECT 175.535 95.895 175.795 96.215 ;
        RECT 176.975 95.955 177.115 104.655 ;
        RECT 179.675 104.395 179.935 104.715 ;
        RECT 177.645 103.520 179.185 103.890 ;
        RECT 179.735 99.615 179.875 104.395 ;
        RECT 180.195 100.635 180.335 109.225 ;
        RECT 182.495 107.515 182.635 109.225 ;
        RECT 182.495 107.375 183.095 107.515 ;
        RECT 180.945 106.240 182.485 106.610 ;
        RECT 181.055 105.475 181.315 105.735 ;
        RECT 180.655 105.415 181.315 105.475 ;
        RECT 180.655 105.335 181.255 105.415 ;
        RECT 180.135 100.315 180.395 100.635 ;
        RECT 180.135 99.635 180.395 99.955 ;
        RECT 179.675 99.295 179.935 99.615 ;
        RECT 177.645 98.080 179.185 98.450 ;
        RECT 179.735 97.235 179.875 99.295 ;
        RECT 179.675 96.915 179.935 97.235 ;
        RECT 180.195 96.555 180.335 99.635 ;
        RECT 180.135 96.235 180.395 96.555 ;
        RECT 175.595 94.175 175.735 95.895 ;
        RECT 176.055 95.815 177.115 95.955 ;
        RECT 177.375 95.895 177.635 96.215 ;
        RECT 180.655 95.955 180.795 105.335 ;
        RECT 180.945 100.800 182.485 101.170 ;
        RECT 182.955 100.635 183.095 107.375 ;
        RECT 184.275 105.075 184.535 105.395 ;
        RECT 182.895 100.315 183.155 100.635 ;
        RECT 182.895 99.635 183.155 99.955 ;
        RECT 183.815 99.635 184.075 99.955 ;
        RECT 182.435 96.750 182.695 96.895 ;
        RECT 182.425 96.380 182.705 96.750 ;
        RECT 175.535 93.855 175.795 94.175 ;
        RECT 175.075 90.455 175.335 90.775 ;
        RECT 175.135 89.755 175.275 90.455 ;
        RECT 175.075 89.435 175.335 89.755 ;
        RECT 174.615 86.035 174.875 86.355 ;
        RECT 174.675 84.315 174.815 86.035 ;
        RECT 176.055 85.675 176.195 95.815 ;
        RECT 177.435 95.195 177.575 95.895 ;
        RECT 180.195 95.815 180.795 95.955 ;
        RECT 176.915 94.875 177.175 95.195 ;
        RECT 177.375 94.875 177.635 95.195 ;
        RECT 176.455 90.455 176.715 90.775 ;
        RECT 176.515 89.415 176.655 90.455 ;
        RECT 176.975 89.415 177.115 94.875 ;
        RECT 177.645 92.640 179.185 93.010 ;
        RECT 178.295 90.455 178.555 90.775 ;
        RECT 176.455 89.095 176.715 89.415 ;
        RECT 176.915 89.095 177.175 89.415 ;
        RECT 175.995 85.355 176.255 85.675 ;
        RECT 175.535 85.015 175.795 85.335 ;
        RECT 174.155 83.995 174.415 84.315 ;
        RECT 174.615 83.995 174.875 84.315 ;
        RECT 173.695 78.215 173.955 78.535 ;
        RECT 173.755 72.415 173.895 78.215 ;
        RECT 174.155 77.875 174.415 78.195 ;
        RECT 174.215 74.875 174.355 77.875 ;
        RECT 174.675 75.475 174.815 83.995 ;
        RECT 175.595 83.295 175.735 85.015 ;
        RECT 175.535 82.975 175.795 83.295 ;
        RECT 176.055 82.615 176.195 85.355 ;
        RECT 175.995 82.295 176.255 82.615 ;
        RECT 176.975 80.915 177.115 89.095 ;
        RECT 178.355 89.075 178.495 90.455 ;
        RECT 178.295 88.755 178.555 89.075 ;
        RECT 177.645 87.200 179.185 87.570 ;
        RECT 179.675 85.015 179.935 85.335 ;
        RECT 177.645 81.760 179.185 82.130 ;
        RECT 179.735 81.255 179.875 85.015 ;
        RECT 179.675 80.935 179.935 81.255 ;
        RECT 176.915 80.595 177.175 80.915 ;
        RECT 176.975 78.875 177.115 80.595 ;
        RECT 180.195 79.805 180.335 95.815 ;
        RECT 180.945 95.360 182.485 95.730 ;
        RECT 180.945 89.920 182.485 90.290 ;
        RECT 180.945 84.480 182.485 84.850 ;
        RECT 182.955 81.255 183.095 99.635 ;
        RECT 183.355 96.575 183.615 96.895 ;
        RECT 183.415 94.515 183.555 96.575 ;
        RECT 183.875 95.195 184.015 99.635 ;
        RECT 183.815 94.875 184.075 95.195 ;
        RECT 183.355 94.195 183.615 94.515 ;
        RECT 183.355 91.475 183.615 91.795 ;
        RECT 183.415 88.735 183.555 91.475 ;
        RECT 183.875 89.270 184.015 94.875 ;
        RECT 183.805 88.900 184.085 89.270 ;
        RECT 183.355 88.415 183.615 88.735 ;
        RECT 183.415 86.355 183.555 88.415 ;
        RECT 183.355 86.035 183.615 86.355 ;
        RECT 183.415 84.315 183.555 86.035 ;
        RECT 183.815 85.355 184.075 85.675 ;
        RECT 183.875 84.315 184.015 85.355 ;
        RECT 183.355 83.995 183.615 84.315 ;
        RECT 183.815 83.995 184.075 84.315 ;
        RECT 183.875 81.595 184.015 83.995 ;
        RECT 183.815 81.275 184.075 81.595 ;
        RECT 182.895 80.935 183.155 81.255 ;
        RECT 179.735 79.665 180.335 79.805 ;
        RECT 176.915 78.555 177.175 78.875 ;
        RECT 176.975 78.195 177.115 78.555 ;
        RECT 179.735 78.535 179.875 79.665 ;
        RECT 180.595 79.575 180.855 79.895 ;
        RECT 179.675 78.390 179.935 78.535 ;
        RECT 176.915 77.875 177.175 78.195 ;
        RECT 179.665 78.020 179.945 78.390 ;
        RECT 180.655 77.855 180.795 79.575 ;
        RECT 180.945 79.040 182.485 79.410 ;
        RECT 180.595 77.535 180.855 77.855 ;
        RECT 181.975 77.535 182.235 77.855 ;
        RECT 175.995 76.855 176.255 77.175 ;
        RECT 180.135 76.855 180.395 77.175 ;
        RECT 175.535 75.835 175.795 76.155 ;
        RECT 174.615 75.155 174.875 75.475 ;
        RECT 174.215 74.735 174.815 74.875 ;
        RECT 174.155 74.135 174.415 74.455 ;
        RECT 174.215 73.435 174.355 74.135 ;
        RECT 174.155 73.115 174.415 73.435 ;
        RECT 173.695 72.095 173.955 72.415 ;
        RECT 173.235 70.395 173.495 70.715 ;
        RECT 174.675 70.375 174.815 74.735 ;
        RECT 175.075 74.135 175.335 74.455 ;
        RECT 175.135 73.630 175.275 74.135 ;
        RECT 175.065 73.260 175.345 73.630 ;
        RECT 175.595 72.415 175.735 75.835 ;
        RECT 176.055 73.095 176.195 76.855 ;
        RECT 177.645 76.320 179.185 76.690 ;
        RECT 175.995 72.775 176.255 73.095 ;
        RECT 180.195 72.835 180.335 76.855 ;
        RECT 180.595 74.475 180.855 74.795 ;
        RECT 180.655 73.435 180.795 74.475 ;
        RECT 182.035 74.455 182.175 77.535 ;
        RECT 182.955 76.235 183.095 80.935 ;
        RECT 183.355 80.595 183.615 80.915 ;
        RECT 183.415 77.175 183.555 80.595 ;
        RECT 183.355 76.855 183.615 77.175 ;
        RECT 182.955 76.095 184.015 76.235 ;
        RECT 184.335 76.155 184.475 105.075 ;
        RECT 184.795 100.635 184.935 109.225 ;
        RECT 187.095 107.775 187.235 109.225 ;
        RECT 187.035 107.455 187.295 107.775 ;
        RECT 187.035 106.775 187.295 107.095 ;
        RECT 185.195 105.075 185.455 105.395 ;
        RECT 184.735 100.315 184.995 100.635 ;
        RECT 185.255 100.035 185.395 105.075 ;
        RECT 187.095 104.375 187.235 106.775 ;
        RECT 189.395 106.075 189.535 109.225 ;
        RECT 189.335 105.755 189.595 106.075 ;
        RECT 189.795 105.755 190.055 106.075 ;
        RECT 186.575 104.055 186.835 104.375 ;
        RECT 187.035 104.055 187.295 104.375 ;
        RECT 189.335 104.055 189.595 104.375 ;
        RECT 186.635 103.435 186.775 104.055 ;
        RECT 186.635 103.295 187.235 103.435 ;
        RECT 186.115 102.355 186.375 102.675 ;
        RECT 186.175 100.295 186.315 102.355 ;
        RECT 184.795 99.895 185.395 100.035 ;
        RECT 186.115 99.975 186.375 100.295 ;
        RECT 184.795 80.915 184.935 99.895 ;
        RECT 186.575 99.635 186.835 99.955 ;
        RECT 186.635 99.275 186.775 99.635 ;
        RECT 186.575 98.955 186.835 99.275 ;
        RECT 185.195 96.235 185.455 96.555 ;
        RECT 185.655 96.235 185.915 96.555 ;
        RECT 185.255 94.515 185.395 96.235 ;
        RECT 185.715 95.195 185.855 96.235 ;
        RECT 186.115 95.895 186.375 96.215 ;
        RECT 185.655 94.875 185.915 95.195 ;
        RECT 186.175 94.855 186.315 95.895 ;
        RECT 186.115 94.535 186.375 94.855 ;
        RECT 185.195 94.195 185.455 94.515 ;
        RECT 185.255 91.195 185.395 94.195 ;
        RECT 185.255 91.055 185.855 91.195 ;
        RECT 185.195 90.455 185.455 90.775 ;
        RECT 185.255 83.635 185.395 90.455 ;
        RECT 185.715 83.635 185.855 91.055 ;
        RECT 186.175 87.035 186.315 94.535 ;
        RECT 186.635 89.755 186.775 98.955 ;
        RECT 187.095 97.315 187.235 103.295 ;
        RECT 187.495 101.675 187.755 101.995 ;
        RECT 187.555 97.915 187.695 101.675 ;
        RECT 188.875 101.335 189.135 101.655 ;
        RECT 187.955 98.615 188.215 98.935 ;
        RECT 187.495 97.595 187.755 97.915 ;
        RECT 187.095 97.235 187.695 97.315 ;
        RECT 187.095 97.175 187.755 97.235 ;
        RECT 187.495 96.915 187.755 97.175 ;
        RECT 187.025 96.380 187.305 96.750 ;
        RECT 186.575 89.435 186.835 89.755 ;
        RECT 186.115 86.715 186.375 87.035 ;
        RECT 186.175 85.335 186.315 86.715 ;
        RECT 186.115 85.015 186.375 85.335 ;
        RECT 185.195 83.315 185.455 83.635 ;
        RECT 185.655 83.315 185.915 83.635 ;
        RECT 184.735 80.595 184.995 80.915 ;
        RECT 184.735 79.915 184.995 80.235 ;
        RECT 182.495 74.735 183.555 74.875 ;
        RECT 182.495 74.455 182.635 74.735 ;
        RECT 181.975 74.135 182.235 74.455 ;
        RECT 182.435 74.135 182.695 74.455 ;
        RECT 180.945 73.600 182.485 73.970 ;
        RECT 180.595 73.115 180.855 73.435 ;
        RECT 182.885 73.260 183.165 73.630 ;
        RECT 177.375 72.435 177.635 72.755 ;
        RECT 179.215 72.435 179.475 72.755 ;
        RECT 180.195 72.695 180.795 72.835 ;
        RECT 175.535 72.095 175.795 72.415 ;
        RECT 177.435 72.155 177.575 72.435 ;
        RECT 176.975 72.015 177.575 72.155 ;
        RECT 175.995 71.415 176.255 71.735 ;
        RECT 174.155 70.055 174.415 70.375 ;
        RECT 174.615 70.055 174.875 70.375 ;
        RECT 174.215 67.655 174.355 70.055 ;
        RECT 176.055 69.695 176.195 71.415 ;
        RECT 175.995 69.550 176.255 69.695 ;
        RECT 175.985 69.180 176.265 69.550 ;
        RECT 175.535 68.695 175.795 69.015 ;
        RECT 172.305 67.140 172.585 67.510 ;
        RECT 172.775 67.335 173.035 67.655 ;
        RECT 174.155 67.335 174.415 67.655 ;
        RECT 169.555 65.185 169.815 65.275 ;
        RECT 169.155 65.045 169.815 65.185 ;
        RECT 146.290 58.035 148.395 63.305 ;
        RECT 169.155 62.555 169.295 65.045 ;
        RECT 169.555 64.955 169.815 65.045 ;
        RECT 175.595 64.935 175.735 68.695 ;
        RECT 175.535 64.615 175.795 64.935 ;
        RECT 173.235 63.595 173.495 63.915 ;
        RECT 169.095 62.235 169.355 62.555 ;
        RECT 173.295 62.215 173.435 63.595 ;
        RECT 176.055 62.555 176.195 69.180 ;
        RECT 176.975 67.315 177.115 72.015 ;
        RECT 179.275 71.735 179.415 72.435 ;
        RECT 180.655 72.415 180.795 72.695 ;
        RECT 180.595 72.095 180.855 72.415 ;
        RECT 179.675 71.755 179.935 72.075 ;
        RECT 179.215 71.415 179.475 71.735 ;
        RECT 177.645 70.880 179.185 71.250 ;
        RECT 179.735 70.910 179.875 71.755 ;
        RECT 179.665 70.540 179.945 70.910 ;
        RECT 177.375 70.055 177.635 70.375 ;
        RECT 177.435 69.015 177.575 70.055 ;
        RECT 179.675 69.715 179.935 70.035 ;
        RECT 177.375 68.695 177.635 69.015 ;
        RECT 176.915 66.995 177.175 67.315 ;
        RECT 176.975 64.595 177.115 66.995 ;
        RECT 177.645 65.440 179.185 65.810 ;
        RECT 179.735 64.595 179.875 69.715 ;
        RECT 182.955 69.015 183.095 73.260 ;
        RECT 182.895 68.695 183.155 69.015 ;
        RECT 180.945 68.160 182.485 68.530 ;
        RECT 181.055 67.335 181.315 67.655 ;
        RECT 180.595 65.975 180.855 66.295 ;
        RECT 180.655 65.275 180.795 65.975 ;
        RECT 180.595 64.955 180.855 65.275 ;
        RECT 176.915 64.275 177.175 64.595 ;
        RECT 179.675 64.275 179.935 64.595 ;
        RECT 176.455 63.255 176.715 63.575 ;
        RECT 175.995 62.235 176.255 62.555 ;
        RECT 173.235 61.895 173.495 62.215 ;
        RECT 176.515 61.535 176.655 63.255 ;
        RECT 176.975 62.215 177.115 64.275 ;
        RECT 179.665 63.740 179.945 64.110 ;
        RECT 180.135 63.935 180.395 64.255 ;
        RECT 181.115 63.995 181.255 67.335 ;
        RECT 176.915 61.895 177.175 62.215 ;
        RECT 175.075 61.275 175.335 61.535 ;
        RECT 175.075 61.215 176.195 61.275 ;
        RECT 176.455 61.215 176.715 61.535 ;
        RECT 175.135 61.135 176.195 61.215 ;
        RECT 176.055 60.855 176.195 61.135 ;
        RECT 164.035 60.710 164.295 60.855 ;
        RECT 164.025 60.340 164.305 60.710 ;
        RECT 175.995 60.535 176.255 60.855 ;
        RECT 176.055 59.495 176.195 60.535 ;
        RECT 177.645 60.000 179.185 60.370 ;
        RECT 175.995 59.175 176.255 59.495 ;
        RECT 172.315 58.835 172.575 59.155 ;
        RECT 167.715 57.815 167.975 58.135 ;
        RECT 146.290 53.355 148.395 57.455 ;
        RECT 167.775 56.775 167.915 57.815 ;
        RECT 167.715 56.455 167.975 56.775 ;
        RECT 166.335 55.775 166.595 56.095 ;
        RECT 165.875 53.115 166.135 53.375 ;
        RECT 166.395 53.115 166.535 55.775 ;
        RECT 165.875 53.055 166.535 53.115 ;
        RECT 165.935 52.975 166.535 53.055 ;
        RECT 146.290 48.675 148.395 52.775 ;
        RECT 166.395 50.655 166.535 52.975 ;
        RECT 172.375 51.675 172.515 58.835 ;
        RECT 177.375 58.495 177.635 58.815 ;
        RECT 176.915 56.795 177.175 57.115 ;
        RECT 174.155 56.455 174.415 56.775 ;
        RECT 174.215 53.035 174.355 56.455 ;
        RECT 175.075 56.115 175.335 56.435 ;
        RECT 174.155 52.715 174.415 53.035 ;
        RECT 172.315 51.355 172.575 51.675 ;
        RECT 166.335 50.335 166.595 50.655 ;
        RECT 170.935 50.335 171.195 50.655 ;
        RECT 146.290 43.995 148.395 48.095 ;
        RECT 166.395 45.215 166.535 50.335 ;
        RECT 170.995 48.955 171.135 50.335 ;
        RECT 170.935 48.635 171.195 48.955 ;
        RECT 172.375 48.275 172.515 51.355 ;
        RECT 174.215 51.335 174.355 52.715 ;
        RECT 174.155 51.015 174.415 51.335 ;
        RECT 172.775 49.655 173.035 49.975 ;
        RECT 172.315 47.955 172.575 48.275 ;
        RECT 172.835 47.255 172.975 49.655 ;
        RECT 175.135 47.935 175.275 56.115 ;
        RECT 175.535 55.095 175.795 55.415 ;
        RECT 175.595 54.055 175.735 55.095 ;
        RECT 176.975 54.055 177.115 56.795 ;
        RECT 177.435 55.755 177.575 58.495 ;
        RECT 177.835 57.815 178.095 58.135 ;
        RECT 177.895 56.775 178.035 57.815 ;
        RECT 179.735 57.115 179.875 63.740 ;
        RECT 180.195 59.835 180.335 63.935 ;
        RECT 180.655 63.915 181.255 63.995 ;
        RECT 180.655 63.855 181.315 63.915 ;
        RECT 180.655 60.855 180.795 63.855 ;
        RECT 181.055 63.595 181.315 63.855 ;
        RECT 180.945 62.720 182.485 63.090 ;
        RECT 181.055 61.215 181.315 61.535 ;
        RECT 180.595 60.535 180.855 60.855 ;
        RECT 180.135 59.515 180.395 59.835 ;
        RECT 180.595 59.515 180.855 59.835 ;
        RECT 180.655 59.065 180.795 59.515 ;
        RECT 181.115 59.155 181.255 61.215 ;
        RECT 180.195 58.925 180.795 59.065 ;
        RECT 179.675 56.795 179.935 57.115 ;
        RECT 177.835 56.455 178.095 56.775 ;
        RECT 179.675 55.775 179.935 56.095 ;
        RECT 177.375 55.435 177.635 55.755 ;
        RECT 177.645 54.560 179.185 54.930 ;
        RECT 175.535 53.735 175.795 54.055 ;
        RECT 176.915 53.735 177.175 54.055 ;
        RECT 179.735 51.675 179.875 55.775 ;
        RECT 179.675 51.355 179.935 51.675 ;
        RECT 180.195 51.335 180.335 58.925 ;
        RECT 181.055 58.835 181.315 59.155 ;
        RECT 182.435 58.670 182.695 58.815 ;
        RECT 180.595 58.155 180.855 58.475 ;
        RECT 182.425 58.300 182.705 58.670 ;
        RECT 180.655 56.435 180.795 58.155 ;
        RECT 180.945 57.280 182.485 57.650 ;
        RECT 182.955 57.115 183.095 68.695 ;
        RECT 183.415 64.255 183.555 74.735 ;
        RECT 183.875 69.015 184.015 76.095 ;
        RECT 184.275 75.835 184.535 76.155 ;
        RECT 184.265 75.300 184.545 75.670 ;
        RECT 183.815 68.695 184.075 69.015 ;
        RECT 183.815 65.975 184.075 66.295 ;
        RECT 183.875 64.595 184.015 65.975 ;
        RECT 183.815 64.275 184.075 64.595 ;
        RECT 183.355 63.935 183.615 64.255 ;
        RECT 184.335 61.535 184.475 75.300 ;
        RECT 184.795 74.455 184.935 79.915 ;
        RECT 184.735 74.135 184.995 74.455 ;
        RECT 184.725 72.580 185.005 72.950 ;
        RECT 184.735 72.435 184.995 72.580 ;
        RECT 184.795 63.915 184.935 72.435 ;
        RECT 185.255 67.655 185.395 83.315 ;
        RECT 187.095 83.295 187.235 96.380 ;
        RECT 187.495 95.895 187.755 96.215 ;
        RECT 187.555 93.495 187.695 95.895 ;
        RECT 187.495 93.175 187.755 93.495 ;
        RECT 188.015 89.415 188.155 98.615 ;
        RECT 187.955 89.095 188.215 89.415 ;
        RECT 188.015 86.695 188.155 89.095 ;
        RECT 187.955 86.375 188.215 86.695 ;
        RECT 187.955 85.695 188.215 86.015 ;
        RECT 187.035 82.975 187.295 83.295 ;
        RECT 187.495 82.975 187.755 83.295 ;
        RECT 186.115 81.275 186.375 81.595 ;
        RECT 185.655 79.575 185.915 79.895 ;
        RECT 185.715 77.710 185.855 79.575 ;
        RECT 185.645 77.340 185.925 77.710 ;
        RECT 185.655 77.195 185.915 77.340 ;
        RECT 185.655 75.495 185.915 75.815 ;
        RECT 186.175 75.670 186.315 81.275 ;
        RECT 186.575 77.535 186.835 77.855 ;
        RECT 185.715 72.415 185.855 75.495 ;
        RECT 186.105 75.300 186.385 75.670 ;
        RECT 186.115 75.045 186.375 75.135 ;
        RECT 186.635 75.045 186.775 77.535 ;
        RECT 187.035 76.855 187.295 77.175 ;
        RECT 187.095 76.155 187.235 76.855 ;
        RECT 187.035 75.835 187.295 76.155 ;
        RECT 186.115 74.905 186.775 75.045 ;
        RECT 186.115 74.815 186.375 74.905 ;
        RECT 186.575 73.395 186.835 73.435 ;
        RECT 187.095 73.395 187.235 75.835 ;
        RECT 186.575 73.255 187.235 73.395 ;
        RECT 186.575 73.115 186.835 73.255 ;
        RECT 185.655 72.095 185.915 72.415 ;
        RECT 185.655 69.375 185.915 69.695 ;
        RECT 187.035 69.375 187.295 69.695 ;
        RECT 185.195 67.335 185.455 67.655 ;
        RECT 185.255 65.275 185.395 67.335 ;
        RECT 185.195 64.955 185.455 65.275 ;
        RECT 185.715 64.595 185.855 69.375 ;
        RECT 186.115 68.695 186.375 69.015 ;
        RECT 186.175 66.295 186.315 68.695 ;
        RECT 186.115 65.975 186.375 66.295 ;
        RECT 185.655 64.275 185.915 64.595 ;
        RECT 184.735 63.595 184.995 63.915 ;
        RECT 184.795 62.555 184.935 63.595 ;
        RECT 184.735 62.235 184.995 62.555 ;
        RECT 184.275 61.215 184.535 61.535 ;
        RECT 184.735 60.535 184.995 60.855 ;
        RECT 183.815 58.835 184.075 59.155 ;
        RECT 183.355 57.815 183.615 58.135 ;
        RECT 182.895 56.795 183.155 57.115 ;
        RECT 181.515 56.630 181.775 56.775 ;
        RECT 180.595 56.115 180.855 56.435 ;
        RECT 181.505 56.260 181.785 56.630 ;
        RECT 183.415 56.345 183.555 57.815 ;
        RECT 182.955 56.205 183.555 56.345 ;
        RECT 182.435 56.005 182.695 56.095 ;
        RECT 182.955 56.005 183.095 56.205 ;
        RECT 182.435 55.865 183.095 56.005 ;
        RECT 182.435 55.775 182.695 55.865 ;
        RECT 183.345 55.580 183.625 55.950 ;
        RECT 183.875 55.755 184.015 58.835 ;
        RECT 184.795 57.310 184.935 60.535 ;
        RECT 185.715 59.835 185.855 64.275 ;
        RECT 186.175 63.575 186.315 65.975 ;
        RECT 187.095 64.255 187.235 69.375 ;
        RECT 187.035 64.110 187.295 64.255 ;
        RECT 187.025 63.740 187.305 64.110 ;
        RECT 186.115 63.255 186.375 63.575 ;
        RECT 187.035 63.255 187.295 63.575 ;
        RECT 186.175 61.535 186.315 63.255 ;
        RECT 186.575 61.555 186.835 61.875 ;
        RECT 186.115 61.215 186.375 61.535 ;
        RECT 186.115 60.535 186.375 60.855 ;
        RECT 185.655 59.515 185.915 59.835 ;
        RECT 186.175 58.815 186.315 60.535 ;
        RECT 186.635 58.815 186.775 61.555 ;
        RECT 187.095 61.195 187.235 63.255 ;
        RECT 187.555 61.875 187.695 82.975 ;
        RECT 188.015 80.915 188.155 85.695 ;
        RECT 188.415 82.635 188.675 82.955 ;
        RECT 187.955 80.595 188.215 80.915 ;
        RECT 188.475 80.315 188.615 82.635 ;
        RECT 188.015 80.175 188.615 80.315 ;
        RECT 188.015 62.215 188.155 80.175 ;
        RECT 188.415 77.875 188.675 78.195 ;
        RECT 188.475 75.475 188.615 77.875 ;
        RECT 188.935 77.855 189.075 101.335 ;
        RECT 189.395 100.295 189.535 104.055 ;
        RECT 189.335 99.975 189.595 100.295 ;
        RECT 189.855 98.935 189.995 105.755 ;
        RECT 191.695 105.735 191.835 109.225 ;
        RECT 191.635 105.415 191.895 105.735 ;
        RECT 193.475 105.075 193.735 105.395 ;
        RECT 192.555 104.735 192.815 105.055 ;
        RECT 191.175 104.055 191.435 104.375 ;
        RECT 189.795 98.615 190.055 98.935 ;
        RECT 191.235 95.955 191.375 104.055 ;
        RECT 192.615 103.015 192.755 104.735 ;
        RECT 193.535 104.375 193.675 105.075 ;
        RECT 193.995 104.715 194.135 109.225 ;
        RECT 196.295 107.095 196.435 109.225 ;
        RECT 197.615 107.115 197.875 107.435 ;
        RECT 196.235 106.775 196.495 107.095 ;
        RECT 194.855 105.075 195.115 105.395 ;
        RECT 195.775 105.075 196.035 105.395 ;
        RECT 193.935 104.395 194.195 104.715 ;
        RECT 193.475 104.055 193.735 104.375 ;
        RECT 192.555 102.695 192.815 103.015 ;
        RECT 192.615 97.235 192.755 102.695 ;
        RECT 193.015 99.295 193.275 99.615 ;
        RECT 192.555 96.915 192.815 97.235 ;
        RECT 191.235 95.815 192.295 95.955 ;
        RECT 191.175 93.515 191.435 93.835 ;
        RECT 189.795 88.755 190.055 89.075 ;
        RECT 189.855 86.015 189.995 88.755 ;
        RECT 190.715 88.415 190.975 88.735 ;
        RECT 189.795 85.695 190.055 86.015 ;
        RECT 190.255 85.695 190.515 86.015 ;
        RECT 189.855 83.635 189.995 85.695 ;
        RECT 189.795 83.315 190.055 83.635 ;
        RECT 188.875 77.535 189.135 77.855 ;
        RECT 188.415 75.155 188.675 75.475 ;
        RECT 188.475 70.035 188.615 75.155 ;
        RECT 189.335 74.475 189.595 74.795 ;
        RECT 188.415 69.715 188.675 70.035 ;
        RECT 189.395 67.655 189.535 74.475 ;
        RECT 189.335 67.335 189.595 67.655 ;
        RECT 189.335 66.655 189.595 66.975 ;
        RECT 187.955 61.895 188.215 62.215 ;
        RECT 187.495 61.555 187.755 61.875 ;
        RECT 188.415 61.555 188.675 61.875 ;
        RECT 187.035 60.875 187.295 61.195 ;
        RECT 185.655 58.495 185.915 58.815 ;
        RECT 186.115 58.495 186.375 58.815 ;
        RECT 186.575 58.495 186.835 58.815 ;
        RECT 185.195 58.155 185.455 58.475 ;
        RECT 184.725 56.940 185.005 57.310 ;
        RECT 185.255 57.115 185.395 58.155 ;
        RECT 185.195 56.795 185.455 57.115 ;
        RECT 185.715 56.095 185.855 58.495 ;
        RECT 186.635 57.115 186.775 58.495 ;
        RECT 187.555 57.195 187.695 61.555 ;
        RECT 186.575 56.795 186.835 57.115 ;
        RECT 187.555 57.055 188.155 57.195 ;
        RECT 184.735 55.775 184.995 56.095 ;
        RECT 185.655 55.775 185.915 56.095 ;
        RECT 183.355 55.435 183.615 55.580 ;
        RECT 183.815 55.435 184.075 55.755 ;
        RECT 182.895 53.055 183.155 53.375 ;
        RECT 180.945 51.840 182.485 52.210 ;
        RECT 176.455 51.015 176.715 51.335 ;
        RECT 180.135 51.015 180.395 51.335 ;
        RECT 175.995 50.675 176.255 50.995 ;
        RECT 176.055 50.510 176.195 50.675 ;
        RECT 175.985 50.140 176.265 50.510 ;
        RECT 175.075 47.615 175.335 47.935 ;
        RECT 170.935 46.935 171.195 47.255 ;
        RECT 172.775 46.935 173.035 47.255 ;
        RECT 166.335 45.125 166.595 45.215 ;
        RECT 165.935 44.985 166.595 45.125 ;
        RECT 143.435 41.655 145.540 42.245 ;
        RECT 143.835 41.605 145.135 41.655 ;
        RECT 7.065 36.430 8.665 39.630 ;
        RECT 10.170 37.965 74.550 38.965 ;
        RECT 79.810 38.185 127.975 39.285 ;
        RECT 10.170 35.440 74.550 36.940 ;
        RECT 79.810 36.685 127.975 37.785 ;
        RECT 79.810 35.185 127.975 36.285 ;
        RECT 136.295 35.805 138.400 39.905 ;
        RECT 146.290 38.145 148.395 43.415 ;
        RECT 165.935 42.495 166.075 44.985 ;
        RECT 166.335 44.895 166.595 44.985 ;
        RECT 165.875 42.175 166.135 42.495 ;
        RECT 10.170 33.440 74.550 34.940 ;
        RECT 79.810 33.685 127.975 34.785 ;
        RECT 10.170 31.440 74.550 32.940 ;
        RECT 79.810 32.185 127.975 33.285 ;
        RECT 79.810 30.685 127.975 31.785 ;
        RECT 136.295 31.125 138.400 35.225 ;
        RECT 146.290 33.465 148.395 37.565 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 165.935 31.955 166.075 42.175 ;
        RECT 167.255 41.835 167.515 42.155 ;
        RECT 167.315 40.795 167.455 41.835 ;
        RECT 167.255 40.475 167.515 40.795 ;
        RECT 165.875 31.635 166.135 31.955 ;
        RECT 10.170 28.035 74.550 30.415 ;
        RECT 79.810 28.165 127.975 30.285 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 170.995 29.235 171.135 46.935 ;
        RECT 176.515 46.235 176.655 51.015 ;
        RECT 182.955 50.995 183.095 53.055 ;
        RECT 183.355 52.715 183.615 53.035 ;
        RECT 183.415 50.995 183.555 52.715 ;
        RECT 183.875 52.695 184.015 55.435 ;
        RECT 184.795 54.055 184.935 55.775 ;
        RECT 186.635 55.755 186.775 56.795 ;
        RECT 187.035 56.115 187.295 56.435 ;
        RECT 186.575 55.435 186.835 55.755 ;
        RECT 184.735 53.735 184.995 54.055 ;
        RECT 183.815 52.375 184.075 52.695 ;
        RECT 184.795 51.245 184.935 53.735 ;
        RECT 187.095 53.375 187.235 56.115 ;
        RECT 188.015 54.475 188.155 57.055 ;
        RECT 188.475 55.415 188.615 61.555 ;
        RECT 188.875 60.875 189.135 61.195 ;
        RECT 188.415 55.095 188.675 55.415 ;
        RECT 188.015 54.335 188.615 54.475 ;
        RECT 188.935 54.395 189.075 60.875 ;
        RECT 189.395 59.495 189.535 66.655 ;
        RECT 189.855 62.555 189.995 83.315 ;
        RECT 190.315 82.955 190.455 85.695 ;
        RECT 190.255 82.635 190.515 82.955 ;
        RECT 190.315 81.595 190.455 82.635 ;
        RECT 190.775 82.615 190.915 88.415 ;
        RECT 190.715 82.295 190.975 82.615 ;
        RECT 190.255 81.275 190.515 81.595 ;
        RECT 190.775 80.575 190.915 82.295 ;
        RECT 190.715 80.255 190.975 80.575 ;
        RECT 190.255 78.215 190.515 78.535 ;
        RECT 190.315 72.755 190.455 78.215 ;
        RECT 190.715 75.155 190.975 75.475 ;
        RECT 190.255 72.435 190.515 72.755 ;
        RECT 190.315 69.355 190.455 72.435 ;
        RECT 190.775 70.715 190.915 75.155 ;
        RECT 191.235 75.135 191.375 93.515 ;
        RECT 191.635 80.595 191.895 80.915 ;
        RECT 191.175 74.815 191.435 75.135 ;
        RECT 191.175 74.135 191.435 74.455 ;
        RECT 191.235 71.735 191.375 74.135 ;
        RECT 191.175 71.415 191.435 71.735 ;
        RECT 190.715 70.395 190.975 70.715 ;
        RECT 190.255 69.035 190.515 69.355 ;
        RECT 189.795 62.235 190.055 62.555 ;
        RECT 189.795 61.215 190.055 61.535 ;
        RECT 189.335 59.175 189.595 59.495 ;
        RECT 189.855 59.155 189.995 61.215 ;
        RECT 189.795 58.835 190.055 59.155 ;
        RECT 189.335 56.455 189.595 56.775 ;
        RECT 187.955 53.395 188.215 53.715 ;
        RECT 187.035 53.055 187.295 53.375 ;
        RECT 187.495 52.945 187.755 53.035 ;
        RECT 188.015 52.945 188.155 53.395 ;
        RECT 187.495 52.805 188.155 52.945 ;
        RECT 187.495 52.715 187.755 52.805 ;
        RECT 185.195 52.550 185.455 52.695 ;
        RECT 185.185 52.180 185.465 52.550 ;
        RECT 185.195 51.245 185.455 51.335 ;
        RECT 184.795 51.105 185.455 51.245 ;
        RECT 185.195 51.015 185.455 51.105 ;
        RECT 182.895 50.675 183.155 50.995 ;
        RECT 183.355 50.675 183.615 50.995 ;
        RECT 177.645 49.120 179.185 49.490 ;
        RECT 180.135 47.615 180.395 47.935 ;
        RECT 176.915 46.935 177.175 47.255 ;
        RECT 179.675 46.935 179.935 47.255 ;
        RECT 176.455 45.915 176.715 46.235 ;
        RECT 175.535 44.215 175.795 44.535 ;
        RECT 175.595 42.835 175.735 44.215 ;
        RECT 175.535 42.515 175.795 42.835 ;
        RECT 172.315 41.495 172.575 41.815 ;
        RECT 172.375 40.455 172.515 41.495 ;
        RECT 172.315 40.135 172.575 40.455 ;
        RECT 171.395 36.735 171.655 37.055 ;
        RECT 171.455 35.355 171.595 36.735 ;
        RECT 172.375 35.355 172.515 40.135 ;
        RECT 175.075 39.455 175.335 39.775 ;
        RECT 175.135 38.075 175.275 39.455 ;
        RECT 175.075 37.755 175.335 38.075 ;
        RECT 175.075 36.735 175.335 37.055 ;
        RECT 171.395 35.035 171.655 35.355 ;
        RECT 172.315 35.035 172.575 35.355 ;
        RECT 175.135 32.295 175.275 36.735 ;
        RECT 175.595 34.675 175.735 42.515 ;
        RECT 176.975 42.155 177.115 46.935 ;
        RECT 177.645 43.680 179.185 44.050 ;
        RECT 176.915 41.835 177.175 42.155 ;
        RECT 176.915 39.455 177.175 39.775 ;
        RECT 176.975 36.715 177.115 39.455 ;
        RECT 179.735 39.095 179.875 46.935 ;
        RECT 180.195 43.515 180.335 47.615 ;
        RECT 182.955 47.595 183.095 50.675 ;
        RECT 182.895 47.275 183.155 47.595 ;
        RECT 180.945 46.400 182.485 46.770 ;
        RECT 182.955 43.515 183.095 47.275 ;
        RECT 183.415 46.235 183.555 50.675 ;
        RECT 187.035 50.335 187.295 50.655 ;
        RECT 184.735 47.955 184.995 48.275 ;
        RECT 183.815 46.935 184.075 47.255 ;
        RECT 183.355 45.915 183.615 46.235 ;
        RECT 183.875 45.215 184.015 46.935 ;
        RECT 184.275 45.235 184.535 45.555 ;
        RECT 183.815 44.895 184.075 45.215 ;
        RECT 180.135 43.195 180.395 43.515 ;
        RECT 182.895 43.195 183.155 43.515 ;
        RECT 180.945 40.960 182.485 41.330 ;
        RECT 183.875 40.795 184.015 44.895 ;
        RECT 184.335 42.155 184.475 45.235 ;
        RECT 184.795 45.215 184.935 47.955 ;
        RECT 184.735 44.895 184.995 45.215 ;
        RECT 184.275 41.835 184.535 42.155 ;
        RECT 186.115 41.835 186.375 42.155 ;
        RECT 183.815 40.475 184.075 40.795 ;
        RECT 180.135 39.455 180.395 39.775 ;
        RECT 179.675 38.775 179.935 39.095 ;
        RECT 177.645 38.240 179.185 38.610 ;
        RECT 178.755 37.075 179.015 37.395 ;
        RECT 176.915 36.395 177.175 36.715 ;
        RECT 176.975 35.355 177.115 36.395 ;
        RECT 176.915 35.035 177.175 35.355 ;
        RECT 178.815 34.675 178.955 37.075 ;
        RECT 179.735 36.715 179.875 38.775 ;
        RECT 180.195 37.395 180.335 39.455 ;
        RECT 180.135 37.075 180.395 37.395 ;
        RECT 182.895 36.735 183.155 37.055 ;
        RECT 179.675 36.395 179.935 36.715 ;
        RECT 180.945 35.520 182.485 35.890 ;
        RECT 180.135 34.695 180.395 35.015 ;
        RECT 175.535 34.355 175.795 34.675 ;
        RECT 176.915 34.355 177.175 34.675 ;
        RECT 178.755 34.355 179.015 34.675 ;
        RECT 175.075 31.975 175.335 32.295 ;
        RECT 175.135 29.235 175.275 31.975 ;
        RECT 176.975 31.955 177.115 34.355 ;
        RECT 179.675 34.015 179.935 34.335 ;
        RECT 177.645 32.800 179.185 33.170 ;
        RECT 179.735 32.295 179.875 34.015 ;
        RECT 179.675 31.975 179.935 32.295 ;
        RECT 176.915 31.635 177.175 31.955 ;
        RECT 176.975 29.915 177.115 31.635 ;
        RECT 179.675 31.295 179.935 31.615 ;
        RECT 176.915 29.595 177.175 29.915 ;
        RECT 170.935 28.915 171.195 29.235 ;
        RECT 175.075 28.915 175.335 29.235 ;
        RECT 164.035 28.070 164.295 28.215 ;
        RECT 10.170 25.510 74.550 27.010 ;
        RECT 79.810 26.665 127.975 27.765 ;
        RECT 164.025 27.700 164.305 28.070 ;
        RECT 177.645 27.360 179.185 27.730 ;
        RECT 179.735 27.195 179.875 31.295 ;
        RECT 180.195 28.895 180.335 34.695 ;
        RECT 182.955 32.635 183.095 36.735 ;
        RECT 183.355 33.335 183.615 33.655 ;
        RECT 182.895 32.315 183.155 32.635 ;
        RECT 180.945 30.080 182.485 30.450 ;
        RECT 180.135 28.575 180.395 28.895 ;
        RECT 179.675 26.875 179.935 27.195 ;
        RECT 180.195 26.515 180.335 28.575 ;
        RECT 183.415 26.515 183.555 33.335 ;
        RECT 184.335 30.935 184.475 41.835 ;
        RECT 186.175 40.795 186.315 41.835 ;
        RECT 186.115 40.475 186.375 40.795 ;
        RECT 185.655 40.135 185.915 40.455 ;
        RECT 185.715 35.355 185.855 40.135 ;
        RECT 187.095 40.115 187.235 50.335 ;
        RECT 188.475 44.535 188.615 54.335 ;
        RECT 188.875 54.075 189.135 54.395 ;
        RECT 189.395 52.695 189.535 56.455 ;
        RECT 189.855 55.415 189.995 58.835 ;
        RECT 189.795 55.095 190.055 55.415 ;
        RECT 189.795 54.075 190.055 54.395 ;
        RECT 189.335 52.375 189.595 52.695 ;
        RECT 189.335 51.015 189.595 51.335 ;
        RECT 189.395 45.555 189.535 51.015 ;
        RECT 189.855 50.315 189.995 54.075 ;
        RECT 190.315 50.995 190.455 69.035 ;
        RECT 191.235 66.635 191.375 71.415 ;
        RECT 191.175 66.545 191.435 66.635 ;
        RECT 190.775 66.405 191.435 66.545 ;
        RECT 190.775 59.155 190.915 66.405 ;
        RECT 191.175 66.315 191.435 66.405 ;
        RECT 191.695 59.745 191.835 80.595 ;
        RECT 192.155 77.175 192.295 95.815 ;
        RECT 192.615 94.175 192.755 96.915 ;
        RECT 193.075 94.855 193.215 99.295 ;
        RECT 193.475 98.615 193.735 98.935 ;
        RECT 193.535 96.750 193.675 98.615 ;
        RECT 193.465 96.380 193.745 96.750 ;
        RECT 193.015 94.535 193.275 94.855 ;
        RECT 193.535 94.515 193.675 96.380 ;
        RECT 193.935 96.125 194.195 96.215 ;
        RECT 194.915 96.125 195.055 105.075 ;
        RECT 195.835 104.795 195.975 105.075 ;
        RECT 195.375 104.655 195.975 104.795 ;
        RECT 195.375 101.655 195.515 104.655 ;
        RECT 196.235 102.015 196.495 102.335 ;
        RECT 195.315 101.335 195.575 101.655 ;
        RECT 195.375 96.215 195.515 101.335 ;
        RECT 196.295 100.295 196.435 102.015 ;
        RECT 197.675 101.995 197.815 107.115 ;
        RECT 198.595 106.075 198.735 109.225 ;
        RECT 198.535 105.755 198.795 106.075 ;
        RECT 198.995 105.075 199.255 105.395 ;
        RECT 199.055 102.335 199.195 105.075 ;
        RECT 200.375 104.735 200.635 105.055 ;
        RECT 200.435 102.335 200.575 104.735 ;
        RECT 200.895 104.715 201.035 109.225 ;
        RECT 200.835 104.395 201.095 104.715 ;
        RECT 203.195 103.355 203.335 109.225 ;
        RECT 204.975 107.455 205.235 107.775 ;
        RECT 204.515 105.075 204.775 105.395 ;
        RECT 203.135 103.035 203.395 103.355 ;
        RECT 198.995 102.015 199.255 102.335 ;
        RECT 200.375 102.015 200.635 102.335 ;
        RECT 197.615 101.675 197.875 101.995 ;
        RECT 197.155 101.335 197.415 101.655 ;
        RECT 196.235 99.975 196.495 100.295 ;
        RECT 195.775 97.595 196.035 97.915 ;
        RECT 195.835 96.895 195.975 97.595 ;
        RECT 197.215 96.895 197.355 101.335 ;
        RECT 200.435 100.635 200.575 102.015 ;
        RECT 204.575 100.715 204.715 105.075 ;
        RECT 205.035 104.375 205.175 107.455 ;
        RECT 205.495 105.055 205.635 109.225 ;
        RECT 207.795 106.075 207.935 109.225 ;
        RECT 208.655 107.115 208.915 107.435 ;
        RECT 207.735 105.755 207.995 106.075 ;
        RECT 208.715 105.735 208.855 107.115 ;
        RECT 208.655 105.415 208.915 105.735 ;
        RECT 207.735 105.075 207.995 105.395 ;
        RECT 205.435 104.735 205.695 105.055 ;
        RECT 204.975 104.055 205.235 104.375 ;
        RECT 205.895 104.055 206.155 104.375 ;
        RECT 205.955 101.995 206.095 104.055 ;
        RECT 207.795 103.355 207.935 105.075 ;
        RECT 207.735 103.035 207.995 103.355 ;
        RECT 205.895 101.675 206.155 101.995 ;
        RECT 207.735 101.675 207.995 101.995 ;
        RECT 200.375 100.315 200.635 100.635 ;
        RECT 204.575 100.575 205.175 100.715 ;
        RECT 198.075 99.975 198.335 100.295 ;
        RECT 198.135 97.235 198.275 99.975 ;
        RECT 198.075 96.915 198.335 97.235 ;
        RECT 195.775 96.575 196.035 96.895 ;
        RECT 193.935 95.985 195.055 96.125 ;
        RECT 193.935 95.895 194.195 95.985 ;
        RECT 195.315 95.895 195.575 96.215 ;
        RECT 193.995 95.195 194.135 95.895 ;
        RECT 193.935 94.875 194.195 95.195 ;
        RECT 193.475 94.195 193.735 94.515 ;
        RECT 192.555 93.855 192.815 94.175 ;
        RECT 193.995 94.030 194.135 94.875 ;
        RECT 195.375 94.710 195.515 95.895 ;
        RECT 195.305 94.340 195.585 94.710 ;
        RECT 193.925 93.660 194.205 94.030 ;
        RECT 194.395 91.135 194.655 91.455 ;
        RECT 195.315 91.135 195.575 91.455 ;
        RECT 193.015 90.795 193.275 91.115 ;
        RECT 193.075 89.075 193.215 90.795 ;
        RECT 193.015 88.755 193.275 89.075 ;
        RECT 194.455 86.015 194.595 91.135 ;
        RECT 194.855 88.755 195.115 89.075 ;
        RECT 194.395 85.695 194.655 86.015 ;
        RECT 193.015 83.655 193.275 83.975 ;
        RECT 192.555 77.535 192.815 77.855 ;
        RECT 192.095 76.855 192.355 77.175 ;
        RECT 192.615 74.795 192.755 77.535 ;
        RECT 192.555 74.475 192.815 74.795 ;
        RECT 192.615 73.095 192.755 74.475 ;
        RECT 192.555 72.775 192.815 73.095 ;
        RECT 192.555 72.095 192.815 72.415 ;
        RECT 192.615 70.035 192.755 72.095 ;
        RECT 192.555 69.715 192.815 70.035 ;
        RECT 192.095 68.925 192.355 69.015 ;
        RECT 192.095 68.785 192.755 68.925 ;
        RECT 192.095 68.695 192.355 68.785 ;
        RECT 192.615 68.190 192.755 68.785 ;
        RECT 192.545 67.820 192.825 68.190 ;
        RECT 192.615 67.655 192.755 67.820 ;
        RECT 192.555 67.335 192.815 67.655 ;
        RECT 192.545 64.420 192.825 64.790 ;
        RECT 192.615 64.255 192.755 64.420 ;
        RECT 192.555 63.935 192.815 64.255 ;
        RECT 192.095 61.215 192.355 61.535 ;
        RECT 191.235 59.605 191.835 59.745 ;
        RECT 190.715 58.835 190.975 59.155 ;
        RECT 191.235 58.135 191.375 59.605 ;
        RECT 192.155 58.815 192.295 61.215 ;
        RECT 193.075 59.835 193.215 83.655 ;
        RECT 194.915 81.595 195.055 88.755 ;
        RECT 195.375 88.055 195.515 91.135 ;
        RECT 195.835 89.415 195.975 96.575 ;
        RECT 196.685 96.380 196.965 96.750 ;
        RECT 197.155 96.575 197.415 96.895 ;
        RECT 196.755 94.175 196.895 96.380 ;
        RECT 198.535 95.895 198.795 96.215 ;
        RECT 196.695 93.855 196.955 94.175 ;
        RECT 198.595 91.455 198.735 95.895 ;
        RECT 200.435 94.855 200.575 100.315 ;
        RECT 204.515 98.615 204.775 98.935 ;
        RECT 203.585 97.060 203.865 97.430 ;
        RECT 203.655 96.895 203.795 97.060 ;
        RECT 203.595 96.575 203.855 96.895 ;
        RECT 204.575 96.555 204.715 98.615 ;
        RECT 204.515 96.235 204.775 96.555 ;
        RECT 200.375 94.535 200.635 94.855 ;
        RECT 204.515 93.515 204.775 93.835 ;
        RECT 203.135 92.155 203.395 92.475 ;
        RECT 203.595 92.155 203.855 92.475 ;
        RECT 198.535 91.135 198.795 91.455 ;
        RECT 200.825 90.940 201.105 91.310 ;
        RECT 198.535 90.455 198.795 90.775 ;
        RECT 195.775 89.095 196.035 89.415 ;
        RECT 195.315 87.735 195.575 88.055 ;
        RECT 198.075 86.035 198.335 86.355 ;
        RECT 195.775 85.695 196.035 86.015 ;
        RECT 195.835 85.335 195.975 85.695 ;
        RECT 198.135 85.335 198.275 86.035 ;
        RECT 195.775 85.015 196.035 85.335 ;
        RECT 198.075 85.015 198.335 85.335 ;
        RECT 194.855 81.275 195.115 81.595 ;
        RECT 194.395 69.715 194.655 70.035 ;
        RECT 193.935 69.435 194.195 69.695 ;
        RECT 193.535 69.375 194.195 69.435 ;
        RECT 193.535 69.295 194.135 69.375 ;
        RECT 193.535 65.275 193.675 69.295 ;
        RECT 194.455 67.315 194.595 69.715 ;
        RECT 195.315 67.675 195.575 67.995 ;
        RECT 194.395 66.995 194.655 67.315 ;
        RECT 193.475 64.955 193.735 65.275 ;
        RECT 193.535 63.915 193.675 64.955 ;
        RECT 193.935 64.110 194.195 64.255 ;
        RECT 193.475 63.595 193.735 63.915 ;
        RECT 193.925 63.740 194.205 64.110 ;
        RECT 193.535 61.390 193.675 63.595 ;
        RECT 195.375 62.555 195.515 67.675 ;
        RECT 195.835 64.935 195.975 85.015 ;
        RECT 197.605 82.780 197.885 83.150 ;
        RECT 197.675 78.195 197.815 82.780 ;
        RECT 197.615 77.875 197.875 78.195 ;
        RECT 198.075 77.535 198.335 77.855 ;
        RECT 196.235 69.375 196.495 69.695 ;
        RECT 197.155 69.375 197.415 69.695 ;
        RECT 195.775 64.615 196.035 64.935 ;
        RECT 196.295 64.790 196.435 69.375 ;
        RECT 196.695 67.335 196.955 67.655 ;
        RECT 196.755 64.935 196.895 67.335 ;
        RECT 196.225 64.420 196.505 64.790 ;
        RECT 196.695 64.615 196.955 64.935 ;
        RECT 195.775 63.935 196.035 64.255 ;
        RECT 195.835 63.575 195.975 63.935 ;
        RECT 196.235 63.595 196.495 63.915 ;
        RECT 195.775 63.255 196.035 63.575 ;
        RECT 195.315 62.235 195.575 62.555 ;
        RECT 193.465 61.020 193.745 61.390 ;
        RECT 193.015 59.515 193.275 59.835 ;
        RECT 192.095 58.725 192.355 58.815 ;
        RECT 191.695 58.585 192.355 58.725 ;
        RECT 191.175 57.815 191.435 58.135 ;
        RECT 191.695 56.095 191.835 58.585 ;
        RECT 192.095 58.495 192.355 58.585 ;
        RECT 193.015 58.495 193.275 58.815 ;
        RECT 192.095 56.115 192.355 56.435 ;
        RECT 191.635 55.775 191.895 56.095 ;
        RECT 191.695 53.375 191.835 55.775 ;
        RECT 192.155 53.375 192.295 56.115 ;
        RECT 193.075 55.755 193.215 58.495 ;
        RECT 195.835 57.115 195.975 63.255 ;
        RECT 196.295 61.195 196.435 63.595 ;
        RECT 196.755 63.575 196.895 64.615 ;
        RECT 197.215 64.110 197.355 69.375 ;
        RECT 197.615 67.225 197.875 67.315 ;
        RECT 198.135 67.225 198.275 77.535 ;
        RECT 197.615 67.085 198.275 67.225 ;
        RECT 197.615 66.995 197.875 67.085 ;
        RECT 197.145 63.740 197.425 64.110 ;
        RECT 197.615 63.935 197.875 64.255 ;
        RECT 196.695 63.255 196.955 63.575 ;
        RECT 196.235 60.875 196.495 61.195 ;
        RECT 196.295 58.815 196.435 60.875 ;
        RECT 196.695 60.535 196.955 60.855 ;
        RECT 196.235 58.495 196.495 58.815 ;
        RECT 195.775 56.795 196.035 57.115 ;
        RECT 193.015 55.435 193.275 55.755 ;
        RECT 193.475 55.435 193.735 55.755 ;
        RECT 194.385 55.580 194.665 55.950 ;
        RECT 191.635 53.055 191.895 53.375 ;
        RECT 192.095 53.055 192.355 53.375 ;
        RECT 191.695 52.550 191.835 53.055 ;
        RECT 191.625 52.180 191.905 52.550 ;
        RECT 190.255 50.675 190.515 50.995 ;
        RECT 189.795 49.995 190.055 50.315 ;
        RECT 190.315 48.955 190.455 50.675 ;
        RECT 190.255 48.635 190.515 48.955 ;
        RECT 189.335 45.235 189.595 45.555 ;
        RECT 188.415 44.215 188.675 44.535 ;
        RECT 189.395 42.835 189.535 45.235 ;
        RECT 189.335 42.515 189.595 42.835 ;
        RECT 187.035 39.795 187.295 40.115 ;
        RECT 187.095 38.075 187.235 39.795 ;
        RECT 187.495 39.455 187.755 39.775 ;
        RECT 187.035 37.755 187.295 38.075 ;
        RECT 187.035 37.075 187.295 37.395 ;
        RECT 185.655 35.035 185.915 35.355 ;
        RECT 187.095 35.015 187.235 37.075 ;
        RECT 187.555 35.355 187.695 39.455 ;
        RECT 187.495 35.035 187.755 35.355 ;
        RECT 187.035 34.695 187.295 35.015 ;
        RECT 186.575 30.955 186.835 31.275 ;
        RECT 187.955 30.955 188.215 31.275 ;
        RECT 184.275 30.615 184.535 30.935 ;
        RECT 186.115 30.615 186.375 30.935 ;
        RECT 184.335 29.915 184.475 30.615 ;
        RECT 184.275 29.595 184.535 29.915 ;
        RECT 186.175 29.575 186.315 30.615 ;
        RECT 186.635 29.915 186.775 30.955 ;
        RECT 186.575 29.595 186.835 29.915 ;
        RECT 186.115 29.255 186.375 29.575 ;
        RECT 188.015 27.195 188.155 30.955 ;
        RECT 189.395 29.235 189.535 42.515 ;
        RECT 190.255 41.495 190.515 41.815 ;
        RECT 190.315 40.795 190.455 41.495 ;
        RECT 191.695 40.795 191.835 52.180 ;
        RECT 192.155 51.675 192.295 53.055 ;
        RECT 192.095 51.355 192.355 51.675 ;
        RECT 192.555 41.835 192.815 42.155 ;
        RECT 190.255 40.475 190.515 40.795 ;
        RECT 191.635 40.475 191.895 40.795 ;
        RECT 192.615 37.395 192.755 41.835 ;
        RECT 193.075 41.815 193.215 55.435 ;
        RECT 193.535 51.335 193.675 55.435 ;
        RECT 194.455 55.415 194.595 55.580 ;
        RECT 193.935 55.095 194.195 55.415 ;
        RECT 194.395 55.095 194.655 55.415 ;
        RECT 193.995 53.035 194.135 55.095 ;
        RECT 196.295 54.055 196.435 58.495 ;
        RECT 196.755 56.775 196.895 60.535 ;
        RECT 197.675 59.835 197.815 63.935 ;
        RECT 198.135 63.915 198.275 67.085 ;
        RECT 198.075 63.595 198.335 63.915 ;
        RECT 198.595 61.875 198.735 90.455 ;
        RECT 199.455 87.735 199.715 88.055 ;
        RECT 198.995 85.015 199.255 85.335 ;
        RECT 199.055 61.875 199.195 85.015 ;
        RECT 199.515 80.575 199.655 87.735 ;
        RECT 200.895 86.015 201.035 90.940 ;
        RECT 203.195 89.415 203.335 92.155 ;
        RECT 203.135 89.095 203.395 89.415 ;
        RECT 203.195 86.015 203.335 89.095 ;
        RECT 203.655 89.075 203.795 92.155 ;
        RECT 204.575 89.075 204.715 93.515 ;
        RECT 203.595 88.755 203.855 89.075 ;
        RECT 204.515 88.755 204.775 89.075 ;
        RECT 200.835 85.695 201.095 86.015 ;
        RECT 203.135 85.695 203.395 86.015 ;
        RECT 202.215 85.355 202.475 85.675 ;
        RECT 202.275 83.295 202.415 85.355 ;
        RECT 202.215 83.205 202.475 83.295 ;
        RECT 202.215 83.065 202.875 83.205 ;
        RECT 202.215 82.975 202.475 83.065 ;
        RECT 199.915 81.275 200.175 81.595 ;
        RECT 199.455 80.255 199.715 80.575 ;
        RECT 199.515 78.195 199.655 80.255 ;
        RECT 199.975 78.195 200.115 81.275 ;
        RECT 202.215 80.255 202.475 80.575 ;
        RECT 199.455 77.875 199.715 78.195 ;
        RECT 199.915 77.875 200.175 78.195 ;
        RECT 199.515 67.995 199.655 77.875 ;
        RECT 199.975 75.725 200.115 77.875 ;
        RECT 201.755 76.855 202.015 77.175 ;
        RECT 200.375 75.725 200.635 75.815 ;
        RECT 199.975 75.585 200.635 75.725 ;
        RECT 200.375 75.495 200.635 75.585 ;
        RECT 200.835 74.475 201.095 74.795 ;
        RECT 200.895 73.095 201.035 74.475 ;
        RECT 200.835 72.775 201.095 73.095 ;
        RECT 201.295 72.095 201.555 72.415 ;
        RECT 201.355 70.715 201.495 72.095 ;
        RECT 201.295 70.395 201.555 70.715 ;
        RECT 199.455 67.675 199.715 67.995 ;
        RECT 199.915 66.995 200.175 67.315 ;
        RECT 200.375 66.995 200.635 67.315 ;
        RECT 199.975 66.830 200.115 66.995 ;
        RECT 199.905 66.460 200.185 66.830 ;
        RECT 199.455 65.975 199.715 66.295 ;
        RECT 199.515 61.875 199.655 65.975 ;
        RECT 200.435 65.275 200.575 66.995 ;
        RECT 200.375 64.955 200.635 65.275 ;
        RECT 201.295 63.255 201.555 63.575 ;
        RECT 198.535 61.555 198.795 61.875 ;
        RECT 198.995 61.555 199.255 61.875 ;
        RECT 199.455 61.555 199.715 61.875 ;
        RECT 200.375 61.555 200.635 61.875 ;
        RECT 197.615 59.515 197.875 59.835 ;
        RECT 200.435 58.815 200.575 61.555 ;
        RECT 201.355 59.495 201.495 63.255 ;
        RECT 201.295 59.175 201.555 59.495 ;
        RECT 201.815 59.155 201.955 76.855 ;
        RECT 202.275 73.435 202.415 80.255 ;
        RECT 202.215 73.115 202.475 73.435 ;
        RECT 202.275 69.015 202.415 73.115 ;
        RECT 202.215 68.695 202.475 69.015 ;
        RECT 202.735 66.635 202.875 83.065 ;
        RECT 204.515 82.635 204.775 82.955 ;
        RECT 203.135 82.295 203.395 82.615 ;
        RECT 203.195 80.235 203.335 82.295 ;
        RECT 204.575 80.575 204.715 82.635 ;
        RECT 204.055 80.255 204.315 80.575 ;
        RECT 204.515 80.255 204.775 80.575 ;
        RECT 203.135 79.915 203.395 80.235 ;
        RECT 203.195 78.195 203.335 79.915 ;
        RECT 204.115 79.895 204.255 80.255 ;
        RECT 204.055 79.575 204.315 79.895 ;
        RECT 204.115 78.875 204.255 79.575 ;
        RECT 204.055 78.555 204.315 78.875 ;
        RECT 203.135 77.875 203.395 78.195 ;
        RECT 203.195 77.595 203.335 77.875 ;
        RECT 203.195 77.455 203.795 77.595 ;
        RECT 203.135 74.135 203.395 74.455 ;
        RECT 203.195 73.630 203.335 74.135 ;
        RECT 203.125 73.260 203.405 73.630 ;
        RECT 203.135 68.870 203.395 69.015 ;
        RECT 203.125 68.500 203.405 68.870 ;
        RECT 202.675 66.315 202.935 66.635 ;
        RECT 202.735 64.165 202.875 66.315 ;
        RECT 203.135 64.165 203.395 64.255 ;
        RECT 202.735 64.025 203.395 64.165 ;
        RECT 203.135 63.935 203.395 64.025 ;
        RECT 201.755 58.835 202.015 59.155 ;
        RECT 198.995 58.495 199.255 58.815 ;
        RECT 200.375 58.495 200.635 58.815 ;
        RECT 203.655 58.670 203.795 77.455 ;
        RECT 204.055 77.195 204.315 77.515 ;
        RECT 204.115 75.475 204.255 77.195 ;
        RECT 204.575 77.175 204.715 80.255 ;
        RECT 204.515 76.855 204.775 77.175 ;
        RECT 204.055 75.155 204.315 75.475 ;
        RECT 205.035 73.395 205.175 100.575 ;
        RECT 207.795 100.295 207.935 101.675 ;
        RECT 208.195 101.335 208.455 101.655 ;
        RECT 207.735 100.150 207.995 100.295 ;
        RECT 207.725 99.780 208.005 100.150 ;
        RECT 205.955 97.175 207.475 97.315 ;
        RECT 205.955 96.895 206.095 97.175 ;
        RECT 205.895 96.575 206.155 96.895 ;
        RECT 206.355 96.805 206.615 96.895 ;
        RECT 206.355 96.665 207.015 96.805 ;
        RECT 206.355 96.575 206.615 96.665 ;
        RECT 205.435 95.895 205.695 96.215 ;
        RECT 205.495 94.515 205.635 95.895 ;
        RECT 205.435 94.195 205.695 94.515 ;
        RECT 205.955 93.915 206.095 96.575 ;
        RECT 205.495 93.775 206.095 93.915 ;
        RECT 205.495 88.475 205.635 93.775 ;
        RECT 206.355 93.175 206.615 93.495 ;
        RECT 206.415 91.455 206.555 93.175 ;
        RECT 206.355 91.135 206.615 91.455 ;
        RECT 206.875 91.365 207.015 96.665 ;
        RECT 207.335 96.555 207.475 97.175 ;
        RECT 207.275 96.235 207.535 96.555 ;
        RECT 208.255 95.195 208.395 101.335 ;
        RECT 210.095 98.935 210.235 109.225 ;
        RECT 211.875 105.075 212.135 105.395 ;
        RECT 210.495 102.355 210.755 102.675 ;
        RECT 210.955 102.355 211.215 102.675 ;
        RECT 210.555 100.295 210.695 102.355 ;
        RECT 210.495 99.975 210.755 100.295 ;
        RECT 209.575 98.615 209.835 98.935 ;
        RECT 210.035 98.615 210.295 98.935 ;
        RECT 209.635 96.895 209.775 98.615 ;
        RECT 209.575 96.575 209.835 96.895 ;
        RECT 208.655 96.465 208.915 96.555 ;
        RECT 208.655 96.325 209.315 96.465 ;
        RECT 208.655 96.235 208.915 96.325 ;
        RECT 208.195 94.875 208.455 95.195 ;
        RECT 208.655 94.875 208.915 95.195 ;
        RECT 208.715 94.515 208.855 94.875 ;
        RECT 209.175 94.515 209.315 96.325 ;
        RECT 210.035 95.895 210.295 96.215 ;
        RECT 210.095 94.515 210.235 95.895 ;
        RECT 208.655 94.195 208.915 94.515 ;
        RECT 209.115 94.195 209.375 94.515 ;
        RECT 210.035 94.195 210.295 94.515 ;
        RECT 207.275 91.365 207.535 91.455 ;
        RECT 206.875 91.225 207.535 91.365 ;
        RECT 207.275 91.135 207.535 91.225 ;
        RECT 208.195 91.135 208.455 91.455 ;
        RECT 205.895 90.455 206.155 90.775 ;
        RECT 206.355 90.455 206.615 90.775 ;
        RECT 205.955 89.075 206.095 90.455 ;
        RECT 206.415 89.755 206.555 90.455 ;
        RECT 206.355 89.435 206.615 89.755 ;
        RECT 207.735 89.435 207.995 89.755 ;
        RECT 207.795 89.155 207.935 89.435 ;
        RECT 205.895 88.755 206.155 89.075 ;
        RECT 206.875 89.015 207.935 89.155 ;
        RECT 205.495 88.335 206.095 88.475 ;
        RECT 206.355 88.415 206.615 88.735 ;
        RECT 205.435 85.695 205.695 86.015 ;
        RECT 205.495 83.635 205.635 85.695 ;
        RECT 205.435 83.315 205.695 83.635 ;
        RECT 205.955 81.595 206.095 88.335 ;
        RECT 206.415 88.055 206.555 88.415 ;
        RECT 206.355 87.735 206.615 88.055 ;
        RECT 206.875 86.015 207.015 89.015 ;
        RECT 207.275 87.735 207.535 88.055 ;
        RECT 207.335 86.015 207.475 87.735 ;
        RECT 206.815 85.695 207.075 86.015 ;
        RECT 207.275 85.695 207.535 86.015 ;
        RECT 207.735 82.295 207.995 82.615 ;
        RECT 205.895 81.275 206.155 81.595 ;
        RECT 205.955 77.515 206.095 81.275 ;
        RECT 207.795 81.255 207.935 82.295 ;
        RECT 208.255 81.255 208.395 91.135 ;
        RECT 207.735 80.935 207.995 81.255 ;
        RECT 208.195 80.935 208.455 81.255 ;
        RECT 206.355 80.595 206.615 80.915 ;
        RECT 206.415 78.875 206.555 80.595 ;
        RECT 206.355 78.555 206.615 78.875 ;
        RECT 205.895 77.195 206.155 77.515 ;
        RECT 206.815 75.155 207.075 75.475 ;
        RECT 205.035 73.255 206.095 73.395 ;
        RECT 205.955 71.735 206.095 73.255 ;
        RECT 206.875 73.095 207.015 75.155 ;
        RECT 206.815 72.775 207.075 73.095 ;
        RECT 205.895 71.415 206.155 71.735 ;
        RECT 206.355 71.415 206.615 71.735 ;
        RECT 205.955 70.715 206.095 71.415 ;
        RECT 205.895 70.395 206.155 70.715 ;
        RECT 206.415 68.190 206.555 71.415 ;
        RECT 206.875 70.035 207.015 72.775 ;
        RECT 207.795 72.755 207.935 80.935 ;
        RECT 208.715 80.235 208.855 94.195 ;
        RECT 209.575 93.515 209.835 93.835 ;
        RECT 209.115 90.455 209.375 90.775 ;
        RECT 209.175 89.075 209.315 90.455 ;
        RECT 209.115 88.755 209.375 89.075 ;
        RECT 209.115 85.015 209.375 85.335 ;
        RECT 208.655 79.915 208.915 80.235 ;
        RECT 207.735 72.435 207.995 72.755 ;
        RECT 207.735 71.755 207.995 72.075 ;
        RECT 206.815 69.715 207.075 70.035 ;
        RECT 207.795 69.550 207.935 71.755 ;
        RECT 208.195 69.715 208.455 70.035 ;
        RECT 207.725 69.180 208.005 69.550 ;
        RECT 206.345 67.820 206.625 68.190 ;
        RECT 207.725 67.140 208.005 67.510 ;
        RECT 208.255 67.315 208.395 69.715 ;
        RECT 207.735 66.995 207.995 67.140 ;
        RECT 208.195 66.995 208.455 67.315 ;
        RECT 204.505 66.460 204.785 66.830 ;
        RECT 204.575 64.255 204.715 66.460 ;
        RECT 208.655 66.315 208.915 66.635 ;
        RECT 208.185 65.100 208.465 65.470 ;
        RECT 208.255 64.255 208.395 65.100 ;
        RECT 204.515 63.935 204.775 64.255 ;
        RECT 208.195 63.935 208.455 64.255 ;
        RECT 204.055 61.215 204.315 61.535 ;
        RECT 198.075 57.815 198.335 58.135 ;
        RECT 197.145 56.940 197.425 57.310 ;
        RECT 197.215 56.775 197.355 56.940 ;
        RECT 196.695 56.455 196.955 56.775 ;
        RECT 197.155 56.455 197.415 56.775 ;
        RECT 196.235 53.735 196.495 54.055 ;
        RECT 193.935 52.715 194.195 53.035 ;
        RECT 193.475 51.015 193.735 51.335 ;
        RECT 193.995 50.655 194.135 52.715 ;
        RECT 197.215 51.675 197.355 56.455 ;
        RECT 197.155 51.355 197.415 51.675 ;
        RECT 193.935 50.335 194.195 50.655 ;
        RECT 195.315 50.565 195.575 50.655 ;
        RECT 195.315 50.425 195.975 50.565 ;
        RECT 195.315 50.335 195.575 50.425 ;
        RECT 195.835 47.595 195.975 50.425 ;
        RECT 195.775 47.275 196.035 47.595 ;
        RECT 193.935 42.515 194.195 42.835 ;
        RECT 193.015 41.495 193.275 41.815 ;
        RECT 192.555 37.075 192.815 37.395 ;
        RECT 193.995 36.795 194.135 42.515 ;
        RECT 195.835 42.495 195.975 47.275 ;
        RECT 197.215 45.555 197.355 51.355 ;
        RECT 198.135 51.335 198.275 57.815 ;
        RECT 199.055 53.375 199.195 58.495 ;
        RECT 203.585 58.300 203.865 58.670 ;
        RECT 203.655 55.835 203.795 58.300 ;
        RECT 204.115 57.115 204.255 61.215 ;
        RECT 205.895 60.535 206.155 60.855 ;
        RECT 204.515 58.495 204.775 58.815 ;
        RECT 204.055 56.795 204.315 57.115 ;
        RECT 203.655 55.695 204.255 55.835 ;
        RECT 198.535 53.055 198.795 53.375 ;
        RECT 198.995 53.055 199.255 53.375 ;
        RECT 198.075 51.015 198.335 51.335 ;
        RECT 198.595 50.565 198.735 53.055 ;
        RECT 203.595 52.715 203.855 53.035 ;
        RECT 198.135 50.425 198.735 50.565 ;
        RECT 197.155 45.235 197.415 45.555 ;
        RECT 197.215 42.835 197.355 45.235 ;
        RECT 197.615 44.895 197.875 45.215 ;
        RECT 197.675 43.515 197.815 44.895 ;
        RECT 198.135 44.535 198.275 50.425 ;
        RECT 203.655 49.975 203.795 52.715 ;
        RECT 203.595 49.655 203.855 49.975 ;
        RECT 204.115 47.595 204.255 55.695 ;
        RECT 204.575 54.395 204.715 58.495 ;
        RECT 204.975 56.795 205.235 57.115 ;
        RECT 205.035 56.630 205.175 56.795 ;
        RECT 204.965 56.260 205.245 56.630 ;
        RECT 204.515 54.075 204.775 54.395 ;
        RECT 205.955 50.655 206.095 60.535 ;
        RECT 208.715 58.475 208.855 66.315 ;
        RECT 209.175 61.535 209.315 85.015 ;
        RECT 209.635 82.615 209.775 93.515 ;
        RECT 210.095 93.495 210.235 94.195 ;
        RECT 210.035 93.175 210.295 93.495 ;
        RECT 210.035 91.135 210.295 91.455 ;
        RECT 210.095 88.735 210.235 91.135 ;
        RECT 210.035 88.415 210.295 88.735 ;
        RECT 210.035 85.355 210.295 85.675 ;
        RECT 209.575 82.295 209.835 82.615 ;
        RECT 210.095 66.975 210.235 85.355 ;
        RECT 210.555 83.975 210.695 99.975 ;
        RECT 211.015 97.915 211.155 102.355 ;
        RECT 211.935 101.655 212.075 105.075 ;
        RECT 212.395 104.715 212.535 109.225 ;
        RECT 214.175 107.795 214.435 108.115 ;
        RECT 212.335 104.395 212.595 104.715 ;
        RECT 214.235 102.675 214.375 107.795 ;
        RECT 214.175 102.355 214.435 102.675 ;
        RECT 211.875 101.335 212.135 101.655 ;
        RECT 212.335 101.335 212.595 101.655 ;
        RECT 214.175 101.335 214.435 101.655 ;
        RECT 210.955 97.595 211.215 97.915 ;
        RECT 211.935 97.235 212.075 101.335 ;
        RECT 212.395 100.635 212.535 101.335 ;
        RECT 212.335 100.315 212.595 100.635 ;
        RECT 213.715 99.635 213.975 99.955 ;
        RECT 213.255 98.955 213.515 99.275 ;
        RECT 211.875 96.915 212.135 97.235 ;
        RECT 213.315 96.215 213.455 98.955 ;
        RECT 213.255 95.895 213.515 96.215 ;
        RECT 213.775 95.275 213.915 99.635 ;
        RECT 214.235 97.915 214.375 101.335 ;
        RECT 214.695 100.635 214.835 109.225 ;
        RECT 216.015 108.135 216.275 108.455 ;
        RECT 216.075 106.075 216.215 108.135 ;
        RECT 216.995 107.775 217.135 109.225 ;
        RECT 216.935 107.455 217.195 107.775 ;
        RECT 216.935 106.775 217.195 107.095 ;
        RECT 216.015 105.755 216.275 106.075 ;
        RECT 216.995 105.395 217.135 106.775 ;
        RECT 219.295 105.735 219.435 109.225 ;
        RECT 221.595 108.455 221.735 109.225 ;
        RECT 221.535 108.135 221.795 108.455 ;
        RECT 220.945 106.240 222.485 106.610 ;
        RECT 223.895 106.075 224.035 109.225 ;
        RECT 223.835 105.755 224.095 106.075 ;
        RECT 219.235 105.415 219.495 105.735 ;
        RECT 216.935 105.075 217.195 105.395 ;
        RECT 217.395 105.075 217.655 105.395 ;
        RECT 217.455 104.795 217.595 105.075 ;
        RECT 216.995 104.655 217.595 104.795 ;
        RECT 221.075 104.735 221.335 105.055 ;
        RECT 215.095 104.055 215.355 104.375 ;
        RECT 215.155 103.355 215.295 104.055 ;
        RECT 215.095 103.035 215.355 103.355 ;
        RECT 215.155 102.675 215.295 103.035 ;
        RECT 216.475 102.695 216.735 103.015 ;
        RECT 215.095 102.355 215.355 102.675 ;
        RECT 214.635 100.315 214.895 100.635 ;
        RECT 215.555 99.635 215.815 99.955 ;
        RECT 214.175 97.595 214.435 97.915 ;
        RECT 213.775 95.135 214.375 95.275 ;
        RECT 210.955 94.195 211.215 94.515 ;
        RECT 211.015 93.835 211.155 94.195 ;
        RECT 210.955 93.515 211.215 93.835 ;
        RECT 211.875 93.175 212.135 93.495 ;
        RECT 211.405 91.620 211.685 91.990 ;
        RECT 211.415 91.475 211.675 91.620 ;
        RECT 211.935 89.075 212.075 93.175 ;
        RECT 212.335 92.155 212.595 92.475 ;
        RECT 212.395 91.795 212.535 92.155 ;
        RECT 212.335 91.475 212.595 91.795 ;
        RECT 212.795 91.135 213.055 91.455 ;
        RECT 211.875 88.755 212.135 89.075 ;
        RECT 210.955 87.735 211.215 88.055 ;
        RECT 211.415 87.735 211.675 88.055 ;
        RECT 210.495 83.655 210.755 83.975 ;
        RECT 210.555 77.855 210.695 83.655 ;
        RECT 210.495 77.535 210.755 77.855 ;
        RECT 210.555 75.135 210.695 77.535 ;
        RECT 210.495 74.815 210.755 75.135 ;
        RECT 210.495 69.035 210.755 69.355 ;
        RECT 210.035 66.655 210.295 66.975 ;
        RECT 209.575 65.975 209.835 66.295 ;
        RECT 209.635 64.255 209.775 65.975 ;
        RECT 210.555 64.255 210.695 69.035 ;
        RECT 209.575 63.935 209.835 64.255 ;
        RECT 210.495 63.935 210.755 64.255 ;
        RECT 211.015 61.875 211.155 87.735 ;
        RECT 211.475 83.635 211.615 87.735 ;
        RECT 212.855 87.035 212.995 91.135 ;
        RECT 213.245 88.220 213.525 88.590 ;
        RECT 212.795 86.715 213.055 87.035 ;
        RECT 211.865 86.180 212.145 86.550 ;
        RECT 211.935 83.635 212.075 86.180 ;
        RECT 212.855 86.015 212.995 86.715 ;
        RECT 212.795 85.695 213.055 86.015 ;
        RECT 212.335 85.015 212.595 85.335 ;
        RECT 212.395 83.975 212.535 85.015 ;
        RECT 212.335 83.655 212.595 83.975 ;
        RECT 211.415 83.315 211.675 83.635 ;
        RECT 211.875 83.315 212.135 83.635 ;
        RECT 212.325 80.740 212.605 81.110 ;
        RECT 212.395 78.195 212.535 80.740 ;
        RECT 212.795 80.595 213.055 80.915 ;
        RECT 212.855 80.430 212.995 80.595 ;
        RECT 212.785 80.060 213.065 80.430 ;
        RECT 212.335 77.875 212.595 78.195 ;
        RECT 211.875 77.535 212.135 77.855 ;
        RECT 211.415 77.195 211.675 77.515 ;
        RECT 211.475 73.395 211.615 77.195 ;
        RECT 211.935 75.475 212.075 77.535 ;
        RECT 212.335 75.835 212.595 76.155 ;
        RECT 211.875 75.155 212.135 75.475 ;
        RECT 212.395 74.990 212.535 75.835 ;
        RECT 211.875 74.475 212.135 74.795 ;
        RECT 212.325 74.620 212.605 74.990 ;
        RECT 212.335 74.475 212.595 74.620 ;
        RECT 211.935 74.195 212.075 74.475 ;
        RECT 211.935 74.055 212.535 74.195 ;
        RECT 211.475 73.255 212.075 73.395 ;
        RECT 211.415 72.095 211.675 72.415 ;
        RECT 211.475 69.695 211.615 72.095 ;
        RECT 211.415 69.375 211.675 69.695 ;
        RECT 211.475 62.070 211.615 69.375 ;
        RECT 211.935 67.315 212.075 73.255 ;
        RECT 212.395 72.415 212.535 74.055 ;
        RECT 212.335 72.095 212.595 72.415 ;
        RECT 212.335 69.375 212.595 69.695 ;
        RECT 212.395 67.655 212.535 69.375 ;
        RECT 212.785 67.820 213.065 68.190 ;
        RECT 212.795 67.675 213.055 67.820 ;
        RECT 212.335 67.335 212.595 67.655 ;
        RECT 211.875 66.995 212.135 67.315 ;
        RECT 212.395 66.975 212.535 67.335 ;
        RECT 213.315 66.975 213.455 88.220 ;
        RECT 213.705 78.700 213.985 79.070 ;
        RECT 213.715 78.555 213.975 78.700 ;
        RECT 213.715 77.875 213.975 78.195 ;
        RECT 213.775 75.815 213.915 77.875 ;
        RECT 214.235 77.175 214.375 95.135 ;
        RECT 215.095 90.455 215.355 90.775 ;
        RECT 215.155 89.415 215.295 90.455 ;
        RECT 215.095 89.095 215.355 89.415 ;
        RECT 215.615 88.645 215.755 99.635 ;
        RECT 215.155 88.505 215.755 88.645 ;
        RECT 214.635 82.295 214.895 82.615 ;
        RECT 214.175 76.855 214.435 77.175 ;
        RECT 213.715 75.495 213.975 75.815 ;
        RECT 214.235 75.670 214.375 76.855 ;
        RECT 213.775 70.375 213.915 75.495 ;
        RECT 214.165 75.300 214.445 75.670 ;
        RECT 214.175 74.815 214.435 75.135 ;
        RECT 214.235 72.755 214.375 74.815 ;
        RECT 214.175 72.435 214.435 72.755 ;
        RECT 213.715 70.055 213.975 70.375 ;
        RECT 213.715 69.375 213.975 69.695 ;
        RECT 213.775 69.015 213.915 69.375 ;
        RECT 213.715 68.925 213.975 69.015 ;
        RECT 213.715 68.785 214.375 68.925 ;
        RECT 213.715 68.695 213.975 68.785 ;
        RECT 214.235 67.315 214.375 68.785 ;
        RECT 214.175 66.995 214.435 67.315 ;
        RECT 212.335 66.655 212.595 66.975 ;
        RECT 213.255 66.655 213.515 66.975 ;
        RECT 213.715 66.655 213.975 66.975 ;
        RECT 213.255 64.615 213.515 64.935 ;
        RECT 213.315 64.255 213.455 64.615 ;
        RECT 213.775 64.255 213.915 66.655 ;
        RECT 214.175 66.315 214.435 66.635 ;
        RECT 213.255 63.935 213.515 64.255 ;
        RECT 213.715 63.935 213.975 64.255 ;
        RECT 211.875 63.255 212.135 63.575 ;
        RECT 213.775 63.430 213.915 63.935 ;
        RECT 210.035 61.555 210.295 61.875 ;
        RECT 210.955 61.555 211.215 61.875 ;
        RECT 211.405 61.700 211.685 62.070 ;
        RECT 209.115 61.215 209.375 61.535 ;
        RECT 208.655 58.155 208.915 58.475 ;
        RECT 208.655 56.115 208.915 56.435 ;
        RECT 207.275 53.395 207.535 53.715 ;
        RECT 207.335 51.335 207.475 53.395 ;
        RECT 208.715 53.375 208.855 56.115 ;
        RECT 210.095 54.395 210.235 61.555 ;
        RECT 211.935 59.835 212.075 63.255 ;
        RECT 213.705 63.060 213.985 63.430 ;
        RECT 212.335 61.555 212.595 61.875 ;
        RECT 211.875 59.515 212.135 59.835 ;
        RECT 212.395 58.815 212.535 61.555 ;
        RECT 214.235 58.815 214.375 66.315 ;
        RECT 214.695 59.495 214.835 82.295 ;
        RECT 215.155 72.325 215.295 88.505 ;
        RECT 216.535 83.830 216.675 102.695 ;
        RECT 216.995 96.555 217.135 104.655 ;
        RECT 219.695 104.055 219.955 104.375 ;
        RECT 217.645 103.520 219.185 103.890 ;
        RECT 219.755 100.635 219.895 104.055 ;
        RECT 221.135 103.355 221.275 104.735 ;
        RECT 221.075 103.035 221.335 103.355 ;
        RECT 221.135 102.755 221.275 103.035 ;
        RECT 220.215 102.615 221.275 102.755 ;
        RECT 219.695 100.315 219.955 100.635 ;
        RECT 217.645 98.080 219.185 98.450 ;
        RECT 220.215 97.915 220.355 102.615 ;
        RECT 226.195 102.335 226.335 109.225 ;
        RECT 228.495 106.075 228.635 109.225 ;
        RECT 228.895 108.135 229.155 108.455 ;
        RECT 228.435 105.755 228.695 106.075 ;
        RECT 228.955 105.395 229.095 108.135 ;
        RECT 229.815 106.775 230.075 107.095 ;
        RECT 228.895 105.075 229.155 105.395 ;
        RECT 229.875 105.055 230.015 106.775 ;
        RECT 230.795 106.075 230.935 109.225 ;
        RECT 233.095 106.075 233.235 109.225 ;
        RECT 235.395 106.075 235.535 109.225 ;
        RECT 230.735 105.755 230.995 106.075 ;
        RECT 233.035 105.755 233.295 106.075 ;
        RECT 235.335 105.755 235.595 106.075 ;
        RECT 234.415 105.075 234.675 105.395 ;
        RECT 235.335 105.305 235.595 105.395 ;
        RECT 234.935 105.165 235.595 105.305 ;
        RECT 229.815 104.735 230.075 105.055 ;
        RECT 228.895 104.395 229.155 104.715 ;
        RECT 226.135 102.015 226.395 102.335 ;
        RECT 223.835 101.675 224.095 101.995 ;
        RECT 220.945 100.800 222.485 101.170 ;
        RECT 221.075 100.150 221.335 100.295 ;
        RECT 223.895 100.150 224.035 101.675 ;
        RECT 228.955 101.655 229.095 104.395 ;
        RECT 228.895 101.335 229.155 101.655 ;
        RECT 229.355 101.335 229.615 101.655 ;
        RECT 229.415 100.150 229.555 101.335 ;
        RECT 229.875 100.635 230.015 104.735 ;
        RECT 234.475 104.375 234.615 105.075 ;
        RECT 234.415 104.055 234.675 104.375 ;
        RECT 232.575 102.015 232.835 102.335 ;
        RECT 232.635 100.635 232.775 102.015 ;
        RECT 229.815 100.315 230.075 100.635 ;
        RECT 232.575 100.315 232.835 100.635 ;
        RECT 221.065 99.780 221.345 100.150 ;
        RECT 223.825 99.780 224.105 100.150 ;
        RECT 220.155 97.595 220.415 97.915 ;
        RECT 221.525 97.740 221.805 98.110 ;
        RECT 221.595 96.895 221.735 97.740 ;
        RECT 221.535 96.575 221.795 96.895 ;
        RECT 222.915 96.750 223.175 96.895 ;
        RECT 216.935 96.235 217.195 96.555 ;
        RECT 222.905 96.380 223.185 96.750 ;
        RECT 220.945 95.360 222.485 95.730 ;
        RECT 217.645 92.640 219.185 93.010 ;
        RECT 216.935 91.135 217.195 91.455 ;
        RECT 216.465 83.460 216.745 83.830 ;
        RECT 215.555 82.635 215.815 82.955 ;
        RECT 215.615 74.875 215.755 82.635 ;
        RECT 216.015 82.295 216.275 82.615 ;
        RECT 216.075 81.595 216.215 82.295 ;
        RECT 216.015 81.275 216.275 81.595 ;
        RECT 216.535 78.875 216.675 83.460 ;
        RECT 216.015 78.555 216.275 78.875 ;
        RECT 216.475 78.555 216.735 78.875 ;
        RECT 216.075 77.595 216.215 78.555 ;
        RECT 216.075 77.455 216.675 77.595 ;
        RECT 216.015 76.855 216.275 77.175 ;
        RECT 216.075 75.475 216.215 76.855 ;
        RECT 216.015 75.155 216.275 75.475 ;
        RECT 215.615 74.735 216.215 74.875 ;
        RECT 215.555 74.135 215.815 74.455 ;
        RECT 215.615 73.095 215.755 74.135 ;
        RECT 215.555 72.775 215.815 73.095 ;
        RECT 215.555 72.325 215.815 72.415 ;
        RECT 215.155 72.185 215.815 72.325 ;
        RECT 215.555 72.095 215.815 72.185 ;
        RECT 215.095 67.675 215.355 67.995 ;
        RECT 214.635 59.175 214.895 59.495 ;
        RECT 215.155 59.155 215.295 67.675 ;
        RECT 215.545 65.100 215.825 65.470 ;
        RECT 215.615 64.935 215.755 65.100 ;
        RECT 215.555 64.615 215.815 64.935 ;
        RECT 215.555 63.935 215.815 64.255 ;
        RECT 215.615 62.555 215.755 63.935 ;
        RECT 215.555 62.235 215.815 62.555 ;
        RECT 216.075 61.875 216.215 74.735 ;
        RECT 216.535 72.950 216.675 77.455 ;
        RECT 216.465 72.580 216.745 72.950 ;
        RECT 216.475 66.995 216.735 67.315 ;
        RECT 216.535 65.275 216.675 66.995 ;
        RECT 216.475 64.955 216.735 65.275 ;
        RECT 216.995 65.185 217.135 91.135 ;
        RECT 220.945 89.920 222.485 90.290 ;
        RECT 217.645 87.200 219.185 87.570 ;
        RECT 223.895 86.435 224.035 99.780 ;
        RECT 226.135 99.635 226.395 99.955 ;
        RECT 228.435 99.635 228.695 99.955 ;
        RECT 229.345 99.780 229.625 100.150 ;
        RECT 226.195 97.915 226.335 99.635 ;
        RECT 228.495 99.470 228.635 99.635 ;
        RECT 228.425 99.100 228.705 99.470 ;
        RECT 226.135 97.595 226.395 97.915 ;
        RECT 228.495 96.895 228.635 99.100 ;
        RECT 229.415 98.935 229.555 99.780 ;
        RECT 229.355 98.615 229.615 98.935 ;
        RECT 229.355 97.595 229.615 97.915 ;
        RECT 225.675 96.575 225.935 96.895 ;
        RECT 226.595 96.575 226.855 96.895 ;
        RECT 228.435 96.575 228.695 96.895 ;
        RECT 225.215 94.875 225.475 95.195 ;
        RECT 224.755 94.535 225.015 94.855 ;
        RECT 224.295 93.175 224.555 93.495 ;
        RECT 224.355 91.115 224.495 93.175 ;
        RECT 224.295 90.795 224.555 91.115 ;
        RECT 222.975 86.295 224.035 86.435 ;
        RECT 217.395 85.355 217.655 85.675 ;
        RECT 217.455 83.635 217.595 85.355 ;
        RECT 220.945 84.480 222.485 84.850 ;
        RECT 220.155 83.655 220.415 83.975 ;
        RECT 217.395 83.315 217.655 83.635 ;
        RECT 217.645 81.760 219.185 82.130 ;
        RECT 217.395 80.430 217.655 80.575 ;
        RECT 217.385 80.315 217.665 80.430 ;
        RECT 217.385 80.175 218.515 80.315 ;
        RECT 217.385 80.060 217.665 80.175 ;
        RECT 217.845 78.700 218.125 79.070 ;
        RECT 217.915 78.535 218.055 78.700 ;
        RECT 217.855 78.215 218.115 78.535 ;
        RECT 218.375 77.515 218.515 80.175 ;
        RECT 219.235 78.555 219.495 78.875 ;
        RECT 218.315 77.195 218.575 77.515 ;
        RECT 219.295 77.085 219.435 78.555 ;
        RECT 220.215 78.195 220.355 83.655 ;
        RECT 220.945 79.040 222.485 79.410 ;
        RECT 220.155 77.875 220.415 78.195 ;
        RECT 219.295 76.945 219.895 77.085 ;
        RECT 217.645 76.320 219.185 76.690 ;
        RECT 219.755 76.155 219.895 76.945 ;
        RECT 219.695 75.835 219.955 76.155 ;
        RECT 218.315 75.155 218.575 75.475 ;
        RECT 218.375 74.795 218.515 75.155 ;
        RECT 222.975 74.795 223.115 86.295 ;
        RECT 223.375 85.695 223.635 86.015 ;
        RECT 223.435 79.895 223.575 85.695 ;
        RECT 224.815 85.675 224.955 94.535 ;
        RECT 225.275 93.835 225.415 94.875 ;
        RECT 225.215 93.515 225.475 93.835 ;
        RECT 225.735 91.115 225.875 96.575 ;
        RECT 226.135 94.195 226.395 94.515 ;
        RECT 226.195 92.475 226.335 94.195 ;
        RECT 226.135 92.155 226.395 92.475 ;
        RECT 225.675 90.795 225.935 91.115 ;
        RECT 225.735 89.075 225.875 90.795 ;
        RECT 225.675 88.755 225.935 89.075 ;
        RECT 224.755 85.355 225.015 85.675 ;
        RECT 224.295 81.275 224.555 81.595 ;
        RECT 223.375 79.575 223.635 79.895 ;
        RECT 218.315 74.475 218.575 74.795 ;
        RECT 222.915 74.475 223.175 74.795 ;
        RECT 220.155 74.135 220.415 74.455 ;
        RECT 220.215 72.950 220.355 74.135 ;
        RECT 220.945 73.600 222.485 73.970 ;
        RECT 222.975 73.095 223.115 74.475 ;
        RECT 220.145 72.580 220.425 72.950 ;
        RECT 222.915 72.775 223.175 73.095 ;
        RECT 217.645 70.880 219.185 71.250 ;
        RECT 219.695 70.395 219.955 70.715 ;
        RECT 217.395 70.055 217.655 70.375 ;
        RECT 217.455 67.315 217.595 70.055 ;
        RECT 218.775 68.695 219.035 69.015 ;
        RECT 219.755 68.870 219.895 70.395 ;
        RECT 220.155 69.715 220.415 70.035 ;
        RECT 217.845 67.820 218.125 68.190 ;
        RECT 217.915 67.315 218.055 67.820 ;
        RECT 218.315 67.675 218.575 67.995 ;
        RECT 218.375 67.510 218.515 67.675 ;
        RECT 217.395 66.995 217.655 67.315 ;
        RECT 217.855 66.995 218.115 67.315 ;
        RECT 218.305 67.140 218.585 67.510 ;
        RECT 218.835 67.315 218.975 68.695 ;
        RECT 219.685 68.500 219.965 68.870 ;
        RECT 218.775 66.995 219.035 67.315 ;
        RECT 219.235 67.225 219.495 67.315 ;
        RECT 219.235 67.085 219.895 67.225 ;
        RECT 219.235 66.995 219.495 67.085 ;
        RECT 217.455 66.635 217.595 66.995 ;
        RECT 217.395 66.315 217.655 66.635 ;
        RECT 217.645 65.440 219.185 65.810 ;
        RECT 216.995 65.045 217.595 65.185 ;
        RECT 217.455 64.675 217.595 65.045 ;
        RECT 217.455 64.535 218.055 64.675 ;
        RECT 219.755 64.595 219.895 67.085 ;
        RECT 217.395 63.935 217.655 64.255 ;
        RECT 216.475 63.255 216.735 63.575 ;
        RECT 217.455 63.430 217.595 63.935 ;
        RECT 215.555 61.555 215.815 61.875 ;
        RECT 216.015 61.555 216.275 61.875 ;
        RECT 216.535 61.785 216.675 63.255 ;
        RECT 217.385 63.060 217.665 63.430 ;
        RECT 216.935 61.785 217.195 61.875 ;
        RECT 216.535 61.645 217.195 61.785 ;
        RECT 216.935 61.555 217.195 61.645 ;
        RECT 215.615 59.235 215.755 61.555 ;
        RECT 216.475 60.875 216.735 61.195 ;
        RECT 216.935 60.875 217.195 61.195 ;
        RECT 215.095 58.835 215.355 59.155 ;
        RECT 215.615 59.095 216.215 59.235 ;
        RECT 212.335 58.495 212.595 58.815 ;
        RECT 214.175 58.495 214.435 58.815 ;
        RECT 214.635 58.495 214.895 58.815 ;
        RECT 213.715 58.155 213.975 58.475 ;
        RECT 212.335 57.815 212.595 58.135 ;
        RECT 210.955 55.775 211.215 56.095 ;
        RECT 211.015 54.395 211.155 55.775 ;
        RECT 210.035 54.075 210.295 54.395 ;
        RECT 210.955 54.075 211.215 54.395 ;
        RECT 208.655 53.055 208.915 53.375 ;
        RECT 212.395 53.035 212.535 57.815 ;
        RECT 210.495 52.715 210.755 53.035 ;
        RECT 212.335 52.715 212.595 53.035 ;
        RECT 210.555 51.675 210.695 52.715 ;
        RECT 213.775 51.675 213.915 58.155 ;
        RECT 214.695 55.415 214.835 58.495 ;
        RECT 215.095 57.815 215.355 58.135 ;
        RECT 214.635 55.095 214.895 55.415 ;
        RECT 214.175 52.375 214.435 52.695 ;
        RECT 210.495 51.355 210.755 51.675 ;
        RECT 213.715 51.355 213.975 51.675 ;
        RECT 214.235 51.335 214.375 52.375 ;
        RECT 207.275 51.015 207.535 51.335 ;
        RECT 210.945 50.820 211.225 51.190 ;
        RECT 212.335 51.015 212.595 51.335 ;
        RECT 214.175 51.015 214.435 51.335 ;
        RECT 214.635 51.015 214.895 51.335 ;
        RECT 205.895 50.335 206.155 50.655 ;
        RECT 211.015 49.975 211.155 50.820 ;
        RECT 210.955 49.655 211.215 49.975 ;
        RECT 211.415 49.655 211.675 49.975 ;
        RECT 204.055 47.275 204.315 47.595 ;
        RECT 211.475 47.255 211.615 49.655 ;
        RECT 212.395 47.595 212.535 51.015 ;
        RECT 214.695 48.955 214.835 51.015 ;
        RECT 214.635 48.635 214.895 48.955 ;
        RECT 214.175 48.355 214.435 48.615 ;
        RECT 215.155 48.355 215.295 57.815 ;
        RECT 216.075 56.775 216.215 59.095 ;
        RECT 216.015 56.455 216.275 56.775 ;
        RECT 215.555 56.115 215.815 56.435 ;
        RECT 215.615 48.955 215.755 56.115 ;
        RECT 215.555 48.635 215.815 48.955 ;
        RECT 214.175 48.295 215.295 48.355 ;
        RECT 214.235 48.215 215.295 48.295 ;
        RECT 216.535 47.675 216.675 60.875 ;
        RECT 216.995 58.815 217.135 60.875 ;
        RECT 217.915 60.855 218.055 64.535 ;
        RECT 219.695 64.275 219.955 64.595 ;
        RECT 218.775 63.935 219.035 64.255 ;
        RECT 218.835 62.555 218.975 63.935 ;
        RECT 219.235 63.255 219.495 63.575 ;
        RECT 219.695 63.255 219.955 63.575 ;
        RECT 218.775 62.235 219.035 62.555 ;
        RECT 219.295 62.215 219.435 63.255 ;
        RECT 219.235 61.895 219.495 62.215 ;
        RECT 219.755 61.535 219.895 63.255 ;
        RECT 219.695 61.215 219.955 61.535 ;
        RECT 220.215 61.275 220.355 69.715 ;
        RECT 220.945 68.160 222.485 68.530 ;
        RECT 220.615 67.335 220.875 67.655 ;
        RECT 220.675 64.255 220.815 67.335 ;
        RECT 222.915 66.315 223.175 66.635 ;
        RECT 221.075 64.955 221.335 65.275 ;
        RECT 221.135 64.595 221.275 64.955 ;
        RECT 221.075 64.275 221.335 64.595 ;
        RECT 220.615 63.935 220.875 64.255 ;
        RECT 220.945 62.720 222.485 63.090 ;
        RECT 222.455 61.555 222.715 61.875 ;
        RECT 220.215 61.135 220.815 61.275 ;
        RECT 217.855 60.535 218.115 60.855 ;
        RECT 220.155 60.535 220.415 60.855 ;
        RECT 217.645 60.000 219.185 60.370 ;
        RECT 216.935 58.495 217.195 58.815 ;
        RECT 218.315 58.155 218.575 58.475 ;
        RECT 217.395 57.815 217.655 58.135 ;
        RECT 217.455 55.835 217.595 57.815 ;
        RECT 218.375 56.095 218.515 58.155 ;
        RECT 220.215 57.195 220.355 60.535 ;
        RECT 220.675 59.835 220.815 61.135 ;
        RECT 222.515 59.835 222.655 61.555 ;
        RECT 220.615 59.515 220.875 59.835 ;
        RECT 222.455 59.515 222.715 59.835 ;
        RECT 221.075 58.835 221.335 59.155 ;
        RECT 220.615 58.385 220.875 58.475 ;
        RECT 221.135 58.385 221.275 58.835 ;
        RECT 222.975 58.475 223.115 66.315 ;
        RECT 220.615 58.245 221.275 58.385 ;
        RECT 220.615 58.155 220.875 58.245 ;
        RECT 222.915 58.155 223.175 58.475 ;
        RECT 220.945 57.280 222.485 57.650 ;
        RECT 220.215 57.055 220.815 57.195 ;
        RECT 220.675 56.775 220.815 57.055 ;
        RECT 220.155 56.455 220.415 56.775 ;
        RECT 220.615 56.455 220.875 56.775 ;
        RECT 218.775 56.115 219.035 56.435 ;
        RECT 216.075 47.595 216.675 47.675 ;
        RECT 212.335 47.275 212.595 47.595 ;
        RECT 216.015 47.535 216.675 47.595 ;
        RECT 216.995 55.695 217.595 55.835 ;
        RECT 218.315 55.775 218.575 56.095 ;
        RECT 216.015 47.275 216.275 47.535 ;
        RECT 204.975 46.935 205.235 47.255 ;
        RECT 211.415 46.935 211.675 47.255 ;
        RECT 216.475 46.935 216.735 47.255 ;
        RECT 205.035 46.235 205.175 46.935 ;
        RECT 204.975 45.915 205.235 46.235 ;
        RECT 208.655 45.575 208.915 45.895 ;
        RECT 205.895 44.895 206.155 45.215 ;
        RECT 202.675 44.555 202.935 44.875 ;
        RECT 198.075 44.215 198.335 44.535 ;
        RECT 197.615 43.195 197.875 43.515 ;
        RECT 197.155 42.515 197.415 42.835 ;
        RECT 195.775 42.175 196.035 42.495 ;
        RECT 194.395 41.495 194.655 41.815 ;
        RECT 193.535 36.655 194.135 36.795 ;
        RECT 194.455 36.715 194.595 41.495 ;
        RECT 195.835 39.775 195.975 42.175 ;
        RECT 196.235 41.495 196.495 41.815 ;
        RECT 196.295 40.795 196.435 41.495 ;
        RECT 197.215 40.795 197.355 42.515 ;
        RECT 196.235 40.475 196.495 40.795 ;
        RECT 197.155 40.475 197.415 40.795 ;
        RECT 197.675 40.455 197.815 43.195 ;
        RECT 198.135 41.815 198.275 44.215 ;
        RECT 202.735 42.835 202.875 44.555 ;
        RECT 202.675 42.515 202.935 42.835 ;
        RECT 198.075 41.495 198.335 41.815 ;
        RECT 197.615 40.135 197.875 40.455 ;
        RECT 198.535 40.135 198.795 40.455 ;
        RECT 195.775 39.455 196.035 39.775 ;
        RECT 197.615 39.455 197.875 39.775 ;
        RECT 195.835 37.395 195.975 39.455 ;
        RECT 197.675 37.395 197.815 39.455 ;
        RECT 198.595 37.735 198.735 40.135 ;
        RECT 202.215 39.115 202.475 39.435 ;
        RECT 198.535 37.415 198.795 37.735 ;
        RECT 195.775 37.075 196.035 37.395 ;
        RECT 197.155 37.075 197.415 37.395 ;
        RECT 197.615 37.075 197.875 37.395 ;
        RECT 195.315 36.735 195.575 37.055 ;
        RECT 193.535 36.375 193.675 36.655 ;
        RECT 194.395 36.395 194.655 36.715 ;
        RECT 193.475 36.055 193.735 36.375 ;
        RECT 193.935 36.055 194.195 36.375 ;
        RECT 193.475 34.695 193.735 35.015 ;
        RECT 193.535 30.935 193.675 34.695 ;
        RECT 193.995 33.655 194.135 36.055 ;
        RECT 193.935 33.335 194.195 33.655 ;
        RECT 193.995 31.275 194.135 33.335 ;
        RECT 193.935 30.955 194.195 31.275 ;
        RECT 193.475 30.615 193.735 30.935 ;
        RECT 193.535 29.915 193.675 30.615 ;
        RECT 195.375 29.915 195.515 36.735 ;
        RECT 197.215 34.335 197.355 37.075 ;
        RECT 197.675 35.355 197.815 37.075 ;
        RECT 197.615 35.035 197.875 35.355 ;
        RECT 197.155 34.015 197.415 34.335 ;
        RECT 197.215 31.615 197.355 34.015 ;
        RECT 197.155 31.295 197.415 31.615 ;
        RECT 198.595 31.275 198.735 37.415 ;
        RECT 202.275 35.015 202.415 39.115 ;
        RECT 205.955 37.055 206.095 44.895 ;
        RECT 208.195 42.175 208.455 42.495 ;
        RECT 207.735 39.455 207.995 39.775 ;
        RECT 207.795 38.075 207.935 39.455 ;
        RECT 207.735 37.755 207.995 38.075 ;
        RECT 205.895 36.735 206.155 37.055 ;
        RECT 205.895 36.055 206.155 36.375 ;
        RECT 205.955 35.355 206.095 36.055 ;
        RECT 205.895 35.035 206.155 35.355 ;
        RECT 202.215 34.695 202.475 35.015 ;
        RECT 199.915 34.015 200.175 34.335 ;
        RECT 198.535 30.955 198.795 31.275 ;
        RECT 199.455 30.615 199.715 30.935 ;
        RECT 193.475 29.595 193.735 29.915 ;
        RECT 195.315 29.595 195.575 29.915 ;
        RECT 199.515 29.575 199.655 30.615 ;
        RECT 199.975 29.915 200.115 34.015 ;
        RECT 205.955 32.635 206.095 35.035 ;
        RECT 208.255 35.015 208.395 42.175 ;
        RECT 208.715 36.715 208.855 45.575 ;
        RECT 211.475 45.555 211.615 46.935 ;
        RECT 216.535 45.555 216.675 46.935 ;
        RECT 216.995 45.635 217.135 55.695 ;
        RECT 218.835 55.415 218.975 56.115 ;
        RECT 218.775 55.095 219.035 55.415 ;
        RECT 219.695 55.095 219.955 55.415 ;
        RECT 217.645 54.560 219.185 54.930 ;
        RECT 219.755 54.395 219.895 55.095 ;
        RECT 219.695 54.075 219.955 54.395 ;
        RECT 220.215 53.715 220.355 56.455 ;
        RECT 220.155 53.395 220.415 53.715 ;
        RECT 223.435 53.625 223.575 79.575 ;
        RECT 223.835 76.855 224.095 77.175 ;
        RECT 223.895 61.535 224.035 76.855 ;
        RECT 224.355 73.395 224.495 81.275 ;
        RECT 226.195 81.255 226.335 92.155 ;
        RECT 226.655 91.365 226.795 96.575 ;
        RECT 228.895 96.235 229.155 96.555 ;
        RECT 227.055 95.895 227.315 96.215 ;
        RECT 227.115 92.135 227.255 95.895 ;
        RECT 227.515 94.195 227.775 94.515 ;
        RECT 227.575 93.835 227.715 94.195 ;
        RECT 227.515 93.515 227.775 93.835 ;
        RECT 228.435 93.515 228.695 93.835 ;
        RECT 227.055 91.815 227.315 92.135 ;
        RECT 228.495 91.455 228.635 93.515 ;
        RECT 228.955 92.475 229.095 96.235 ;
        RECT 228.895 92.155 229.155 92.475 ;
        RECT 229.415 91.795 229.555 97.595 ;
        RECT 229.875 92.135 230.015 100.315 ;
        RECT 230.275 99.635 230.535 99.955 ;
        RECT 230.335 99.470 230.475 99.635 ;
        RECT 230.265 99.100 230.545 99.470 ;
        RECT 230.335 94.515 230.475 99.100 ;
        RECT 231.195 98.615 231.455 98.935 ;
        RECT 230.275 94.195 230.535 94.515 ;
        RECT 230.275 93.175 230.535 93.495 ;
        RECT 229.815 91.815 230.075 92.135 ;
        RECT 229.355 91.475 229.615 91.795 ;
        RECT 226.655 91.225 227.255 91.365 ;
        RECT 226.585 88.900 226.865 89.270 ;
        RECT 226.655 83.635 226.795 88.900 ;
        RECT 226.595 83.315 226.855 83.635 ;
        RECT 225.215 80.935 225.475 81.255 ;
        RECT 226.135 80.935 226.395 81.255 ;
        RECT 225.275 80.575 225.415 80.935 ;
        RECT 227.115 80.575 227.255 91.225 ;
        RECT 228.435 91.135 228.695 91.455 ;
        RECT 228.895 90.795 229.155 91.115 ;
        RECT 228.955 85.335 229.095 90.795 ;
        RECT 229.415 87.115 229.555 91.475 ;
        RECT 229.875 91.455 230.015 91.815 ;
        RECT 229.815 91.135 230.075 91.455 ;
        RECT 230.335 88.055 230.475 93.175 ;
        RECT 231.255 91.310 231.395 98.615 ;
        RECT 232.565 98.420 232.845 98.790 ;
        RECT 232.635 97.235 232.775 98.420 ;
        RECT 232.575 96.915 232.835 97.235 ;
        RECT 232.115 94.875 232.375 95.195 ;
        RECT 231.185 90.940 231.465 91.310 ;
        RECT 231.655 91.135 231.915 91.455 ;
        RECT 230.735 90.455 230.995 90.775 ;
        RECT 231.195 90.455 231.455 90.775 ;
        RECT 230.795 89.075 230.935 90.455 ;
        RECT 231.255 89.075 231.395 90.455 ;
        RECT 230.735 88.755 230.995 89.075 ;
        RECT 231.195 88.755 231.455 89.075 ;
        RECT 230.275 87.735 230.535 88.055 ;
        RECT 229.415 86.975 230.475 87.115 ;
        RECT 229.355 85.355 229.615 85.675 ;
        RECT 228.895 85.015 229.155 85.335 ;
        RECT 228.955 84.395 229.095 85.015 ;
        RECT 228.035 84.255 229.095 84.395 ;
        RECT 227.515 83.655 227.775 83.975 ;
        RECT 225.215 80.255 225.475 80.575 ;
        RECT 227.055 80.255 227.315 80.575 ;
        RECT 227.115 79.750 227.255 80.255 ;
        RECT 227.575 80.235 227.715 83.655 ;
        RECT 228.035 83.635 228.175 84.255 ;
        RECT 227.975 83.315 228.235 83.635 ;
        RECT 228.425 83.460 228.705 83.830 ;
        RECT 229.415 83.635 229.555 85.355 ;
        RECT 229.815 85.015 230.075 85.335 ;
        RECT 228.435 83.315 228.695 83.460 ;
        RECT 229.355 83.315 229.615 83.635 ;
        RECT 228.435 82.635 228.695 82.955 ;
        RECT 227.975 82.295 228.235 82.615 ;
        RECT 227.515 79.915 227.775 80.235 ;
        RECT 227.045 79.380 227.325 79.750 ;
        RECT 227.575 78.535 227.715 79.915 ;
        RECT 227.515 78.215 227.775 78.535 ;
        RECT 225.215 74.815 225.475 75.135 ;
        RECT 224.355 73.255 224.955 73.395 ;
        RECT 223.835 61.215 224.095 61.535 ;
        RECT 223.835 60.535 224.095 60.855 ;
        RECT 223.895 58.815 224.035 60.535 ;
        RECT 223.835 58.495 224.095 58.815 ;
        RECT 224.295 55.270 224.555 55.415 ;
        RECT 224.285 54.900 224.565 55.270 ;
        RECT 222.975 53.485 223.575 53.625 ;
        RECT 218.775 53.055 219.035 53.375 ;
        RECT 218.835 51.335 218.975 53.055 ;
        RECT 218.775 51.015 219.035 51.335 ;
        RECT 219.695 51.015 219.955 51.335 ;
        RECT 217.645 49.120 219.185 49.490 ;
        RECT 219.235 48.185 219.495 48.275 ;
        RECT 219.755 48.185 219.895 51.015 ;
        RECT 220.215 50.995 220.355 53.395 ;
        RECT 220.945 51.840 222.485 52.210 ;
        RECT 220.155 50.675 220.415 50.995 ;
        RECT 219.235 48.045 219.895 48.185 ;
        RECT 219.235 47.955 219.495 48.045 ;
        RECT 211.415 45.235 211.675 45.555 ;
        RECT 216.475 45.235 216.735 45.555 ;
        RECT 216.995 45.495 218.055 45.635 ;
        RECT 217.915 45.215 218.055 45.495 ;
        RECT 214.635 44.895 214.895 45.215 ;
        RECT 217.855 44.895 218.115 45.215 ;
        RECT 212.795 44.555 213.055 44.875 ;
        RECT 210.035 44.215 210.295 44.535 ;
        RECT 210.095 43.175 210.235 44.215 ;
        RECT 212.855 43.515 212.995 44.555 ;
        RECT 213.255 44.215 213.515 44.535 ;
        RECT 213.315 43.515 213.455 44.215 ;
        RECT 212.795 43.195 213.055 43.515 ;
        RECT 213.255 43.195 213.515 43.515 ;
        RECT 210.035 42.855 210.295 43.175 ;
        RECT 211.875 42.855 212.135 43.175 ;
        RECT 211.935 40.795 212.075 42.855 ;
        RECT 212.855 41.815 212.995 43.195 ;
        RECT 212.795 41.495 213.055 41.815 ;
        RECT 211.875 40.475 212.135 40.795 ;
        RECT 214.695 39.095 214.835 44.895 ;
        RECT 217.645 43.680 219.185 44.050 ;
        RECT 219.755 42.915 219.895 48.045 ;
        RECT 220.215 47.255 220.355 50.675 ;
        RECT 220.615 49.655 220.875 49.975 ;
        RECT 220.675 47.255 220.815 49.655 ;
        RECT 220.155 46.935 220.415 47.255 ;
        RECT 220.615 46.935 220.875 47.255 ;
        RECT 220.945 46.400 222.485 46.770 ;
        RECT 222.975 43.515 223.115 53.485 ;
        RECT 223.375 52.715 223.635 53.035 ;
        RECT 223.435 51.335 223.575 52.715 ;
        RECT 223.375 51.015 223.635 51.335 ;
        RECT 222.915 43.195 223.175 43.515 ;
        RECT 218.835 42.835 219.895 42.915 ;
        RECT 218.775 42.775 219.895 42.835 ;
        RECT 218.775 42.515 219.035 42.775 ;
        RECT 217.455 42.155 218.055 42.235 ;
        RECT 217.395 42.095 218.115 42.155 ;
        RECT 217.395 41.835 217.655 42.095 ;
        RECT 217.855 41.835 218.115 42.095 ;
        RECT 217.915 40.455 218.055 41.835 ;
        RECT 219.755 40.795 219.895 42.775 ;
        RECT 222.975 42.495 223.115 43.195 ;
        RECT 222.915 42.175 223.175 42.495 ;
        RECT 220.945 40.960 222.485 41.330 ;
        RECT 224.815 40.795 224.955 73.255 ;
        RECT 225.275 61.955 225.415 74.815 ;
        RECT 228.035 72.270 228.175 82.295 ;
        RECT 228.495 77.175 228.635 82.635 ;
        RECT 229.345 81.420 229.625 81.790 ;
        RECT 229.415 81.255 229.555 81.420 ;
        RECT 229.875 81.255 230.015 85.015 ;
        RECT 229.355 80.935 229.615 81.255 ;
        RECT 229.815 80.935 230.075 81.255 ;
        RECT 228.895 79.575 229.155 79.895 ;
        RECT 228.955 77.515 229.095 79.575 ;
        RECT 229.415 78.875 229.555 80.935 ;
        RECT 229.805 80.060 230.085 80.430 ;
        RECT 230.335 80.145 230.475 86.975 ;
        RECT 231.715 85.075 231.855 91.135 ;
        RECT 232.175 91.115 232.315 94.875 ;
        RECT 232.635 91.455 232.775 96.915 ;
        RECT 233.955 92.155 234.215 92.475 ;
        RECT 233.495 91.815 233.755 92.135 ;
        RECT 233.555 91.455 233.695 91.815 ;
        RECT 232.575 91.135 232.835 91.455 ;
        RECT 233.495 91.135 233.755 91.455 ;
        RECT 232.115 90.795 232.375 91.115 ;
        RECT 232.175 88.055 232.315 90.795 ;
        RECT 232.115 87.735 232.375 88.055 ;
        RECT 231.255 84.935 231.855 85.075 ;
        RECT 231.255 82.955 231.395 84.935 ;
        RECT 231.655 83.995 231.915 84.315 ;
        RECT 231.195 82.635 231.455 82.955 ;
        RECT 230.735 80.145 230.995 80.235 ;
        RECT 229.815 79.915 230.075 80.060 ;
        RECT 230.335 80.005 230.995 80.145 ;
        RECT 230.735 79.915 230.995 80.005 ;
        RECT 229.355 78.555 229.615 78.875 ;
        RECT 228.895 77.195 229.155 77.515 ;
        RECT 228.435 76.855 228.695 77.175 ;
        RECT 229.355 75.495 229.615 75.815 ;
        RECT 228.895 72.775 229.155 73.095 ;
        RECT 227.965 71.900 228.245 72.270 ;
        RECT 228.035 67.315 228.175 71.900 ;
        RECT 228.955 70.375 229.095 72.775 ;
        RECT 228.895 70.055 229.155 70.375 ;
        RECT 229.415 69.355 229.555 75.495 ;
        RECT 229.875 72.755 230.015 79.915 ;
        RECT 230.795 79.070 230.935 79.915 ;
        RECT 230.725 78.700 231.005 79.070 ;
        RECT 230.795 77.175 230.935 78.700 ;
        RECT 231.195 78.215 231.455 78.535 ;
        RECT 230.735 76.855 230.995 77.175 ;
        RECT 231.255 74.455 231.395 78.215 ;
        RECT 231.195 74.135 231.455 74.455 ;
        RECT 229.815 72.435 230.075 72.755 ;
        RECT 230.735 72.435 230.995 72.755 ;
        RECT 230.795 72.075 230.935 72.435 ;
        RECT 230.735 71.755 230.995 72.075 ;
        RECT 230.275 70.395 230.535 70.715 ;
        RECT 229.355 69.035 229.615 69.355 ;
        RECT 227.975 66.995 228.235 67.315 ;
        RECT 228.435 66.655 228.695 66.975 ;
        RECT 226.135 65.975 226.395 66.295 ;
        RECT 226.195 64.255 226.335 65.975 ;
        RECT 228.495 65.275 228.635 66.655 ;
        RECT 228.435 64.955 228.695 65.275 ;
        RECT 226.135 63.935 226.395 64.255 ;
        RECT 230.335 62.215 230.475 70.395 ;
        RECT 230.795 67.995 230.935 71.755 ;
        RECT 230.735 67.675 230.995 67.995 ;
        RECT 231.255 62.555 231.395 74.135 ;
        RECT 231.715 70.375 231.855 83.995 ;
        RECT 232.115 79.575 232.375 79.895 ;
        RECT 232.175 77.855 232.315 79.575 ;
        RECT 232.115 77.535 232.375 77.855 ;
        RECT 232.635 75.385 232.775 91.135 ;
        RECT 234.015 85.925 234.155 92.155 ;
        RECT 234.415 88.075 234.675 88.395 ;
        RECT 234.475 86.550 234.615 88.075 ;
        RECT 234.405 86.180 234.685 86.550 ;
        RECT 234.015 85.785 234.615 85.925 ;
        RECT 233.035 82.295 233.295 82.615 ;
        RECT 233.495 82.295 233.755 82.615 ;
        RECT 233.095 80.575 233.235 82.295 ;
        RECT 233.555 80.915 233.695 82.295 ;
        RECT 233.495 80.595 233.755 80.915 ;
        RECT 234.475 80.575 234.615 85.785 ;
        RECT 234.935 84.315 235.075 105.165 ;
        RECT 235.335 105.075 235.595 105.165 ;
        RECT 235.855 96.555 235.995 109.495 ;
        RECT 237.625 109.225 237.905 128.720 ;
        RECT 239.925 109.225 240.205 129.300 ;
        RECT 242.225 109.225 242.505 129.880 ;
        RECT 237.695 106.075 237.835 109.225 ;
        RECT 239.015 107.795 239.275 108.115 ;
        RECT 237.635 105.755 237.895 106.075 ;
        RECT 239.075 105.395 239.215 107.795 ;
        RECT 239.015 105.075 239.275 105.395 ;
        RECT 238.555 104.735 238.815 105.055 ;
        RECT 237.175 104.055 237.435 104.375 ;
        RECT 238.095 104.055 238.355 104.375 ;
        RECT 235.795 96.235 236.055 96.555 ;
        RECT 234.875 83.995 235.135 84.315 ;
        RECT 233.035 80.255 233.295 80.575 ;
        RECT 233.955 80.255 234.215 80.575 ;
        RECT 234.415 80.255 234.675 80.575 ;
        RECT 233.495 79.915 233.755 80.235 ;
        RECT 233.035 77.195 233.295 77.515 ;
        RECT 232.175 75.245 232.775 75.385 ;
        RECT 232.175 72.755 232.315 75.245 ;
        RECT 232.575 74.475 232.835 74.795 ;
        RECT 232.635 73.435 232.775 74.475 ;
        RECT 232.575 73.115 232.835 73.435 ;
        RECT 232.115 72.435 232.375 72.755 ;
        RECT 231.655 70.055 231.915 70.375 ;
        RECT 231.195 62.235 231.455 62.555 ;
        RECT 225.275 61.815 226.335 61.955 ;
        RECT 230.275 61.895 230.535 62.215 ;
        RECT 231.715 61.875 231.855 70.055 ;
        RECT 233.095 69.015 233.235 77.195 ;
        RECT 233.555 77.175 233.695 79.915 ;
        RECT 233.495 76.855 233.755 77.175 ;
        RECT 234.015 73.395 234.155 80.255 ;
        RECT 236.715 75.835 236.975 76.155 ;
        RECT 236.255 74.135 236.515 74.455 ;
        RECT 234.015 73.255 234.615 73.395 ;
        RECT 233.495 72.435 233.755 72.755 ;
        RECT 233.555 70.715 233.695 72.435 ;
        RECT 234.475 70.910 234.615 73.255 ;
        RECT 233.495 70.395 233.755 70.715 ;
        RECT 234.405 70.540 234.685 70.910 ;
        RECT 234.475 69.355 234.615 70.540 ;
        RECT 235.335 70.055 235.595 70.375 ;
        RECT 235.395 69.355 235.535 70.055 ;
        RECT 234.415 69.035 234.675 69.355 ;
        RECT 235.335 69.035 235.595 69.355 ;
        RECT 233.035 68.695 233.295 69.015 ;
        RECT 236.315 63.915 236.455 74.135 ;
        RECT 236.775 72.755 236.915 75.835 ;
        RECT 237.235 75.475 237.375 104.055 ;
        RECT 238.155 102.675 238.295 104.055 ;
        RECT 238.095 102.355 238.355 102.675 ;
        RECT 238.085 83.460 238.365 83.830 ;
        RECT 237.175 75.155 237.435 75.475 ;
        RECT 237.635 74.815 237.895 75.135 ;
        RECT 237.695 73.435 237.835 74.815 ;
        RECT 237.635 73.115 237.895 73.435 ;
        RECT 237.175 72.775 237.435 73.095 ;
        RECT 236.715 72.435 236.975 72.755 ;
        RECT 237.235 71.735 237.375 72.775 ;
        RECT 237.635 72.665 237.895 72.755 ;
        RECT 238.155 72.665 238.295 83.460 ;
        RECT 238.615 80.575 238.755 104.735 ;
        RECT 239.995 102.675 240.135 109.225 ;
        RECT 242.295 107.095 242.435 109.225 ;
        RECT 242.695 109.155 242.955 109.475 ;
        RECT 244.525 109.225 244.805 130.460 ;
        RECT 246.825 109.225 247.105 131.040 ;
        RECT 249.125 109.225 249.405 131.620 ;
        RECT 251.425 109.225 251.705 132.200 ;
        RECT 253.725 109.225 254.005 132.780 ;
        RECT 256.025 109.225 256.305 133.360 ;
        RECT 258.325 109.225 258.605 133.940 ;
        RECT 258.855 109.415 259.915 109.555 ;
        RECT 242.235 106.775 242.495 107.095 ;
        RECT 242.755 106.075 242.895 109.155 ;
        RECT 242.695 105.755 242.955 106.075 ;
        RECT 244.595 104.625 244.735 109.225 ;
        RECT 245.455 108.815 245.715 109.135 ;
        RECT 244.995 107.115 245.255 107.435 ;
        RECT 245.055 105.395 245.195 107.115 ;
        RECT 244.995 105.075 245.255 105.395 ;
        RECT 244.995 104.625 245.255 104.715 ;
        RECT 244.595 104.485 245.255 104.625 ;
        RECT 244.995 104.395 245.255 104.485 ;
        RECT 241.315 103.035 241.575 103.355 ;
        RECT 239.935 102.355 240.195 102.675 ;
        RECT 239.935 101.335 240.195 101.655 ;
        RECT 239.995 99.955 240.135 101.335 ;
        RECT 241.375 100.295 241.515 103.035 ;
        RECT 241.315 99.975 241.575 100.295 ;
        RECT 239.935 99.635 240.195 99.955 ;
        RECT 244.075 99.295 244.335 99.615 ;
        RECT 243.155 97.430 243.415 97.575 ;
        RECT 243.145 97.060 243.425 97.430 ;
        RECT 241.315 96.575 241.575 96.895 ;
        RECT 241.775 96.575 242.035 96.895 ;
        RECT 241.375 95.195 241.515 96.575 ;
        RECT 241.315 94.875 241.575 95.195 ;
        RECT 239.475 94.195 239.735 94.515 ;
        RECT 239.015 88.415 239.275 88.735 ;
        RECT 238.555 80.255 238.815 80.575 ;
        RECT 237.635 72.525 238.295 72.665 ;
        RECT 237.635 72.435 237.895 72.525 ;
        RECT 237.175 71.415 237.435 71.735 ;
        RECT 236.715 64.275 236.975 64.595 ;
        RECT 236.255 63.595 236.515 63.915 ;
        RECT 236.775 62.215 236.915 64.275 ;
        RECT 236.715 61.895 236.975 62.215 ;
        RECT 225.215 61.215 225.475 61.535 ;
        RECT 225.275 50.315 225.415 61.215 ;
        RECT 225.675 58.155 225.935 58.475 ;
        RECT 225.735 55.415 225.875 58.155 ;
        RECT 226.195 57.310 226.335 61.815 ;
        RECT 231.655 61.555 231.915 61.875 ;
        RECT 234.875 61.555 235.135 61.875 ;
        RECT 230.275 60.535 230.535 60.855 ;
        RECT 233.955 60.535 234.215 60.855 ;
        RECT 227.515 58.835 227.775 59.155 ;
        RECT 226.125 56.940 226.405 57.310 ;
        RECT 227.575 56.095 227.715 58.835 ;
        RECT 228.435 58.495 228.695 58.815 ;
        RECT 228.495 56.435 228.635 58.495 ;
        RECT 229.815 57.815 230.075 58.135 ;
        RECT 228.435 56.115 228.695 56.435 ;
        RECT 227.515 55.775 227.775 56.095 ;
        RECT 226.135 55.435 226.395 55.755 ;
        RECT 225.675 55.095 225.935 55.415 ;
        RECT 225.675 52.605 225.935 52.695 ;
        RECT 226.195 52.605 226.335 55.435 ;
        RECT 229.875 54.395 230.015 57.815 ;
        RECT 230.335 56.775 230.475 60.535 ;
        RECT 232.575 58.495 232.835 58.815 ;
        RECT 232.115 58.155 232.375 58.475 ;
        RECT 230.275 56.455 230.535 56.775 ;
        RECT 231.655 55.095 231.915 55.415 ;
        RECT 231.715 54.590 231.855 55.095 ;
        RECT 229.815 54.075 230.075 54.395 ;
        RECT 231.645 54.220 231.925 54.590 ;
        RECT 227.975 53.735 228.235 54.055 ;
        RECT 225.675 52.465 226.335 52.605 ;
        RECT 225.675 52.375 225.935 52.465 ;
        RECT 225.215 49.995 225.475 50.315 ;
        RECT 225.275 45.215 225.415 49.995 ;
        RECT 226.195 47.935 226.335 52.465 ;
        RECT 226.135 47.615 226.395 47.935 ;
        RECT 226.195 45.895 226.335 47.615 ;
        RECT 227.515 47.275 227.775 47.595 ;
        RECT 226.595 46.935 226.855 47.255 ;
        RECT 226.135 45.575 226.395 45.895 ;
        RECT 225.215 44.895 225.475 45.215 ;
        RECT 226.135 44.215 226.395 44.535 ;
        RECT 226.195 42.835 226.335 44.215 ;
        RECT 226.655 43.515 226.795 46.935 ;
        RECT 227.045 45.380 227.325 45.750 ;
        RECT 227.055 45.235 227.315 45.380 ;
        RECT 227.575 43.515 227.715 47.275 ;
        RECT 228.035 45.555 228.175 53.735 ;
        RECT 229.815 53.395 230.075 53.715 ;
        RECT 230.275 53.395 230.535 53.715 ;
        RECT 229.875 45.555 230.015 53.395 ;
        RECT 230.335 50.995 230.475 53.395 ;
        RECT 232.175 53.035 232.315 58.155 ;
        RECT 232.635 53.715 232.775 58.495 ;
        RECT 234.015 58.475 234.155 60.535 ;
        RECT 233.955 58.155 234.215 58.475 ;
        RECT 234.935 55.755 235.075 61.555 ;
        RECT 238.615 61.535 238.755 80.255 ;
        RECT 239.075 74.455 239.215 88.415 ;
        RECT 239.535 83.635 239.675 94.195 ;
        RECT 241.835 90.775 241.975 96.575 ;
        RECT 242.685 94.340 242.965 94.710 ;
        RECT 244.135 94.515 244.275 99.295 ;
        RECT 244.995 98.675 245.255 98.935 ;
        RECT 245.515 98.675 245.655 108.815 ;
        RECT 246.375 108.475 246.635 108.795 ;
        RECT 246.435 104.965 246.575 108.475 ;
        RECT 246.895 105.735 247.035 109.225 ;
        RECT 248.215 107.115 248.475 107.435 ;
        RECT 246.835 105.415 247.095 105.735 ;
        RECT 246.435 104.825 247.035 104.965 ;
        RECT 246.375 103.265 246.635 103.355 ;
        RECT 245.975 103.125 246.635 103.265 ;
        RECT 245.975 101.655 246.115 103.125 ;
        RECT 246.375 103.035 246.635 103.125 ;
        RECT 246.375 102.015 246.635 102.335 ;
        RECT 245.915 101.335 246.175 101.655 ;
        RECT 244.995 98.615 245.655 98.675 ;
        RECT 245.055 98.535 245.655 98.615 ;
        RECT 245.515 96.895 245.655 98.535 ;
        RECT 245.455 96.575 245.715 96.895 ;
        RECT 244.535 96.235 244.795 96.555 ;
        RECT 244.595 95.195 244.735 96.235 ;
        RECT 244.535 94.875 244.795 95.195 ;
        RECT 243.155 94.425 243.415 94.515 ;
        RECT 242.695 94.195 242.955 94.340 ;
        RECT 243.155 94.285 243.815 94.425 ;
        RECT 243.155 94.195 243.415 94.285 ;
        RECT 243.155 93.175 243.415 93.495 ;
        RECT 243.215 92.135 243.355 93.175 ;
        RECT 243.155 91.815 243.415 92.135 ;
        RECT 242.235 91.135 242.495 91.455 ;
        RECT 242.695 91.310 242.955 91.455 ;
        RECT 241.775 90.455 242.035 90.775 ;
        RECT 240.855 85.015 241.115 85.335 ;
        RECT 240.915 83.975 241.055 85.015 ;
        RECT 241.835 84.315 241.975 90.455 ;
        RECT 241.775 83.995 242.035 84.315 ;
        RECT 240.855 83.655 241.115 83.975 ;
        RECT 239.475 83.315 239.735 83.635 ;
        RECT 239.535 80.915 239.675 83.315 ;
        RECT 241.775 82.635 242.035 82.955 ;
        RECT 241.835 82.470 241.975 82.635 ;
        RECT 241.765 82.100 242.045 82.470 ;
        RECT 239.935 80.935 240.195 81.255 ;
        RECT 239.475 80.595 239.735 80.915 ;
        RECT 239.995 80.575 240.135 80.935 ;
        RECT 241.765 80.740 242.045 81.110 ;
        RECT 241.835 80.575 241.975 80.740 ;
        RECT 239.935 80.255 240.195 80.575 ;
        RECT 240.395 80.255 240.655 80.575 ;
        RECT 241.775 80.255 242.035 80.575 ;
        RECT 242.295 80.315 242.435 91.135 ;
        RECT 242.685 90.940 242.965 91.310 ;
        RECT 243.675 89.755 243.815 94.285 ;
        RECT 244.075 94.195 244.335 94.515 ;
        RECT 244.535 94.195 244.795 94.515 ;
        RECT 245.455 94.195 245.715 94.515 ;
        RECT 243.615 89.435 243.875 89.755 ;
        RECT 244.135 89.075 244.275 94.195 ;
        RECT 244.595 92.475 244.735 94.195 ;
        RECT 245.515 93.915 245.655 94.195 ;
        RECT 245.055 93.775 245.655 93.915 ;
        RECT 245.055 93.495 245.195 93.775 ;
        RECT 244.995 93.175 245.255 93.495 ;
        RECT 244.535 92.155 244.795 92.475 ;
        RECT 245.975 91.310 246.115 101.335 ;
        RECT 246.435 100.295 246.575 102.015 ;
        RECT 246.895 101.655 247.035 104.825 ;
        RECT 247.295 104.230 247.555 104.375 ;
        RECT 247.285 103.860 247.565 104.230 ;
        RECT 247.755 104.055 248.015 104.375 ;
        RECT 247.815 102.675 247.955 104.055 ;
        RECT 247.755 102.355 248.015 102.675 ;
        RECT 246.835 101.335 247.095 101.655 ;
        RECT 246.375 99.975 246.635 100.295 ;
        RECT 247.755 99.635 248.015 99.955 ;
        RECT 247.815 98.675 247.955 99.635 ;
        RECT 248.275 99.615 248.415 107.115 ;
        RECT 248.675 101.335 248.935 101.655 ;
        RECT 248.215 99.295 248.475 99.615 ;
        RECT 247.815 98.535 248.415 98.675 ;
        RECT 248.275 96.895 248.415 98.535 ;
        RECT 248.735 97.315 248.875 101.335 ;
        RECT 249.195 99.275 249.335 109.225 ;
        RECT 251.495 106.075 251.635 109.225 ;
        RECT 252.815 108.475 253.075 108.795 ;
        RECT 252.355 108.135 252.615 108.455 ;
        RECT 251.435 105.755 251.695 106.075 ;
        RECT 249.595 104.735 249.855 105.055 ;
        RECT 250.975 104.735 251.235 105.055 ;
        RECT 249.655 102.675 249.795 104.735 ;
        RECT 251.035 103.355 251.175 104.735 ;
        RECT 250.975 103.035 251.235 103.355 ;
        RECT 249.595 102.355 249.855 102.675 ;
        RECT 249.655 99.615 249.795 102.355 ;
        RECT 250.055 102.015 250.315 102.335 ;
        RECT 250.115 101.655 250.255 102.015 ;
        RECT 250.055 101.335 250.315 101.655 ;
        RECT 250.515 100.315 250.775 100.635 ;
        RECT 250.575 99.955 250.715 100.315 ;
        RECT 250.055 99.635 250.315 99.955 ;
        RECT 250.515 99.635 250.775 99.955 ;
        RECT 250.975 99.635 251.235 99.955 ;
        RECT 249.595 99.295 249.855 99.615 ;
        RECT 250.115 99.470 250.255 99.635 ;
        RECT 249.135 98.955 249.395 99.275 ;
        RECT 250.045 99.100 250.325 99.470 ;
        RECT 248.735 97.175 249.795 97.315 ;
        RECT 246.375 96.575 246.635 96.895 ;
        RECT 248.215 96.575 248.475 96.895 ;
        RECT 246.435 92.475 246.575 96.575 ;
        RECT 247.755 96.465 248.015 96.555 ;
        RECT 246.895 96.325 248.015 96.465 ;
        RECT 246.375 92.155 246.635 92.475 ;
        RECT 245.455 90.795 245.715 91.115 ;
        RECT 245.905 90.940 246.185 91.310 ;
        RECT 246.895 91.115 247.035 96.325 ;
        RECT 247.755 96.235 248.015 96.325 ;
        RECT 247.745 95.700 248.025 96.070 ;
        RECT 247.815 94.515 247.955 95.700 ;
        RECT 248.215 94.875 248.475 95.195 ;
        RECT 247.755 94.195 248.015 94.515 ;
        RECT 247.295 93.855 247.555 94.175 ;
        RECT 247.355 91.795 247.495 93.855 ;
        RECT 247.755 93.175 248.015 93.495 ;
        RECT 247.295 91.475 247.555 91.795 ;
        RECT 246.835 90.795 247.095 91.115 ;
        RECT 247.285 90.940 247.565 91.310 ;
        RECT 247.295 90.795 247.555 90.940 ;
        RECT 242.695 88.755 242.955 89.075 ;
        RECT 244.075 88.755 244.335 89.075 ;
        RECT 244.535 88.755 244.795 89.075 ;
        RECT 242.755 86.695 242.895 88.755 ;
        RECT 243.155 88.475 243.415 88.735 ;
        RECT 244.595 88.475 244.735 88.755 ;
        RECT 243.155 88.415 244.735 88.475 ;
        RECT 243.215 88.335 244.735 88.415 ;
        RECT 244.525 87.540 244.805 87.910 ;
        RECT 242.695 86.375 242.955 86.695 ;
        RECT 244.075 86.375 244.335 86.695 ;
        RECT 244.135 86.015 244.275 86.375 ;
        RECT 242.695 85.695 242.955 86.015 ;
        RECT 243.155 85.695 243.415 86.015 ;
        RECT 244.075 85.925 244.335 86.015 ;
        RECT 243.675 85.785 244.335 85.925 ;
        RECT 242.755 83.635 242.895 85.695 ;
        RECT 242.695 83.315 242.955 83.635 ;
        RECT 239.995 78.875 240.135 80.255 ;
        RECT 239.935 78.555 240.195 78.875 ;
        RECT 239.015 74.135 239.275 74.455 ;
        RECT 239.075 64.935 239.215 74.135 ;
        RECT 240.455 68.190 240.595 80.255 ;
        RECT 242.295 80.175 242.895 80.315 ;
        RECT 241.315 79.575 241.575 79.895 ;
        RECT 241.775 79.575 242.035 79.895 ;
        RECT 242.235 79.575 242.495 79.895 ;
        RECT 241.375 77.765 241.515 79.575 ;
        RECT 241.835 78.535 241.975 79.575 ;
        RECT 241.775 78.215 242.035 78.535 ;
        RECT 242.295 77.855 242.435 79.575 ;
        RECT 241.375 77.625 241.975 77.765 ;
        RECT 241.315 75.835 241.575 76.155 ;
        RECT 241.375 73.435 241.515 75.835 ;
        RECT 241.315 73.115 241.575 73.435 ;
        RECT 241.315 72.435 241.575 72.755 ;
        RECT 241.375 70.715 241.515 72.435 ;
        RECT 241.315 70.395 241.575 70.715 ;
        RECT 241.835 69.695 241.975 77.625 ;
        RECT 242.235 77.535 242.495 77.855 ;
        RECT 242.755 73.395 242.895 80.175 ;
        RECT 242.295 73.255 242.895 73.395 ;
        RECT 242.295 72.755 242.435 73.255 ;
        RECT 242.235 72.435 242.495 72.755 ;
        RECT 241.775 69.375 242.035 69.695 ;
        RECT 240.855 68.695 241.115 69.015 ;
        RECT 241.315 68.695 241.575 69.015 ;
        RECT 242.295 68.755 242.435 72.435 ;
        RECT 242.685 69.860 242.965 70.230 ;
        RECT 242.755 69.355 242.895 69.860 ;
        RECT 242.695 69.035 242.955 69.355 ;
        RECT 240.385 67.820 240.665 68.190 ;
        RECT 240.455 67.315 240.595 67.820 ;
        RECT 240.915 67.315 241.055 68.695 ;
        RECT 240.395 66.995 240.655 67.315 ;
        RECT 240.855 66.995 241.115 67.315 ;
        RECT 241.375 65.275 241.515 68.695 ;
        RECT 242.295 68.615 242.895 68.755 ;
        RECT 242.755 66.635 242.895 68.615 ;
        RECT 242.235 66.315 242.495 66.635 ;
        RECT 242.695 66.315 242.955 66.635 ;
        RECT 241.315 64.955 241.575 65.275 ;
        RECT 239.015 64.615 239.275 64.935 ;
        RECT 238.555 61.215 238.815 61.535 ;
        RECT 241.315 61.215 241.575 61.535 ;
        RECT 241.375 59.495 241.515 61.215 ;
        RECT 241.315 59.175 241.575 59.495 ;
        RECT 236.715 58.155 236.975 58.475 ;
        RECT 236.775 56.775 236.915 58.155 ;
        RECT 237.175 57.815 237.435 58.135 ;
        RECT 236.715 56.455 236.975 56.775 ;
        RECT 234.875 55.435 235.135 55.755 ;
        RECT 233.035 55.095 233.295 55.415 ;
        RECT 233.095 54.055 233.235 55.095 ;
        RECT 234.405 54.900 234.685 55.270 ;
        RECT 233.485 54.220 233.765 54.590 ;
        RECT 234.475 54.395 234.615 54.900 ;
        RECT 233.555 54.055 233.695 54.220 ;
        RECT 234.415 54.075 234.675 54.395 ;
        RECT 233.035 53.735 233.295 54.055 ;
        RECT 233.495 53.735 233.755 54.055 ;
        RECT 232.575 53.395 232.835 53.715 ;
        RECT 236.255 53.055 236.515 53.375 ;
        RECT 232.115 52.715 232.375 53.035 ;
        RECT 233.035 52.715 233.295 53.035 ;
        RECT 235.335 52.715 235.595 53.035 ;
        RECT 230.275 50.675 230.535 50.995 ;
        RECT 230.335 48.275 230.475 50.675 ;
        RECT 231.655 49.655 231.915 49.975 ;
        RECT 230.275 47.955 230.535 48.275 ;
        RECT 227.975 45.235 228.235 45.555 ;
        RECT 229.815 45.235 230.075 45.555 ;
        RECT 231.715 45.215 231.855 49.655 ;
        RECT 233.095 47.110 233.235 52.715 ;
        RECT 233.025 46.740 233.305 47.110 ;
        RECT 233.095 46.235 233.235 46.740 ;
        RECT 233.035 45.915 233.295 46.235 ;
        RECT 228.435 44.895 228.695 45.215 ;
        RECT 230.275 44.895 230.535 45.215 ;
        RECT 231.655 44.895 231.915 45.215 ;
        RECT 228.495 43.515 228.635 44.895 ;
        RECT 226.595 43.195 226.855 43.515 ;
        RECT 227.515 43.195 227.775 43.515 ;
        RECT 228.435 43.195 228.695 43.515 ;
        RECT 226.135 42.515 226.395 42.835 ;
        RECT 230.335 42.495 230.475 44.895 ;
        RECT 235.395 42.835 235.535 52.715 ;
        RECT 236.315 50.995 236.455 53.055 ;
        RECT 236.255 50.675 236.515 50.995 ;
        RECT 236.315 45.750 236.455 50.675 ;
        RECT 236.775 49.715 236.915 56.455 ;
        RECT 237.235 53.375 237.375 57.815 ;
        RECT 239.475 56.115 239.735 56.435 ;
        RECT 239.015 55.095 239.275 55.415 ;
        RECT 239.075 53.375 239.215 55.095 ;
        RECT 237.175 53.055 237.435 53.375 ;
        RECT 238.095 53.285 238.355 53.375 ;
        RECT 237.695 53.145 238.355 53.285 ;
        RECT 236.775 49.575 237.375 49.715 ;
        RECT 236.715 48.635 236.975 48.955 ;
        RECT 236.245 45.380 236.525 45.750 ;
        RECT 236.775 42.835 236.915 48.635 ;
        RECT 235.335 42.515 235.595 42.835 ;
        RECT 236.715 42.515 236.975 42.835 ;
        RECT 227.055 42.175 227.315 42.495 ;
        RECT 230.275 42.175 230.535 42.495 ;
        RECT 226.135 41.495 226.395 41.815 ;
        RECT 219.695 40.475 219.955 40.795 ;
        RECT 224.755 40.475 225.015 40.795 ;
        RECT 217.855 40.135 218.115 40.455 ;
        RECT 217.915 39.515 218.055 40.135 ;
        RECT 226.195 39.775 226.335 41.495 ;
        RECT 227.115 40.115 227.255 42.175 ;
        RECT 227.975 40.475 228.235 40.795 ;
        RECT 227.055 39.795 227.315 40.115 ;
        RECT 216.995 39.375 218.055 39.515 ;
        RECT 221.535 39.455 221.795 39.775 ;
        RECT 226.135 39.455 226.395 39.775 ;
        RECT 214.635 38.775 214.895 39.095 ;
        RECT 216.475 38.775 216.735 39.095 ;
        RECT 216.535 37.055 216.675 38.775 ;
        RECT 209.115 36.735 209.375 37.055 ;
        RECT 216.475 36.735 216.735 37.055 ;
        RECT 208.655 36.395 208.915 36.715 ;
        RECT 209.175 35.355 209.315 36.735 ;
        RECT 216.015 36.055 216.275 36.375 ;
        RECT 216.075 35.355 216.215 36.055 ;
        RECT 209.115 35.035 209.375 35.355 ;
        RECT 216.015 35.035 216.275 35.355 ;
        RECT 208.195 34.695 208.455 35.015 ;
        RECT 205.895 32.315 206.155 32.635 ;
        RECT 204.975 30.955 205.235 31.275 ;
        RECT 202.675 30.615 202.935 30.935 ;
        RECT 199.915 29.595 200.175 29.915 ;
        RECT 202.735 29.575 202.875 30.615 ;
        RECT 205.035 29.915 205.175 30.955 ;
        RECT 204.975 29.595 205.235 29.915 ;
        RECT 199.455 29.255 199.715 29.575 ;
        RECT 202.675 29.255 202.935 29.575 ;
        RECT 205.955 29.235 206.095 32.315 ;
        RECT 208.255 31.615 208.395 34.695 ;
        RECT 210.955 34.015 211.215 34.335 ;
        RECT 211.015 32.635 211.155 34.015 ;
        RECT 213.255 33.335 213.515 33.655 ;
        RECT 213.315 32.635 213.455 33.335 ;
        RECT 210.955 32.315 211.215 32.635 ;
        RECT 213.255 32.315 213.515 32.635 ;
        RECT 216.075 31.615 216.215 35.035 ;
        RECT 216.995 35.015 217.135 39.375 ;
        RECT 217.645 38.240 219.185 38.610 ;
        RECT 221.595 38.075 221.735 39.455 ;
        RECT 221.535 37.755 221.795 38.075 ;
        RECT 227.115 37.055 227.255 39.795 ;
        RECT 227.515 39.115 227.775 39.435 ;
        RECT 227.575 37.395 227.715 39.115 ;
        RECT 228.035 37.395 228.175 40.475 ;
        RECT 235.335 40.135 235.595 40.455 ;
        RECT 234.875 39.795 235.135 40.115 ;
        RECT 231.195 39.455 231.455 39.775 ;
        RECT 230.735 37.985 230.995 38.075 ;
        RECT 231.255 37.985 231.395 39.455 ;
        RECT 231.655 38.775 231.915 39.095 ;
        RECT 232.115 38.775 232.375 39.095 ;
        RECT 230.735 37.845 231.395 37.985 ;
        RECT 230.735 37.755 230.995 37.845 ;
        RECT 227.515 37.075 227.775 37.395 ;
        RECT 227.975 37.075 228.235 37.395 ;
        RECT 227.055 36.735 227.315 37.055 ;
        RECT 225.675 36.395 225.935 36.715 ;
        RECT 220.945 35.520 222.485 35.890 ;
        RECT 225.735 35.355 225.875 36.395 ;
        RECT 226.135 36.055 226.395 36.375 ;
        RECT 225.675 35.035 225.935 35.355 ;
        RECT 216.935 34.695 217.195 35.015 ;
        RECT 220.615 34.015 220.875 34.335 ;
        RECT 225.675 34.015 225.935 34.335 ;
        RECT 217.645 32.800 219.185 33.170 ;
        RECT 220.675 32.635 220.815 34.015 ;
        RECT 225.735 32.635 225.875 34.015 ;
        RECT 226.195 32.635 226.335 36.055 ;
        RECT 227.115 34.335 227.255 36.735 ;
        RECT 231.255 36.715 231.395 37.845 ;
        RECT 231.715 36.715 231.855 38.775 ;
        RECT 231.195 36.395 231.455 36.715 ;
        RECT 231.655 36.395 231.915 36.715 ;
        RECT 228.435 36.055 228.695 36.375 ;
        RECT 227.055 34.015 227.315 34.335 ;
        RECT 220.615 32.315 220.875 32.635 ;
        RECT 225.675 32.315 225.935 32.635 ;
        RECT 226.135 32.315 226.395 32.635 ;
        RECT 227.115 31.615 227.255 34.015 ;
        RECT 228.495 33.655 228.635 36.055 ;
        RECT 232.175 35.015 232.315 38.775 ;
        RECT 234.935 35.355 235.075 39.795 ;
        RECT 234.415 35.035 234.675 35.355 ;
        RECT 234.875 35.035 235.135 35.355 ;
        RECT 228.895 34.695 229.155 35.015 ;
        RECT 232.115 34.695 232.375 35.015 ;
        RECT 228.435 33.335 228.695 33.655 ;
        RECT 228.495 31.955 228.635 33.335 ;
        RECT 228.955 31.955 229.095 34.695 ;
        RECT 234.475 32.635 234.615 35.035 ;
        RECT 234.415 32.315 234.675 32.635 ;
        RECT 228.435 31.635 228.695 31.955 ;
        RECT 228.895 31.635 229.155 31.955 ;
        RECT 208.195 31.295 208.455 31.615 ;
        RECT 216.015 31.295 216.275 31.615 ;
        RECT 227.055 31.295 227.315 31.615 ;
        RECT 220.945 30.080 222.485 30.450 ;
        RECT 234.935 29.235 235.075 35.035 ;
        RECT 235.395 31.615 235.535 40.135 ;
        RECT 235.795 39.455 236.055 39.775 ;
        RECT 236.715 39.455 236.975 39.775 ;
        RECT 235.335 31.295 235.595 31.615 ;
        RECT 235.855 30.935 235.995 39.455 ;
        RECT 236.775 36.375 236.915 39.455 ;
        RECT 237.235 37.735 237.375 49.575 ;
        RECT 237.695 44.535 237.835 53.145 ;
        RECT 238.095 53.055 238.355 53.145 ;
        RECT 239.015 53.055 239.275 53.375 ;
        RECT 239.015 50.335 239.275 50.655 ;
        RECT 238.095 47.275 238.355 47.595 ;
        RECT 237.635 44.215 237.895 44.535 ;
        RECT 238.155 42.155 238.295 47.275 ;
        RECT 238.555 46.935 238.815 47.255 ;
        RECT 238.095 42.065 238.355 42.155 ;
        RECT 237.695 41.925 238.355 42.065 ;
        RECT 237.175 37.415 237.435 37.735 ;
        RECT 236.715 36.055 236.975 36.375 ;
        RECT 237.695 35.015 237.835 41.925 ;
        RECT 238.095 41.835 238.355 41.925 ;
        RECT 238.615 40.115 238.755 46.935 ;
        RECT 239.075 43.515 239.215 50.335 ;
        RECT 239.015 43.195 239.275 43.515 ;
        RECT 239.535 41.815 239.675 56.115 ;
        RECT 242.295 53.715 242.435 66.315 ;
        RECT 242.695 63.935 242.955 64.255 ;
        RECT 242.755 62.555 242.895 63.935 ;
        RECT 242.695 62.235 242.955 62.555 ;
        RECT 243.215 59.595 243.355 85.695 ;
        RECT 243.675 81.595 243.815 85.785 ;
        RECT 244.075 85.695 244.335 85.785 ;
        RECT 244.075 85.015 244.335 85.335 ;
        RECT 244.135 83.295 244.275 85.015 ;
        RECT 244.075 82.975 244.335 83.295 ;
        RECT 243.615 81.275 243.875 81.595 ;
        RECT 244.135 80.575 244.275 82.975 ;
        RECT 244.595 80.575 244.735 87.540 ;
        RECT 244.995 83.830 245.255 83.975 ;
        RECT 244.985 83.460 245.265 83.830 ;
        RECT 244.995 82.975 245.255 83.295 ;
        RECT 244.075 80.255 244.335 80.575 ;
        RECT 244.535 80.255 244.795 80.575 ;
        RECT 244.535 79.575 244.795 79.895 ;
        RECT 244.595 77.175 244.735 79.575 ;
        RECT 243.615 76.855 243.875 77.175 ;
        RECT 244.535 76.855 244.795 77.175 ;
        RECT 243.675 72.665 243.815 76.855 ;
        RECT 245.055 73.435 245.195 82.975 ;
        RECT 244.995 73.115 245.255 73.435 ;
        RECT 244.070 72.665 244.330 72.755 ;
        RECT 243.675 72.525 244.330 72.665 ;
        RECT 243.675 65.470 243.815 72.525 ;
        RECT 244.070 72.435 244.330 72.525 ;
        RECT 245.515 70.795 245.655 90.795 ;
        RECT 246.895 89.755 247.035 90.795 ;
        RECT 246.835 89.435 247.095 89.755 ;
        RECT 245.915 86.715 246.175 87.035 ;
        RECT 245.975 84.315 246.115 86.715 ;
        RECT 246.895 85.335 247.035 89.435 ;
        RECT 247.815 89.075 247.955 93.175 ;
        RECT 248.275 91.990 248.415 94.875 ;
        RECT 249.135 94.195 249.395 94.515 ;
        RECT 248.205 91.620 248.485 91.990 ;
        RECT 248.215 91.135 248.475 91.455 ;
        RECT 247.755 88.755 248.015 89.075 ;
        RECT 246.835 85.015 247.095 85.335 ;
        RECT 248.275 84.315 248.415 91.135 ;
        RECT 249.195 90.775 249.335 94.195 ;
        RECT 249.135 90.455 249.395 90.775 ;
        RECT 249.195 85.335 249.335 90.455 ;
        RECT 249.655 89.755 249.795 97.175 ;
        RECT 250.115 96.635 250.255 99.100 ;
        RECT 251.035 98.790 251.175 99.635 ;
        RECT 250.965 98.420 251.245 98.790 ;
        RECT 250.115 96.495 252.095 96.635 ;
        RECT 251.435 95.895 251.695 96.215 ;
        RECT 251.495 94.515 251.635 95.895 ;
        RECT 250.055 94.195 250.315 94.515 ;
        RECT 250.975 94.195 251.235 94.515 ;
        RECT 251.435 94.195 251.695 94.515 ;
        RECT 250.115 90.775 250.255 94.195 ;
        RECT 251.035 91.990 251.175 94.195 ;
        RECT 250.965 91.620 251.245 91.990 ;
        RECT 250.055 90.455 250.315 90.775 ;
        RECT 249.595 89.435 249.855 89.755 ;
        RECT 250.115 86.945 250.255 90.455 ;
        RECT 251.035 89.415 251.175 91.620 ;
        RECT 250.975 89.095 251.235 89.415 ;
        RECT 250.515 88.755 250.775 89.075 ;
        RECT 250.575 87.035 250.715 88.755 ;
        RECT 249.655 86.805 250.255 86.945 ;
        RECT 248.675 85.015 248.935 85.335 ;
        RECT 249.135 85.015 249.395 85.335 ;
        RECT 245.915 83.995 246.175 84.315 ;
        RECT 246.375 83.995 246.635 84.315 ;
        RECT 248.215 83.995 248.475 84.315 ;
        RECT 245.915 83.545 246.175 83.635 ;
        RECT 246.435 83.545 246.575 83.995 ;
        RECT 248.735 83.975 248.875 85.015 ;
        RECT 248.675 83.655 248.935 83.975 ;
        RECT 245.915 83.405 246.575 83.545 ;
        RECT 245.915 83.315 246.175 83.405 ;
        RECT 246.835 83.315 247.095 83.635 ;
        RECT 245.975 80.575 246.115 83.315 ;
        RECT 246.375 82.865 246.635 82.955 ;
        RECT 246.895 82.865 247.035 83.315 ;
        RECT 249.195 82.955 249.335 85.015 ;
        RECT 246.375 82.725 247.035 82.865 ;
        RECT 246.375 82.635 246.635 82.725 ;
        RECT 249.135 82.635 249.395 82.955 ;
        RECT 247.295 82.295 247.555 82.615 ;
        RECT 247.355 81.790 247.495 82.295 ;
        RECT 247.285 81.420 247.565 81.790 ;
        RECT 249.195 80.575 249.335 82.635 ;
        RECT 249.655 81.110 249.795 86.805 ;
        RECT 250.515 86.715 250.775 87.035 ;
        RECT 250.055 86.035 250.315 86.355 ;
        RECT 250.115 83.635 250.255 86.035 ;
        RECT 250.055 83.315 250.315 83.635 ;
        RECT 249.585 80.740 249.865 81.110 ;
        RECT 245.915 80.255 246.175 80.575 ;
        RECT 246.835 80.255 247.095 80.575 ;
        RECT 248.675 80.430 248.935 80.575 ;
        RECT 246.895 79.750 247.035 80.255 ;
        RECT 247.295 79.915 247.555 80.235 ;
        RECT 248.665 80.060 248.945 80.430 ;
        RECT 249.135 80.255 249.395 80.575 ;
        RECT 250.975 80.255 251.235 80.575 ;
        RECT 246.825 79.380 247.105 79.750 ;
        RECT 245.915 74.135 246.175 74.455 ;
        RECT 245.975 73.435 246.115 74.135 ;
        RECT 245.915 73.115 246.175 73.435 ;
        RECT 245.975 72.755 246.115 73.115 ;
        RECT 247.355 73.005 247.495 79.915 ;
        RECT 248.215 79.575 248.475 79.895 ;
        RECT 249.135 79.575 249.395 79.895 ;
        RECT 249.595 79.750 249.855 79.895 ;
        RECT 248.275 79.070 248.415 79.575 ;
        RECT 248.205 78.700 248.485 79.070 ;
        RECT 249.195 78.195 249.335 79.575 ;
        RECT 249.585 79.380 249.865 79.750 ;
        RECT 249.135 77.875 249.395 78.195 ;
        RECT 246.895 72.865 247.495 73.005 ;
        RECT 245.915 72.435 246.175 72.755 ;
        RECT 245.055 70.655 245.655 70.795 ;
        RECT 245.055 69.355 245.195 70.655 ;
        RECT 245.455 70.055 245.715 70.375 ;
        RECT 246.895 70.230 247.035 72.865 ;
        RECT 247.295 71.415 247.555 71.735 ;
        RECT 244.535 69.035 244.795 69.355 ;
        RECT 244.995 69.035 245.255 69.355 ;
        RECT 244.075 66.995 244.335 67.315 ;
        RECT 243.605 65.100 243.885 65.470 ;
        RECT 244.135 64.935 244.275 66.995 ;
        RECT 244.075 64.615 244.335 64.935 ;
        RECT 244.135 62.215 244.275 64.615 ;
        RECT 244.595 63.485 244.735 69.035 ;
        RECT 245.055 67.315 245.195 69.035 ;
        RECT 244.995 66.995 245.255 67.315 ;
        RECT 244.995 66.315 245.255 66.635 ;
        RECT 245.055 64.255 245.195 66.315 ;
        RECT 245.515 66.295 245.655 70.055 ;
        RECT 246.825 69.860 247.105 70.230 ;
        RECT 247.355 69.695 247.495 71.415 ;
        RECT 245.915 69.375 246.175 69.695 ;
        RECT 247.295 69.375 247.555 69.695 ;
        RECT 247.755 69.550 248.015 69.695 ;
        RECT 251.035 69.550 251.175 80.255 ;
        RECT 251.955 73.095 252.095 96.495 ;
        RECT 252.415 78.195 252.555 108.135 ;
        RECT 252.875 100.295 253.015 108.475 ;
        RECT 253.275 107.455 253.535 107.775 ;
        RECT 252.815 99.975 253.075 100.295 ;
        RECT 253.335 100.205 253.475 107.455 ;
        RECT 253.795 105.735 253.935 109.225 ;
        RECT 256.095 107.095 256.235 109.225 ;
        RECT 258.395 108.875 258.535 109.225 ;
        RECT 258.855 108.875 258.995 109.415 ;
        RECT 258.395 108.735 258.995 108.875 ;
        RECT 256.495 107.795 256.755 108.115 ;
        RECT 255.575 106.775 255.835 107.095 ;
        RECT 256.035 106.775 256.295 107.095 ;
        RECT 253.735 105.415 253.995 105.735 ;
        RECT 255.115 104.735 255.375 105.055 ;
        RECT 254.655 104.055 254.915 104.375 ;
        RECT 254.195 101.675 254.455 101.995 ;
        RECT 254.255 100.635 254.395 101.675 ;
        RECT 254.715 100.635 254.855 104.055 ;
        RECT 255.175 103.355 255.315 104.735 ;
        RECT 255.635 104.375 255.775 106.775 ;
        RECT 255.575 104.055 255.835 104.375 ;
        RECT 256.025 103.860 256.305 104.230 ;
        RECT 255.115 103.035 255.375 103.355 ;
        RECT 254.195 100.315 254.455 100.635 ;
        RECT 254.655 100.315 254.915 100.635 ;
        RECT 253.335 100.065 253.935 100.205 ;
        RECT 253.795 100.035 253.935 100.065 ;
        RECT 253.795 99.955 254.395 100.035 ;
        RECT 253.795 99.895 254.455 99.955 ;
        RECT 254.195 99.635 254.455 99.895 ;
        RECT 255.175 99.355 255.315 103.035 ;
        RECT 254.255 99.215 255.315 99.355 ;
        RECT 255.575 99.295 255.835 99.615 ;
        RECT 256.095 99.525 256.235 103.860 ;
        RECT 256.555 100.295 256.695 107.795 ;
        RECT 257.415 107.115 257.675 107.435 ;
        RECT 257.475 105.395 257.615 107.115 ;
        RECT 257.415 105.075 257.675 105.395 ;
        RECT 257.645 103.520 259.185 103.890 ;
        RECT 259.255 100.315 259.515 100.635 ;
        RECT 256.495 99.975 256.755 100.295 ;
        RECT 256.955 99.635 257.215 99.955 ;
        RECT 256.095 99.385 256.695 99.525 ;
        RECT 254.255 96.555 254.395 99.215 ;
        RECT 255.635 97.915 255.775 99.295 ;
        RECT 256.035 98.615 256.295 98.935 ;
        RECT 255.575 97.595 255.835 97.915 ;
        RECT 256.095 96.895 256.235 98.615 ;
        RECT 255.575 96.575 255.835 96.895 ;
        RECT 256.035 96.575 256.295 96.895 ;
        RECT 254.195 96.235 254.455 96.555 ;
        RECT 252.815 95.895 253.075 96.215 ;
        RECT 253.275 96.070 253.535 96.215 ;
        RECT 252.875 88.395 253.015 95.895 ;
        RECT 253.265 95.700 253.545 96.070 ;
        RECT 255.635 94.855 255.775 96.575 ;
        RECT 256.555 95.955 256.695 99.385 ;
        RECT 256.095 95.815 256.695 95.955 ;
        RECT 255.575 94.535 255.835 94.855 ;
        RECT 254.195 94.195 254.455 94.515 ;
        RECT 252.815 88.075 253.075 88.395 ;
        RECT 253.725 87.540 254.005 87.910 ;
        RECT 252.815 83.315 253.075 83.635 ;
        RECT 252.875 82.470 253.015 83.315 ;
        RECT 253.275 82.635 253.535 82.955 ;
        RECT 252.805 82.100 253.085 82.470 ;
        RECT 253.335 80.235 253.475 82.635 ;
        RECT 253.275 79.915 253.535 80.235 ;
        RECT 252.355 77.875 252.615 78.195 ;
        RECT 253.795 75.385 253.935 87.540 ;
        RECT 254.255 80.915 254.395 94.195 ;
        RECT 256.095 92.135 256.235 95.815 ;
        RECT 256.495 94.195 256.755 94.515 ;
        RECT 256.035 91.815 256.295 92.135 ;
        RECT 256.035 86.035 256.295 86.355 ;
        RECT 254.655 83.995 254.915 84.315 ;
        RECT 254.195 80.595 254.455 80.915 ;
        RECT 254.715 75.815 254.855 83.995 ;
        RECT 255.115 82.975 255.375 83.295 ;
        RECT 255.175 81.595 255.315 82.975 ;
        RECT 256.095 81.675 256.235 86.035 ;
        RECT 256.555 83.975 256.695 94.195 ;
        RECT 257.015 87.910 257.155 99.635 ;
        RECT 259.315 98.935 259.455 100.315 ;
        RECT 259.775 100.295 259.915 109.415 ;
        RECT 260.625 109.225 260.905 134.520 ;
        RECT 261.095 109.495 261.355 109.815 ;
        RECT 260.695 107.435 260.835 109.225 ;
        RECT 260.635 107.115 260.895 107.435 ;
        RECT 261.155 107.095 261.295 109.495 ;
        RECT 262.925 109.225 263.205 135.100 ;
        RECT 265.225 109.225 265.505 135.680 ;
        RECT 267.525 109.225 267.805 136.260 ;
        RECT 269.825 109.225 270.105 136.840 ;
        RECT 272.125 109.225 272.405 137.420 ;
        RECT 274.425 109.225 274.705 138.000 ;
        RECT 276.725 109.225 277.005 138.580 ;
        RECT 279.025 109.225 279.305 139.160 ;
        RECT 281.325 109.225 281.605 139.740 ;
        RECT 262.995 107.775 263.135 109.225 ;
        RECT 262.935 107.455 263.195 107.775 ;
        RECT 260.175 106.775 260.435 107.095 ;
        RECT 261.095 106.775 261.355 107.095 ;
        RECT 260.235 104.375 260.375 106.775 ;
        RECT 260.945 106.240 262.485 106.610 ;
        RECT 260.635 105.075 260.895 105.395 ;
        RECT 263.395 105.075 263.655 105.395 ;
        RECT 264.775 105.075 265.035 105.395 ;
        RECT 260.175 104.055 260.435 104.375 ;
        RECT 260.695 103.355 260.835 105.075 ;
        RECT 260.635 103.035 260.895 103.355 ;
        RECT 260.635 101.905 260.895 101.995 ;
        RECT 260.235 101.765 260.895 101.905 ;
        RECT 260.235 100.635 260.375 101.765 ;
        RECT 260.635 101.675 260.895 101.765 ;
        RECT 260.945 100.800 262.485 101.170 ;
        RECT 260.175 100.315 260.435 100.635 ;
        RECT 259.715 99.975 259.975 100.295 ;
        RECT 260.625 99.780 260.905 100.150 ;
        RECT 260.635 99.635 260.895 99.780 ;
        RECT 259.715 99.295 259.975 99.615 ;
        RECT 259.255 98.615 259.515 98.935 ;
        RECT 257.645 98.080 259.185 98.450 ;
        RECT 259.775 97.995 259.915 99.295 ;
        RECT 259.315 97.855 259.915 97.995 ;
        RECT 257.405 97.060 257.685 97.430 ;
        RECT 257.475 96.895 257.615 97.060 ;
        RECT 257.415 96.575 257.675 96.895 ;
        RECT 257.415 95.895 257.675 96.215 ;
        RECT 257.475 94.710 257.615 95.895 ;
        RECT 257.405 94.340 257.685 94.710 ;
        RECT 259.315 94.515 259.455 97.855 ;
        RECT 259.715 97.255 259.975 97.575 ;
        RECT 259.775 96.895 259.915 97.255 ;
        RECT 260.695 96.895 260.835 99.635 ;
        RECT 259.715 96.575 259.975 96.895 ;
        RECT 260.175 96.750 260.435 96.895 ;
        RECT 259.255 94.195 259.515 94.515 ;
        RECT 259.775 93.235 259.915 96.575 ;
        RECT 260.165 96.380 260.445 96.750 ;
        RECT 260.635 96.575 260.895 96.895 ;
        RECT 260.945 95.360 262.485 95.730 ;
        RECT 262.475 94.535 262.735 94.855 ;
        RECT 260.175 94.195 260.435 94.515 ;
        RECT 260.635 94.195 260.895 94.515 ;
        RECT 260.235 94.030 260.375 94.195 ;
        RECT 260.165 93.660 260.445 94.030 ;
        RECT 259.775 93.095 260.375 93.235 ;
        RECT 257.645 92.640 259.185 93.010 ;
        RECT 258.795 92.155 259.055 92.475 ;
        RECT 258.325 90.940 258.605 91.310 ;
        RECT 258.395 89.755 258.535 90.940 ;
        RECT 258.335 89.435 258.595 89.755 ;
        RECT 258.855 87.965 258.995 92.155 ;
        RECT 259.255 90.795 259.515 91.115 ;
        RECT 259.315 88.305 259.455 90.795 ;
        RECT 259.705 89.580 259.985 89.950 ;
        RECT 259.775 89.415 259.915 89.580 ;
        RECT 259.715 89.095 259.975 89.415 ;
        RECT 260.235 88.395 260.375 93.095 ;
        RECT 260.695 92.475 260.835 94.195 ;
        RECT 261.555 93.175 261.815 93.495 ;
        RECT 261.615 92.475 261.755 93.175 ;
        RECT 260.635 92.155 260.895 92.475 ;
        RECT 261.555 92.155 261.815 92.475 ;
        RECT 262.535 92.135 262.675 94.535 ;
        RECT 262.935 94.195 263.195 94.515 ;
        RECT 262.475 91.815 262.735 92.135 ;
        RECT 260.945 89.920 262.485 90.290 ;
        RECT 261.555 88.755 261.815 89.075 ;
        RECT 262.475 88.755 262.735 89.075 ;
        RECT 259.315 88.165 259.915 88.305 ;
        RECT 256.945 87.540 257.225 87.910 ;
        RECT 258.855 87.825 259.455 87.965 ;
        RECT 259.315 87.795 259.455 87.825 ;
        RECT 259.315 87.655 259.500 87.795 ;
        RECT 257.645 87.200 259.185 87.570 ;
        RECT 259.360 87.115 259.500 87.655 ;
        RECT 259.775 87.230 259.915 88.165 ;
        RECT 260.175 88.075 260.435 88.395 ;
        RECT 259.315 86.975 259.500 87.115 ;
        RECT 259.315 86.605 259.455 86.975 ;
        RECT 259.705 86.860 259.985 87.230 ;
        RECT 260.235 86.695 260.375 88.075 ;
        RECT 259.315 86.465 259.915 86.605 ;
        RECT 256.955 85.695 257.215 86.015 ;
        RECT 256.495 83.655 256.755 83.975 ;
        RECT 255.115 81.275 255.375 81.595 ;
        RECT 255.635 81.535 256.235 81.675 ;
        RECT 255.635 79.895 255.775 81.535 ;
        RECT 256.555 81.255 256.695 83.655 ;
        RECT 256.495 80.935 256.755 81.255 ;
        RECT 256.555 80.575 256.695 80.935 ;
        RECT 257.015 80.575 257.155 85.695 ;
        RECT 259.775 83.975 259.915 86.465 ;
        RECT 260.175 86.375 260.435 86.695 ;
        RECT 261.615 85.335 261.755 88.755 ;
        RECT 262.535 86.355 262.675 88.755 ;
        RECT 262.475 86.035 262.735 86.355 ;
        RECT 261.555 85.015 261.815 85.335 ;
        RECT 260.945 84.480 262.485 84.850 ;
        RECT 259.715 83.655 259.975 83.975 ;
        RECT 262.995 83.715 263.135 94.195 ;
        RECT 263.455 84.225 263.595 105.075 ;
        RECT 264.315 99.635 264.575 99.955 ;
        RECT 263.855 98.615 264.115 98.935 ;
        RECT 263.915 94.515 264.055 98.615 ;
        RECT 264.375 94.855 264.515 99.635 ;
        RECT 264.315 94.535 264.575 94.855 ;
        RECT 263.855 94.195 264.115 94.515 ;
        RECT 263.915 92.670 264.055 94.195 ;
        RECT 264.375 94.175 264.515 94.535 ;
        RECT 264.315 93.855 264.575 94.175 ;
        RECT 263.845 92.300 264.125 92.670 ;
        RECT 263.855 91.135 264.115 91.455 ;
        RECT 263.915 89.075 264.055 91.135 ;
        RECT 264.315 90.795 264.575 91.115 ;
        RECT 263.855 88.755 264.115 89.075 ;
        RECT 263.455 84.085 264.055 84.225 ;
        RECT 259.255 83.315 259.515 83.635 ;
        RECT 261.095 83.315 261.355 83.635 ;
        RECT 262.995 83.575 263.595 83.715 ;
        RECT 259.315 82.355 259.455 83.315 ;
        RECT 259.315 82.215 259.500 82.355 ;
        RECT 257.645 81.760 259.185 82.130 ;
        RECT 259.360 81.675 259.500 82.215 ;
        RECT 258.795 81.275 259.055 81.595 ;
        RECT 259.315 81.535 259.500 81.675 ;
        RECT 258.855 80.575 258.995 81.275 ;
        RECT 256.495 80.255 256.755 80.575 ;
        RECT 256.955 80.485 257.215 80.575 ;
        RECT 258.335 80.485 258.595 80.575 ;
        RECT 256.955 80.345 257.615 80.485 ;
        RECT 256.955 80.255 257.215 80.345 ;
        RECT 255.575 79.575 255.835 79.895 ;
        RECT 256.035 78.215 256.295 78.535 ;
        RECT 255.115 77.875 255.375 78.195 ;
        RECT 255.175 76.155 255.315 77.875 ;
        RECT 255.115 75.835 255.375 76.155 ;
        RECT 254.655 75.495 254.915 75.815 ;
        RECT 253.795 75.245 254.395 75.385 ;
        RECT 253.725 74.620 254.005 74.990 ;
        RECT 251.895 72.775 252.155 73.095 ;
        RECT 245.455 65.975 245.715 66.295 ;
        RECT 245.445 64.420 245.725 64.790 ;
        RECT 245.515 64.255 245.655 64.420 ;
        RECT 244.995 63.935 245.255 64.255 ;
        RECT 245.455 63.935 245.715 64.255 ;
        RECT 244.595 63.345 245.195 63.485 ;
        RECT 244.075 61.895 244.335 62.215 ;
        RECT 245.055 61.535 245.195 63.345 ;
        RECT 244.535 61.215 244.795 61.535 ;
        RECT 244.995 61.215 245.255 61.535 ;
        RECT 244.595 59.835 244.735 61.215 ;
        RECT 243.215 59.455 243.815 59.595 ;
        RECT 244.535 59.515 244.795 59.835 ;
        RECT 245.975 59.495 246.115 69.375 ;
        RECT 247.745 69.180 248.025 69.550 ;
        RECT 250.965 69.180 251.245 69.550 ;
        RECT 249.135 68.695 249.395 69.015 ;
        RECT 249.195 67.655 249.335 68.695 ;
        RECT 250.045 68.500 250.325 68.870 ;
        RECT 249.135 67.335 249.395 67.655 ;
        RECT 248.675 66.995 248.935 67.315 ;
        RECT 248.735 66.830 248.875 66.995 ;
        RECT 248.665 66.460 248.945 66.830 ;
        RECT 246.375 65.975 246.635 66.295 ;
        RECT 246.435 59.835 246.575 65.975 ;
        RECT 250.115 64.935 250.255 68.500 ;
        RECT 250.055 64.615 250.315 64.935 ;
        RECT 246.835 63.255 247.095 63.575 ;
        RECT 246.895 61.875 247.035 63.255 ;
        RECT 246.835 61.555 247.095 61.875 ;
        RECT 247.295 61.555 247.555 61.875 ;
        RECT 248.665 61.700 248.945 62.070 ;
        RECT 250.115 61.875 250.255 64.615 ;
        RECT 251.435 62.235 251.695 62.555 ;
        RECT 248.675 61.555 248.935 61.700 ;
        RECT 250.055 61.555 250.315 61.875 ;
        RECT 246.375 59.515 246.635 59.835 ;
        RECT 243.675 57.195 243.815 59.455 ;
        RECT 244.065 58.980 244.345 59.350 ;
        RECT 245.915 59.175 246.175 59.495 ;
        RECT 246.895 59.235 247.035 61.555 ;
        RECT 246.435 59.095 247.035 59.235 ;
        RECT 244.075 58.835 244.335 58.980 ;
        RECT 246.435 58.135 246.575 59.095 ;
        RECT 246.375 57.815 246.635 58.135 ;
        RECT 243.675 57.055 244.275 57.195 ;
        RECT 243.155 56.685 243.415 56.775 ;
        RECT 243.155 56.545 243.815 56.685 ;
        RECT 243.155 56.455 243.415 56.545 ;
        RECT 243.155 55.095 243.415 55.415 ;
        RECT 242.235 53.395 242.495 53.715 ;
        RECT 241.315 52.375 241.575 52.695 ;
        RECT 240.395 47.615 240.655 47.935 ;
        RECT 240.455 45.895 240.595 47.615 ;
        RECT 240.395 45.805 240.655 45.895 ;
        RECT 240.395 45.665 241.055 45.805 ;
        RECT 240.395 45.575 240.655 45.665 ;
        RECT 239.935 45.235 240.195 45.555 ;
        RECT 239.475 41.495 239.735 41.815 ;
        RECT 239.995 40.795 240.135 45.235 ;
        RECT 240.385 44.020 240.665 44.390 ;
        RECT 240.455 42.495 240.595 44.020 ;
        RECT 240.395 42.175 240.655 42.495 ;
        RECT 239.935 40.475 240.195 40.795 ;
        RECT 238.555 39.795 238.815 40.115 ;
        RECT 240.915 37.395 241.055 45.665 ;
        RECT 241.375 45.215 241.515 52.375 ;
        RECT 242.225 49.460 242.505 49.830 ;
        RECT 242.695 49.655 242.955 49.975 ;
        RECT 241.765 46.740 242.045 47.110 ;
        RECT 241.835 45.215 241.975 46.740 ;
        RECT 242.295 45.555 242.435 49.460 ;
        RECT 242.755 48.275 242.895 49.655 ;
        RECT 242.695 47.955 242.955 48.275 ;
        RECT 242.695 47.275 242.955 47.595 ;
        RECT 242.755 46.235 242.895 47.275 ;
        RECT 242.695 45.915 242.955 46.235 ;
        RECT 242.235 45.235 242.495 45.555 ;
        RECT 242.685 45.380 242.965 45.750 ;
        RECT 242.695 45.235 242.955 45.380 ;
        RECT 241.315 44.895 241.575 45.215 ;
        RECT 241.775 44.895 242.035 45.215 ;
        RECT 242.295 42.495 242.435 45.235 ;
        RECT 242.695 44.215 242.955 44.535 ;
        RECT 242.755 42.835 242.895 44.215 ;
        RECT 242.695 42.515 242.955 42.835 ;
        RECT 243.215 42.495 243.355 55.095 ;
        RECT 243.675 53.375 243.815 56.545 ;
        RECT 243.615 53.055 243.875 53.375 ;
        RECT 243.675 44.875 243.815 53.055 ;
        RECT 243.615 44.555 243.875 44.875 ;
        RECT 242.235 42.175 242.495 42.495 ;
        RECT 243.155 42.175 243.415 42.495 ;
        RECT 241.775 41.495 242.035 41.815 ;
        RECT 241.835 40.115 241.975 41.495 ;
        RECT 244.135 40.795 244.275 57.055 ;
        RECT 245.445 56.940 245.725 57.310 ;
        RECT 244.535 50.335 244.795 50.655 ;
        RECT 244.595 46.235 244.735 50.335 ;
        RECT 244.995 47.275 245.255 47.595 ;
        RECT 244.535 45.915 244.795 46.235 ;
        RECT 245.055 45.895 245.195 47.275 ;
        RECT 244.995 45.575 245.255 45.895 ;
        RECT 244.075 40.475 244.335 40.795 ;
        RECT 241.775 39.795 242.035 40.115 ;
        RECT 242.235 38.775 242.495 39.095 ;
        RECT 243.155 38.775 243.415 39.095 ;
        RECT 242.295 37.395 242.435 38.775 ;
        RECT 240.855 37.305 241.115 37.395 ;
        RECT 240.455 37.165 241.115 37.305 ;
        RECT 237.635 34.695 237.895 35.015 ;
        RECT 237.695 31.275 237.835 34.695 ;
        RECT 240.455 34.675 240.595 37.165 ;
        RECT 240.855 37.075 241.115 37.165 ;
        RECT 242.235 37.075 242.495 37.395 ;
        RECT 241.775 36.395 242.035 36.715 ;
        RECT 240.395 34.355 240.655 34.675 ;
        RECT 241.835 31.275 241.975 36.395 ;
        RECT 243.215 35.015 243.355 38.775 ;
        RECT 245.055 37.395 245.195 45.575 ;
        RECT 244.995 37.075 245.255 37.395 ;
        RECT 245.055 36.715 245.195 37.075 ;
        RECT 244.995 36.395 245.255 36.715 ;
        RECT 245.055 35.015 245.195 36.395 ;
        RECT 243.155 34.695 243.415 35.015 ;
        RECT 244.995 34.695 245.255 35.015 ;
        RECT 245.515 31.615 245.655 56.940 ;
        RECT 245.915 55.775 246.175 56.095 ;
        RECT 245.975 48.955 246.115 55.775 ;
        RECT 247.355 50.510 247.495 61.555 ;
        RECT 248.215 61.215 248.475 61.535 ;
        RECT 248.275 60.855 248.415 61.215 ;
        RECT 249.595 60.875 249.855 61.195 ;
        RECT 248.215 60.535 248.475 60.855 ;
        RECT 248.275 58.475 248.415 60.535 ;
        RECT 249.655 59.155 249.795 60.875 ;
        RECT 249.595 58.835 249.855 59.155 ;
        RECT 248.215 58.155 248.475 58.475 ;
        RECT 249.585 58.300 249.865 58.670 ;
        RECT 248.275 57.990 248.415 58.155 ;
        RECT 249.655 58.135 249.795 58.300 ;
        RECT 248.205 57.620 248.485 57.990 ;
        RECT 249.595 57.815 249.855 58.135 ;
        RECT 249.655 57.115 249.795 57.815 ;
        RECT 249.595 56.795 249.855 57.115 ;
        RECT 250.055 56.795 250.315 57.115 ;
        RECT 247.755 53.735 248.015 54.055 ;
        RECT 247.815 53.375 247.955 53.735 ;
        RECT 247.755 53.055 248.015 53.375 ;
        RECT 250.115 52.695 250.255 56.795 ;
        RECT 251.495 56.775 251.635 62.235 ;
        RECT 253.795 62.070 253.935 74.620 ;
        RECT 254.255 67.655 254.395 75.245 ;
        RECT 255.115 75.155 255.375 75.475 ;
        RECT 255.175 74.990 255.315 75.155 ;
        RECT 255.105 74.620 255.385 74.990 ;
        RECT 254.195 67.335 254.455 67.655 ;
        RECT 254.255 63.915 254.395 67.335 ;
        RECT 255.175 66.975 255.315 74.620 ;
        RECT 256.095 72.755 256.235 78.215 ;
        RECT 256.485 78.020 256.765 78.390 ;
        RECT 256.555 77.855 256.695 78.020 ;
        RECT 256.495 77.535 256.755 77.855 ;
        RECT 256.035 72.435 256.295 72.755 ;
        RECT 256.035 71.755 256.295 72.075 ;
        RECT 256.095 67.995 256.235 71.755 ;
        RECT 256.555 70.035 256.695 77.535 ;
        RECT 257.475 77.085 257.615 80.345 ;
        RECT 257.935 80.345 258.595 80.485 ;
        RECT 257.935 78.535 258.075 80.345 ;
        RECT 258.335 80.255 258.595 80.345 ;
        RECT 258.795 80.255 259.055 80.575 ;
        RECT 258.795 79.575 259.055 79.895 ;
        RECT 258.855 78.875 258.995 79.575 ;
        RECT 258.335 78.555 258.595 78.875 ;
        RECT 258.795 78.555 259.055 78.875 ;
        RECT 257.875 78.215 258.135 78.535 ;
        RECT 258.395 78.390 258.535 78.555 ;
        RECT 258.325 78.020 258.605 78.390 ;
        RECT 259.315 78.275 259.455 81.535 ;
        RECT 261.155 80.995 261.295 83.315 ;
        RECT 262.935 82.975 263.195 83.295 ;
        RECT 262.005 81.420 262.285 81.790 ;
        RECT 262.995 81.595 263.135 82.975 ;
        RECT 259.775 80.855 261.295 80.995 ;
        RECT 259.775 78.875 259.915 80.855 ;
        RECT 261.545 80.740 261.825 81.110 ;
        RECT 260.635 80.485 260.895 80.575 ;
        RECT 260.235 80.345 260.895 80.485 ;
        RECT 259.715 78.555 259.975 78.875 ;
        RECT 258.335 77.875 258.595 78.020 ;
        RECT 258.795 77.875 259.055 78.195 ;
        RECT 259.315 78.135 259.915 78.275 ;
        RECT 257.875 77.595 258.135 77.855 ;
        RECT 258.855 77.595 258.995 77.875 ;
        RECT 257.875 77.535 258.995 77.595 ;
        RECT 257.935 77.455 258.995 77.535 ;
        RECT 259.245 77.340 259.525 77.710 ;
        RECT 259.315 77.175 259.455 77.340 ;
        RECT 257.020 76.945 257.615 77.085 ;
        RECT 257.020 76.065 257.160 76.945 ;
        RECT 259.255 76.855 259.515 77.175 ;
        RECT 257.645 76.320 259.185 76.690 ;
        RECT 259.775 76.350 259.915 78.135 ;
        RECT 257.020 75.925 257.615 76.065 ;
        RECT 257.475 75.475 257.615 75.925 ;
        RECT 258.335 75.835 258.595 76.155 ;
        RECT 258.795 75.835 259.055 76.155 ;
        RECT 259.705 75.980 259.985 76.350 ;
        RECT 257.415 75.155 257.675 75.475 ;
        RECT 257.875 74.815 258.135 75.135 ;
        RECT 257.415 74.475 257.675 74.795 ;
        RECT 256.955 74.135 257.215 74.455 ;
        RECT 257.015 72.075 257.155 74.135 ;
        RECT 257.475 73.630 257.615 74.475 ;
        RECT 257.935 74.310 258.075 74.815 ;
        RECT 257.865 73.940 258.145 74.310 ;
        RECT 257.405 73.260 257.685 73.630 ;
        RECT 257.935 73.435 258.075 73.940 ;
        RECT 257.875 73.115 258.135 73.435 ;
        RECT 258.395 72.325 258.535 75.835 ;
        RECT 258.855 73.095 258.995 75.835 ;
        RECT 259.715 75.495 259.975 75.815 ;
        RECT 259.775 74.310 259.915 75.495 ;
        RECT 260.235 74.365 260.375 80.345 ;
        RECT 260.635 80.255 260.895 80.345 ;
        RECT 261.615 80.235 261.755 80.740 ;
        RECT 262.075 80.235 262.215 81.420 ;
        RECT 262.935 81.275 263.195 81.595 ;
        RECT 262.925 80.740 263.205 81.110 ;
        RECT 261.555 79.915 261.815 80.235 ;
        RECT 262.015 79.915 262.275 80.235 ;
        RECT 260.945 79.040 262.485 79.410 ;
        RECT 261.095 78.555 261.355 78.875 ;
        RECT 262.995 78.785 263.135 80.740 ;
        RECT 261.615 78.645 263.135 78.785 ;
        RECT 260.635 77.875 260.895 78.195 ;
        RECT 260.695 77.710 260.835 77.875 ;
        RECT 261.155 77.855 261.295 78.555 ;
        RECT 261.615 78.195 261.755 78.645 ;
        RECT 263.455 78.275 263.595 83.575 ;
        RECT 263.915 81.790 264.055 84.085 ;
        RECT 263.845 81.420 264.125 81.790 ;
        RECT 264.375 80.995 264.515 90.795 ;
        RECT 264.835 86.015 264.975 105.075 ;
        RECT 265.295 103.355 265.435 109.225 ;
        RECT 267.595 105.735 267.735 109.225 ;
        RECT 269.895 106.155 270.035 109.225 ;
        RECT 271.675 107.795 271.935 108.115 ;
        RECT 271.735 107.095 271.875 107.795 ;
        RECT 272.195 107.095 272.335 109.225 ;
        RECT 272.595 108.135 272.855 108.455 ;
        RECT 271.675 106.775 271.935 107.095 ;
        RECT 272.135 106.775 272.395 107.095 ;
        RECT 269.895 106.015 270.495 106.155 ;
        RECT 267.535 105.415 267.795 105.735 ;
        RECT 268.515 105.395 270.035 105.475 ;
        RECT 268.515 105.335 270.095 105.395 ;
        RECT 267.535 104.735 267.795 105.055 ;
        RECT 267.995 104.735 268.255 105.055 ;
        RECT 265.235 103.035 265.495 103.355 ;
        RECT 266.155 102.355 266.415 102.675 ;
        RECT 265.695 101.675 265.955 101.995 ;
        RECT 265.755 100.635 265.895 101.675 ;
        RECT 265.695 100.315 265.955 100.635 ;
        RECT 265.695 98.615 265.955 98.935 ;
        RECT 265.755 96.555 265.895 98.615 ;
        RECT 265.695 96.235 265.955 96.555 ;
        RECT 265.235 91.310 265.495 91.455 ;
        RECT 265.225 90.940 265.505 91.310 ;
        RECT 265.235 90.455 265.495 90.775 ;
        RECT 264.775 85.695 265.035 86.015 ;
        RECT 264.775 82.295 265.035 82.615 ;
        RECT 264.835 81.255 264.975 82.295 ;
        RECT 261.555 77.875 261.815 78.195 ;
        RECT 262.015 77.875 262.275 78.195 ;
        RECT 262.535 78.135 263.595 78.275 ;
        RECT 263.915 80.855 264.515 80.995 ;
        RECT 264.775 80.935 265.035 81.255 ;
        RECT 265.295 81.110 265.435 90.455 ;
        RECT 266.215 88.735 266.355 102.355 ;
        RECT 267.595 96.895 267.735 104.735 ;
        RECT 268.055 98.935 268.195 104.735 ;
        RECT 268.515 103.015 268.655 105.335 ;
        RECT 269.835 105.075 270.095 105.335 ;
        RECT 270.355 104.715 270.495 106.015 ;
        RECT 270.295 104.395 270.555 104.715 ;
        RECT 270.755 104.055 271.015 104.375 ;
        RECT 268.455 102.695 268.715 103.015 ;
        RECT 267.995 98.615 268.255 98.935 ;
        RECT 267.535 96.575 267.795 96.895 ;
        RECT 268.515 95.195 268.655 102.695 ;
        RECT 269.835 101.335 270.095 101.655 ;
        RECT 269.895 99.615 270.035 101.335 ;
        RECT 269.835 99.295 270.095 99.615 ;
        RECT 269.375 96.575 269.635 96.895 ;
        RECT 268.455 94.875 268.715 95.195 ;
        RECT 269.435 92.475 269.575 96.575 ;
        RECT 267.995 92.155 268.255 92.475 ;
        RECT 269.375 92.155 269.635 92.475 ;
        RECT 267.535 91.135 267.795 91.455 ;
        RECT 266.615 90.455 266.875 90.775 ;
        RECT 266.675 88.735 266.815 90.455 ;
        RECT 267.595 89.755 267.735 91.135 ;
        RECT 267.535 89.435 267.795 89.755 ;
        RECT 266.155 88.415 266.415 88.735 ;
        RECT 266.615 88.415 266.875 88.735 ;
        RECT 266.215 86.015 266.355 88.415 ;
        RECT 268.055 88.395 268.195 92.155 ;
        RECT 268.455 90.795 268.715 91.115 ;
        RECT 267.995 88.075 268.255 88.395 ;
        RECT 266.155 85.695 266.415 86.015 ;
        RECT 266.615 85.015 266.875 85.335 ;
        RECT 266.675 83.635 266.815 85.015 ;
        RECT 266.615 83.545 266.875 83.635 ;
        RECT 266.215 83.405 266.875 83.545 ;
        RECT 260.625 77.340 260.905 77.710 ;
        RECT 261.095 77.535 261.355 77.855 ;
        RECT 262.075 77.175 262.215 77.875 ;
        RECT 262.015 76.855 262.275 77.175 ;
        RECT 262.005 75.980 262.285 76.350 ;
        RECT 262.535 76.155 262.675 78.135 ;
        RECT 263.915 78.105 264.055 80.855 ;
        RECT 265.225 80.740 265.505 81.110 ;
        RECT 264.315 80.430 264.575 80.575 ;
        RECT 265.695 80.485 265.955 80.575 ;
        RECT 266.215 80.485 266.355 83.405 ;
        RECT 266.615 83.315 266.875 83.405 ;
        RECT 267.535 82.975 267.795 83.295 ;
        RECT 267.075 81.275 267.335 81.595 ;
        RECT 264.305 80.060 264.585 80.430 ;
        RECT 265.695 80.345 266.355 80.485 ;
        RECT 265.695 80.255 265.955 80.345 ;
        RECT 264.775 79.575 265.035 79.895 ;
        RECT 263.915 77.965 264.515 78.105 ;
        RECT 263.845 77.340 264.125 77.710 ;
        RECT 262.935 76.855 263.195 77.175 ;
        RECT 261.545 75.300 261.825 75.670 ;
        RECT 261.615 75.135 261.755 75.300 ;
        RECT 262.075 75.135 262.215 75.980 ;
        RECT 262.475 75.835 262.735 76.155 ;
        RECT 262.535 75.135 262.675 75.835 ;
        RECT 262.995 75.135 263.135 76.855 ;
        RECT 261.555 74.815 261.815 75.135 ;
        RECT 262.015 74.815 262.275 75.135 ;
        RECT 262.475 74.815 262.735 75.135 ;
        RECT 262.935 74.815 263.195 75.135 ;
        RECT 259.705 73.940 259.985 74.310 ;
        RECT 260.235 74.225 263.135 74.365 ;
        RECT 259.775 73.345 259.915 73.940 ;
        RECT 260.945 73.600 262.485 73.970 ;
        RECT 259.775 73.205 261.295 73.345 ;
        RECT 258.795 72.775 259.055 73.095 ;
        RECT 260.635 72.435 260.895 72.755 ;
        RECT 258.395 72.185 259.455 72.325 ;
        RECT 256.955 71.755 257.215 72.075 ;
        RECT 259.315 71.475 259.455 72.185 ;
        RECT 260.175 71.755 260.435 72.075 ;
        RECT 259.315 71.335 259.500 71.475 ;
        RECT 259.715 71.415 259.975 71.735 ;
        RECT 256.945 70.540 257.225 70.910 ;
        RECT 257.645 70.880 259.185 71.250 ;
        RECT 259.360 70.795 259.500 71.335 ;
        RECT 259.315 70.655 259.500 70.795 ;
        RECT 256.955 70.395 257.215 70.540 ;
        RECT 258.795 70.055 259.055 70.375 ;
        RECT 256.495 69.715 256.755 70.035 ;
        RECT 256.955 69.375 257.215 69.695 ;
        RECT 256.495 69.035 256.755 69.355 ;
        RECT 256.035 67.675 256.295 67.995 ;
        RECT 256.035 66.995 256.295 67.315 ;
        RECT 255.115 66.655 255.375 66.975 ;
        RECT 255.575 64.955 255.835 65.275 ;
        RECT 254.195 63.595 254.455 63.915 ;
        RECT 253.725 61.700 254.005 62.070 ;
        RECT 253.735 61.555 253.995 61.700 ;
        RECT 255.635 61.390 255.775 64.955 ;
        RECT 255.565 61.020 255.845 61.390 ;
        RECT 256.095 61.195 256.235 66.995 ;
        RECT 255.635 60.855 255.775 61.020 ;
        RECT 256.035 60.875 256.295 61.195 ;
        RECT 255.575 60.535 255.835 60.855 ;
        RECT 252.815 59.405 253.075 59.495 ;
        RECT 252.815 59.265 253.475 59.405 ;
        RECT 252.815 59.175 253.075 59.265 ;
        RECT 252.815 58.495 253.075 58.815 ;
        RECT 251.435 56.455 251.695 56.775 ;
        RECT 252.875 56.095 253.015 58.495 ;
        RECT 253.335 58.385 253.475 59.265 ;
        RECT 256.555 59.155 256.695 69.035 ;
        RECT 257.015 62.215 257.155 69.375 ;
        RECT 258.855 67.315 258.995 70.055 ;
        RECT 259.315 70.035 259.455 70.655 ;
        RECT 259.255 69.715 259.515 70.035 ;
        RECT 259.255 69.035 259.515 69.355 ;
        RECT 259.315 67.995 259.455 69.035 ;
        RECT 259.775 67.995 259.915 71.415 ;
        RECT 259.255 67.675 259.515 67.995 ;
        RECT 259.715 67.675 259.975 67.995 ;
        RECT 259.245 67.395 259.525 67.510 ;
        RECT 258.795 66.995 259.055 67.315 ;
        RECT 259.245 67.255 259.915 67.395 ;
        RECT 259.245 67.140 259.525 67.255 ;
        RECT 257.865 66.460 258.145 66.830 ;
        RECT 259.775 66.635 259.915 67.255 ;
        RECT 260.235 66.975 260.375 71.755 ;
        RECT 260.695 70.035 260.835 72.435 ;
        RECT 260.635 69.715 260.895 70.035 ;
        RECT 261.155 69.695 261.295 73.205 ;
        RECT 261.555 73.115 261.815 73.435 ;
        RECT 261.615 72.950 261.755 73.115 ;
        RECT 261.545 72.580 261.825 72.950 ;
        RECT 262.465 72.580 262.745 72.950 ;
        RECT 262.475 72.435 262.735 72.580 ;
        RECT 262.475 71.415 262.735 71.735 ;
        RECT 261.545 70.540 261.825 70.910 ;
        RECT 261.555 70.395 261.815 70.540 ;
        RECT 262.535 69.695 262.675 71.415 ;
        RECT 261.095 69.375 261.355 69.695 ;
        RECT 262.475 69.375 262.735 69.695 ;
        RECT 260.945 68.160 262.485 68.530 ;
        RECT 262.995 67.395 263.135 74.225 ;
        RECT 263.395 74.135 263.655 74.455 ;
        RECT 263.455 67.655 263.595 74.135 ;
        RECT 263.915 72.415 264.055 77.340 ;
        RECT 264.375 76.350 264.515 77.965 ;
        RECT 264.305 75.980 264.585 76.350 ;
        RECT 264.315 75.155 264.575 75.475 ;
        RECT 263.855 72.095 264.115 72.415 ;
        RECT 264.375 69.695 264.515 75.155 ;
        RECT 264.835 72.755 264.975 79.575 ;
        RECT 267.135 78.875 267.275 81.275 ;
        RECT 267.075 78.555 267.335 78.875 ;
        RECT 266.605 78.020 266.885 78.390 ;
        RECT 266.615 77.875 266.875 78.020 ;
        RECT 265.235 77.535 265.495 77.855 ;
        RECT 265.295 74.990 265.435 77.535 ;
        RECT 267.595 77.175 267.735 82.975 ;
        RECT 267.985 81.420 268.265 81.790 ;
        RECT 267.535 76.855 267.795 77.175 ;
        RECT 265.225 74.620 265.505 74.990 ;
        RECT 265.695 74.815 265.955 75.135 ;
        RECT 265.235 74.135 265.495 74.455 ;
        RECT 264.775 72.435 265.035 72.755 ;
        RECT 265.295 69.695 265.435 74.135 ;
        RECT 265.755 73.435 265.895 74.815 ;
        RECT 268.055 73.435 268.195 81.420 ;
        RECT 268.515 80.995 268.655 90.795 ;
        RECT 268.915 90.455 269.175 90.775 ;
        RECT 268.975 88.590 269.115 90.455 ;
        RECT 268.905 88.220 269.185 88.590 ;
        RECT 270.815 87.035 270.955 104.055 ;
        RECT 272.655 102.675 272.795 108.135 ;
        RECT 273.515 107.115 273.775 107.435 ;
        RECT 273.575 106.075 273.715 107.115 ;
        RECT 273.515 105.755 273.775 106.075 ;
        RECT 274.495 104.375 274.635 109.225 ;
        RECT 275.815 107.455 276.075 107.775 ;
        RECT 275.875 106.075 276.015 107.455 ;
        RECT 275.815 105.755 276.075 106.075 ;
        RECT 276.795 105.055 276.935 109.225 ;
        RECT 279.095 107.435 279.235 109.225 ;
        RECT 279.035 107.115 279.295 107.435 ;
        RECT 281.395 105.735 281.535 109.225 ;
        RECT 282.255 109.155 282.515 109.475 ;
        RECT 283.625 109.225 283.905 140.320 ;
        RECT 285.925 109.225 286.205 140.900 ;
        RECT 288.225 109.225 288.505 141.480 ;
        RECT 290.525 109.225 290.805 142.060 ;
        RECT 292.825 109.225 293.105 142.640 ;
        RECT 295.125 109.225 295.405 143.220 ;
        RECT 297.425 109.225 297.705 143.800 ;
        RECT 299.725 109.225 300.005 144.380 ;
        RECT 302.025 109.225 302.305 144.960 ;
        RECT 304.325 109.225 304.605 145.540 ;
        RECT 306.625 109.225 306.905 146.120 ;
        RECT 308.925 109.225 309.205 146.700 ;
        RECT 281.335 105.415 281.595 105.735 ;
        RECT 279.495 105.075 279.755 105.395 ;
        RECT 281.795 105.075 282.055 105.395 ;
        RECT 276.735 104.735 276.995 105.055 ;
        RECT 273.055 104.055 273.315 104.375 ;
        RECT 274.435 104.055 274.695 104.375 ;
        RECT 272.135 102.355 272.395 102.675 ;
        RECT 272.595 102.355 272.855 102.675 ;
        RECT 272.195 97.235 272.335 102.355 ;
        RECT 273.115 102.335 273.255 104.055 ;
        RECT 279.035 102.355 279.295 102.675 ;
        RECT 273.055 102.015 273.315 102.335 ;
        RECT 277.655 101.675 277.915 101.995 ;
        RECT 274.895 101.335 275.155 101.655 ;
        RECT 274.955 100.295 275.095 101.335 ;
        RECT 274.895 99.975 275.155 100.295 ;
        RECT 276.275 99.295 276.535 99.615 ;
        RECT 276.335 97.915 276.475 99.295 ;
        RECT 276.275 97.595 276.535 97.915 ;
        RECT 272.135 96.915 272.395 97.235 ;
        RECT 277.195 96.915 277.455 97.235 ;
        RECT 277.255 95.195 277.395 96.915 ;
        RECT 277.195 94.875 277.455 95.195 ;
        RECT 276.725 94.340 277.005 94.710 ;
        RECT 276.795 94.175 276.935 94.340 ;
        RECT 276.735 93.855 276.995 94.175 ;
        RECT 277.255 93.495 277.395 94.875 ;
        RECT 275.815 93.175 276.075 93.495 ;
        RECT 277.195 93.175 277.455 93.495 ;
        RECT 275.875 88.735 276.015 93.175 ;
        RECT 277.715 91.115 277.855 101.675 ;
        RECT 279.095 98.935 279.235 102.355 ;
        RECT 279.035 98.615 279.295 98.935 ;
        RECT 278.105 97.060 278.385 97.430 ;
        RECT 279.095 97.235 279.235 98.615 ;
        RECT 278.175 96.215 278.315 97.060 ;
        RECT 279.035 96.915 279.295 97.235 ;
        RECT 278.565 96.380 278.845 96.750 ;
        RECT 278.115 95.895 278.375 96.215 ;
        RECT 278.175 94.515 278.315 95.895 ;
        RECT 278.635 94.515 278.775 96.380 ;
        RECT 278.115 94.195 278.375 94.515 ;
        RECT 278.575 94.195 278.835 94.515 ;
        RECT 278.575 93.515 278.835 93.835 ;
        RECT 278.635 91.795 278.775 93.515 ;
        RECT 278.575 91.475 278.835 91.795 ;
        RECT 278.115 91.135 278.375 91.455 ;
        RECT 277.655 90.795 277.915 91.115 ;
        RECT 276.275 90.455 276.535 90.775 ;
        RECT 275.815 88.415 276.075 88.735 ;
        RECT 276.335 88.055 276.475 90.455 ;
        RECT 277.655 89.435 277.915 89.755 ;
        RECT 277.715 89.270 277.855 89.435 ;
        RECT 276.735 88.755 276.995 89.075 ;
        RECT 277.645 88.900 277.925 89.270 ;
        RECT 276.275 87.735 276.535 88.055 ;
        RECT 276.795 87.035 276.935 88.755 ;
        RECT 270.755 86.715 271.015 87.035 ;
        RECT 276.735 86.715 276.995 87.035 ;
        RECT 270.295 85.355 270.555 85.675 ;
        RECT 269.365 82.780 269.645 83.150 ;
        RECT 269.435 81.595 269.575 82.780 ;
        RECT 269.375 81.275 269.635 81.595 ;
        RECT 268.515 80.855 269.115 80.995 ;
        RECT 268.455 80.255 268.715 80.575 ;
        RECT 268.515 78.875 268.655 80.255 ;
        RECT 268.455 78.555 268.715 78.875 ;
        RECT 268.455 77.195 268.715 77.515 ;
        RECT 268.515 75.135 268.655 77.195 ;
        RECT 268.455 74.815 268.715 75.135 ;
        RECT 265.695 73.345 265.955 73.435 ;
        RECT 265.695 73.205 266.815 73.345 ;
        RECT 265.695 73.115 265.955 73.205 ;
        RECT 265.695 70.055 265.955 70.375 ;
        RECT 265.755 69.695 265.895 70.055 ;
        RECT 266.675 70.035 266.815 73.205 ;
        RECT 267.995 73.115 268.255 73.435 ;
        RECT 266.615 69.715 266.875 70.035 ;
        RECT 264.315 69.375 264.575 69.695 ;
        RECT 265.235 69.375 265.495 69.695 ;
        RECT 265.695 69.375 265.955 69.695 ;
        RECT 264.375 67.655 264.515 69.375 ;
        RECT 268.055 69.355 268.195 73.115 ;
        RECT 268.975 72.950 269.115 80.855 ;
        RECT 269.365 80.060 269.645 80.430 ;
        RECT 269.835 80.255 270.095 80.575 ;
        RECT 268.905 72.580 269.185 72.950 ;
        RECT 267.995 69.035 268.255 69.355 ;
        RECT 262.535 67.255 263.135 67.395 ;
        RECT 263.395 67.335 263.655 67.655 ;
        RECT 264.315 67.335 264.575 67.655 ;
        RECT 260.175 66.655 260.435 66.975 ;
        RECT 257.875 66.315 258.135 66.460 ;
        RECT 259.255 66.315 259.515 66.635 ;
        RECT 259.715 66.315 259.975 66.635 ;
        RECT 259.315 66.035 259.455 66.315 ;
        RECT 259.315 65.895 259.915 66.035 ;
        RECT 257.645 65.440 259.185 65.810 ;
        RECT 259.245 63.740 259.525 64.110 ;
        RECT 259.255 63.595 259.515 63.740 ;
        RECT 257.415 63.255 257.675 63.575 ;
        RECT 256.955 61.895 257.215 62.215 ;
        RECT 257.475 61.875 257.615 63.255 ;
        RECT 259.315 62.555 259.455 63.595 ;
        RECT 258.795 62.235 259.055 62.555 ;
        RECT 259.255 62.235 259.515 62.555 ;
        RECT 258.855 61.955 258.995 62.235 ;
        RECT 259.775 61.955 259.915 65.895 ;
        RECT 260.175 63.935 260.435 64.255 ;
        RECT 257.415 61.555 257.675 61.875 ;
        RECT 258.855 61.815 259.915 61.955 ;
        RECT 260.235 61.875 260.375 63.935 ;
        RECT 262.535 63.485 262.675 67.255 ;
        RECT 264.375 66.830 264.515 67.335 ;
        RECT 264.305 66.460 264.585 66.830 ;
        RECT 268.975 66.635 269.115 72.580 ;
        RECT 269.435 72.075 269.575 80.060 ;
        RECT 269.375 71.755 269.635 72.075 ;
        RECT 269.895 69.695 270.035 80.255 ;
        RECT 270.355 75.815 270.495 85.355 ;
        RECT 270.295 75.495 270.555 75.815 ;
        RECT 270.815 74.795 270.955 86.715 ;
        RECT 276.275 86.375 276.535 86.695 ;
        RECT 271.675 83.655 271.935 83.975 ;
        RECT 270.755 74.475 271.015 74.795 ;
        RECT 271.735 74.455 271.875 83.655 ;
        RECT 276.335 81.595 276.475 86.375 ;
        RECT 276.275 81.275 276.535 81.595 ;
        RECT 275.815 80.255 276.075 80.575 ;
        RECT 275.355 76.855 275.615 77.175 ;
        RECT 275.415 74.795 275.555 76.855 ;
        RECT 275.355 74.475 275.615 74.795 ;
        RECT 270.295 74.135 270.555 74.455 ;
        RECT 271.675 74.135 271.935 74.455 ;
        RECT 272.135 74.135 272.395 74.455 ;
        RECT 270.355 71.735 270.495 74.135 ;
        RECT 272.195 72.415 272.335 74.135 ;
        RECT 272.135 72.095 272.395 72.415 ;
        RECT 275.355 71.755 275.615 72.075 ;
        RECT 270.295 71.415 270.555 71.735 ;
        RECT 269.835 69.375 270.095 69.695 ;
        RECT 268.915 66.315 269.175 66.635 ;
        RECT 269.895 63.575 270.035 69.375 ;
        RECT 262.535 63.345 263.135 63.485 ;
        RECT 260.945 62.720 262.485 63.090 ;
        RECT 262.995 62.555 263.135 63.345 ;
        RECT 269.835 63.255 270.095 63.575 ;
        RECT 262.935 62.235 263.195 62.555 ;
        RECT 257.645 60.000 259.185 60.370 ;
        RECT 256.495 58.835 256.755 59.155 ;
        RECT 253.735 58.385 253.995 58.475 ;
        RECT 253.335 58.245 253.995 58.385 ;
        RECT 253.735 58.155 253.995 58.245 ;
        RECT 259.255 58.155 259.515 58.475 ;
        RECT 254.655 57.990 254.915 58.135 ;
        RECT 254.645 57.620 254.925 57.990 ;
        RECT 256.025 56.940 256.305 57.310 ;
        RECT 256.095 56.775 256.235 56.940 ;
        RECT 256.035 56.455 256.295 56.775 ;
        RECT 252.815 55.775 253.075 56.095 ;
        RECT 254.655 55.775 254.915 56.095 ;
        RECT 253.275 55.095 253.535 55.415 ;
        RECT 252.355 52.715 252.615 53.035 ;
        RECT 253.335 52.945 253.475 55.095 ;
        RECT 254.715 53.715 254.855 55.775 ;
        RECT 256.035 55.095 256.295 55.415 ;
        RECT 259.315 55.155 259.455 58.155 ;
        RECT 259.775 57.115 259.915 61.815 ;
        RECT 260.175 61.555 260.435 61.875 ;
        RECT 262.475 61.555 262.735 61.875 ;
        RECT 262.935 61.555 263.195 61.875 ;
        RECT 269.375 61.555 269.635 61.875 ;
        RECT 262.535 61.390 262.675 61.555 ;
        RECT 262.465 61.020 262.745 61.390 ;
        RECT 262.995 59.835 263.135 61.555 ;
        RECT 263.855 60.875 264.115 61.195 ;
        RECT 262.935 59.515 263.195 59.835 ;
        RECT 263.915 59.155 264.055 60.875 ;
        RECT 269.435 59.155 269.575 61.555 ;
        RECT 263.855 58.835 264.115 59.155 ;
        RECT 269.375 58.835 269.635 59.155 ;
        RECT 263.915 58.135 264.055 58.835 ;
        RECT 269.895 58.815 270.035 63.255 ;
        RECT 269.835 58.495 270.095 58.815 ;
        RECT 263.855 57.815 264.115 58.135 ;
        RECT 260.945 57.280 262.485 57.650 ;
        RECT 270.355 57.115 270.495 71.415 ;
        RECT 275.415 69.695 275.555 71.755 ;
        RECT 270.755 69.375 271.015 69.695 ;
        RECT 275.355 69.375 275.615 69.695 ;
        RECT 270.815 67.315 270.955 69.375 ;
        RECT 273.055 69.035 273.315 69.355 ;
        RECT 273.115 67.315 273.255 69.035 ;
        RECT 270.755 66.995 271.015 67.315 ;
        RECT 273.055 66.995 273.315 67.315 ;
        RECT 270.815 63.915 270.955 66.995 ;
        RECT 272.595 66.315 272.855 66.635 ;
        RECT 272.655 64.255 272.795 66.315 ;
        RECT 273.115 65.275 273.255 66.995 ;
        RECT 275.415 66.295 275.555 69.375 ;
        RECT 275.875 67.655 276.015 80.255 ;
        RECT 276.335 72.755 276.475 81.275 ;
        RECT 276.735 80.595 276.995 80.915 ;
        RECT 276.795 77.515 276.935 80.595 ;
        RECT 278.175 80.575 278.315 91.135 ;
        RECT 279.095 89.075 279.235 96.915 ;
        RECT 279.035 88.755 279.295 89.075 ;
        RECT 279.095 86.015 279.235 88.755 ;
        RECT 279.035 85.695 279.295 86.015 ;
        RECT 278.575 80.935 278.835 81.255 ;
        RECT 278.115 80.255 278.375 80.575 ;
        RECT 278.115 77.535 278.375 77.855 ;
        RECT 276.735 77.195 276.995 77.515 ;
        RECT 278.175 76.155 278.315 77.535 ;
        RECT 278.115 75.835 278.375 76.155 ;
        RECT 278.635 75.555 278.775 80.935 ;
        RECT 279.095 78.875 279.235 85.695 ;
        RECT 279.035 78.555 279.295 78.875 ;
        RECT 276.735 75.155 276.995 75.475 ;
        RECT 278.175 75.415 278.775 75.555 ;
        RECT 276.275 72.435 276.535 72.755 ;
        RECT 276.795 72.415 276.935 75.155 ;
        RECT 277.655 73.115 277.915 73.435 ;
        RECT 277.195 72.435 277.455 72.755 ;
        RECT 276.735 72.095 276.995 72.415 ;
        RECT 277.255 69.695 277.395 72.435 ;
        RECT 277.715 71.735 277.855 73.115 ;
        RECT 277.655 71.415 277.915 71.735 ;
        RECT 278.175 70.375 278.315 75.415 ;
        RECT 278.575 74.815 278.835 75.135 ;
        RECT 278.635 73.435 278.775 74.815 ;
        RECT 278.575 73.115 278.835 73.435 ;
        RECT 279.555 73.395 279.695 105.075 ;
        RECT 281.855 104.285 281.995 105.075 ;
        RECT 281.395 104.145 281.995 104.285 ;
        RECT 280.875 101.335 281.135 101.655 ;
        RECT 279.955 96.235 280.215 96.555 ;
        RECT 280.015 95.195 280.155 96.235 ;
        RECT 279.955 94.875 280.215 95.195 ;
        RECT 280.935 94.425 281.075 101.335 ;
        RECT 280.475 94.285 281.075 94.425 ;
        RECT 280.475 81.595 280.615 94.285 ;
        RECT 280.875 93.515 281.135 93.835 ;
        RECT 280.935 91.115 281.075 93.515 ;
        RECT 280.875 90.795 281.135 91.115 ;
        RECT 280.415 81.275 280.675 81.595 ;
        RECT 280.475 80.915 280.615 81.275 ;
        RECT 280.415 80.595 280.675 80.915 ;
        RECT 280.475 80.315 280.615 80.595 ;
        RECT 280.475 80.175 281.075 80.315 ;
        RECT 281.395 80.235 281.535 104.145 ;
        RECT 281.795 98.615 282.055 98.935 ;
        RECT 281.855 92.475 281.995 98.615 ;
        RECT 282.315 97.915 282.455 109.155 ;
        RECT 283.175 107.115 283.435 107.435 ;
        RECT 282.715 106.775 282.975 107.095 ;
        RECT 282.775 106.075 282.915 106.775 ;
        RECT 283.235 106.075 283.375 107.115 ;
        RECT 282.715 105.755 282.975 106.075 ;
        RECT 283.175 105.755 283.435 106.075 ;
        RECT 282.715 101.675 282.975 101.995 ;
        RECT 282.775 100.295 282.915 101.675 ;
        RECT 282.715 99.975 282.975 100.295 ;
        RECT 282.255 97.595 282.515 97.915 ;
        RECT 282.315 95.195 282.455 97.595 ;
        RECT 282.775 96.555 282.915 99.975 ;
        RECT 283.175 99.635 283.435 99.955 ;
        RECT 282.715 96.235 282.975 96.555 ;
        RECT 283.235 95.955 283.375 99.635 ;
        RECT 283.695 99.615 283.835 109.225 ;
        RECT 285.015 105.075 285.275 105.395 ;
        RECT 285.075 104.115 285.215 105.075 ;
        RECT 285.075 103.975 285.675 104.115 ;
        RECT 285.015 103.035 285.275 103.355 ;
        RECT 284.555 100.315 284.815 100.635 ;
        RECT 283.635 99.295 283.895 99.615 ;
        RECT 284.615 98.935 284.755 100.315 ;
        RECT 285.075 99.955 285.215 103.035 ;
        RECT 285.535 100.035 285.675 103.975 ;
        RECT 285.995 102.755 286.135 109.225 ;
        RECT 286.915 105.395 287.515 105.475 ;
        RECT 286.855 105.335 287.515 105.395 ;
        RECT 286.855 105.075 287.115 105.335 ;
        RECT 285.995 102.615 286.595 102.755 ;
        RECT 285.935 101.675 286.195 101.995 ;
        RECT 285.995 100.635 286.135 101.675 ;
        RECT 285.935 100.315 286.195 100.635 ;
        RECT 285.015 99.635 285.275 99.955 ;
        RECT 285.535 99.895 286.135 100.035 ;
        RECT 285.475 99.295 285.735 99.615 ;
        RECT 284.555 98.615 284.815 98.935 ;
        RECT 285.535 96.750 285.675 99.295 ;
        RECT 285.465 96.380 285.745 96.750 ;
        RECT 282.775 95.815 283.375 95.955 ;
        RECT 284.555 95.895 284.815 96.215 ;
        RECT 285.015 95.895 285.275 96.215 ;
        RECT 282.255 94.875 282.515 95.195 ;
        RECT 282.775 94.175 282.915 95.815 ;
        RECT 283.635 94.875 283.895 95.195 ;
        RECT 283.175 94.195 283.435 94.515 ;
        RECT 282.715 93.855 282.975 94.175 ;
        RECT 281.795 92.155 282.055 92.475 ;
        RECT 281.855 91.795 281.995 92.155 ;
        RECT 283.235 91.795 283.375 94.195 ;
        RECT 281.795 91.475 282.055 91.795 ;
        RECT 283.175 91.475 283.435 91.795 ;
        RECT 282.255 90.455 282.515 90.775 ;
        RECT 281.795 86.035 282.055 86.355 ;
        RECT 281.855 80.915 281.995 86.035 ;
        RECT 281.795 80.595 282.055 80.915 ;
        RECT 280.415 79.575 280.675 79.895 ;
        RECT 280.475 75.475 280.615 79.575 ;
        RECT 280.935 75.475 281.075 80.175 ;
        RECT 281.335 79.915 281.595 80.235 ;
        RECT 280.415 75.155 280.675 75.475 ;
        RECT 280.875 75.155 281.135 75.475 ;
        RECT 280.875 74.475 281.135 74.795 ;
        RECT 279.095 73.255 279.695 73.395 ;
        RECT 278.115 70.055 278.375 70.375 ;
        RECT 277.195 69.375 277.455 69.695 ;
        RECT 275.815 67.335 276.075 67.655 ;
        RECT 277.255 66.975 277.395 69.375 ;
        RECT 277.195 66.655 277.455 66.975 ;
        RECT 275.355 65.975 275.615 66.295 ;
        RECT 273.055 64.955 273.315 65.275 ;
        RECT 272.595 63.935 272.855 64.255 ;
        RECT 270.755 63.595 271.015 63.915 ;
        RECT 275.415 61.535 275.555 65.975 ;
        RECT 277.255 64.935 277.395 66.655 ;
        RECT 277.195 64.615 277.455 64.935 ;
        RECT 277.255 61.875 277.395 64.615 ;
        RECT 277.195 61.555 277.455 61.875 ;
        RECT 278.175 61.535 278.315 70.055 ;
        RECT 278.635 70.035 278.775 73.115 ;
        RECT 278.575 69.715 278.835 70.035 ;
        RECT 279.095 68.870 279.235 73.255 ;
        RECT 279.495 69.035 279.755 69.355 ;
        RECT 279.025 68.500 279.305 68.870 ;
        RECT 279.555 67.995 279.695 69.035 ;
        RECT 279.495 67.675 279.755 67.995 ;
        RECT 279.495 66.995 279.755 67.315 ;
        RECT 279.555 66.830 279.695 66.995 ;
        RECT 279.485 66.460 279.765 66.830 ;
        RECT 279.555 64.595 279.695 66.460 ;
        RECT 279.495 64.275 279.755 64.595 ;
        RECT 279.955 64.275 280.215 64.595 ;
        RECT 279.035 62.235 279.295 62.555 ;
        RECT 275.355 61.215 275.615 61.535 ;
        RECT 278.115 61.215 278.375 61.535 ;
        RECT 272.135 60.875 272.395 61.195 ;
        RECT 272.195 58.475 272.335 60.875 ;
        RECT 279.095 59.835 279.235 62.235 ;
        RECT 279.035 59.515 279.295 59.835 ;
        RECT 272.135 58.155 272.395 58.475 ;
        RECT 274.895 58.155 275.155 58.475 ;
        RECT 279.025 58.300 279.305 58.670 ;
        RECT 274.955 57.115 275.095 58.155 ;
        RECT 279.095 58.135 279.235 58.300 ;
        RECT 279.035 57.815 279.295 58.135 ;
        RECT 259.715 56.795 259.975 57.115 ;
        RECT 270.295 56.795 270.555 57.115 ;
        RECT 274.895 56.795 275.155 57.115 ;
        RECT 264.315 56.455 264.575 56.775 ;
        RECT 262.935 56.115 263.195 56.435 ;
        RECT 261.095 55.775 261.355 56.095 ;
        RECT 255.575 54.075 255.835 54.395 ;
        RECT 254.655 53.395 254.915 53.715 ;
        RECT 254.195 52.945 254.455 53.035 ;
        RECT 253.335 52.805 254.455 52.945 ;
        RECT 250.055 52.375 250.315 52.695 ;
        RECT 251.435 52.375 251.695 52.695 ;
        RECT 252.415 52.550 252.555 52.715 ;
        RECT 251.495 50.995 251.635 52.375 ;
        RECT 252.345 52.180 252.625 52.550 ;
        RECT 252.815 51.355 253.075 51.675 ;
        RECT 252.875 50.995 253.015 51.355 ;
        RECT 249.595 50.675 249.855 50.995 ;
        RECT 251.435 50.675 251.695 50.995 ;
        RECT 252.815 50.675 253.075 50.995 ;
        RECT 247.285 50.140 247.565 50.510 ;
        RECT 246.835 49.655 247.095 49.975 ;
        RECT 249.655 49.830 249.795 50.675 ;
        RECT 245.915 48.635 246.175 48.955 ;
        RECT 245.975 45.215 246.115 48.635 ;
        RECT 245.915 44.895 246.175 45.215 ;
        RECT 246.895 42.835 247.035 49.655 ;
        RECT 249.585 49.460 249.865 49.830 ;
        RECT 251.895 46.935 252.155 47.255 ;
        RECT 251.955 45.895 252.095 46.935 ;
        RECT 252.875 46.235 253.015 50.675 ;
        RECT 252.815 45.915 253.075 46.235 ;
        RECT 251.895 45.575 252.155 45.895 ;
        RECT 251.895 44.895 252.155 45.215 ;
        RECT 251.955 43.515 252.095 44.895 ;
        RECT 251.895 43.195 252.155 43.515 ;
        RECT 246.835 42.515 247.095 42.835 ;
        RECT 249.135 41.835 249.395 42.155 ;
        RECT 253.335 42.065 253.475 52.805 ;
        RECT 254.195 52.715 254.455 52.805 ;
        RECT 253.725 50.820 254.005 51.190 ;
        RECT 253.735 50.675 253.995 50.820 ;
        RECT 254.195 50.675 254.455 50.995 ;
        RECT 254.255 48.955 254.395 50.675 ;
        RECT 254.195 48.635 254.455 48.955 ;
        RECT 254.715 48.275 254.855 53.395 ;
        RECT 255.115 52.550 255.375 52.695 ;
        RECT 255.105 52.180 255.385 52.550 ;
        RECT 255.115 50.335 255.375 50.655 ;
        RECT 254.655 47.955 254.915 48.275 ;
        RECT 255.175 43.175 255.315 50.335 ;
        RECT 255.635 44.875 255.775 54.075 ;
        RECT 256.095 53.375 256.235 55.095 ;
        RECT 259.315 55.015 259.915 55.155 ;
        RECT 257.645 54.560 259.185 54.930 ;
        RECT 256.035 53.055 256.295 53.375 ;
        RECT 256.095 51.335 256.235 53.055 ;
        RECT 259.775 53.035 259.915 55.015 ;
        RECT 261.155 54.395 261.295 55.775 ;
        RECT 261.095 54.075 261.355 54.395 ;
        RECT 259.715 52.715 259.975 53.035 ;
        RECT 256.495 52.375 256.755 52.695 ;
        RECT 256.035 51.015 256.295 51.335 ;
        RECT 256.035 50.335 256.295 50.655 ;
        RECT 256.095 48.275 256.235 50.335 ;
        RECT 256.555 48.275 256.695 52.375 ;
        RECT 256.955 50.675 257.215 50.995 ;
        RECT 256.035 47.955 256.295 48.275 ;
        RECT 256.495 47.955 256.755 48.275 ;
        RECT 256.555 45.215 256.695 47.955 ;
        RECT 256.495 44.895 256.755 45.215 ;
        RECT 255.575 44.555 255.835 44.875 ;
        RECT 257.015 43.515 257.155 50.675 ;
        RECT 257.645 49.120 259.185 49.490 ;
        RECT 257.415 47.275 257.675 47.595 ;
        RECT 257.475 45.895 257.615 47.275 ;
        RECT 259.775 47.255 259.915 52.715 ;
        RECT 260.945 51.840 262.485 52.210 ;
        RECT 262.995 51.335 263.135 56.115 ;
        RECT 263.395 53.735 263.655 54.055 ;
        RECT 262.935 51.015 263.195 51.335 ;
        RECT 262.935 49.995 263.195 50.315 ;
        RECT 260.175 49.655 260.435 49.975 ;
        RECT 259.715 46.935 259.975 47.255 ;
        RECT 257.415 45.575 257.675 45.895 ;
        RECT 260.235 45.555 260.375 49.655 ;
        RECT 260.945 46.400 262.485 46.770 ;
        RECT 260.175 45.235 260.435 45.555 ;
        RECT 257.645 43.680 259.185 44.050 ;
        RECT 256.955 43.195 257.215 43.515 ;
        RECT 255.115 42.855 255.375 43.175 ;
        RECT 262.995 42.835 263.135 49.995 ;
        RECT 263.455 48.275 263.595 53.735 ;
        RECT 263.395 47.955 263.655 48.275 ;
        RECT 263.395 46.935 263.655 47.255 ;
        RECT 263.455 44.535 263.595 46.935 ;
        RECT 264.375 45.215 264.515 56.455 ;
        RECT 276.735 56.115 276.995 56.435 ;
        RECT 267.995 53.395 268.255 53.715 ;
        RECT 267.075 51.015 267.335 51.335 ;
        RECT 266.155 49.655 266.415 49.975 ;
        RECT 266.215 47.595 266.355 49.655 ;
        RECT 266.155 47.275 266.415 47.595 ;
        RECT 264.775 45.915 265.035 46.235 ;
        RECT 264.315 44.895 264.575 45.215 ;
        RECT 263.395 44.215 263.655 44.535 ;
        RECT 262.935 42.515 263.195 42.835 ;
        RECT 263.455 42.495 263.595 44.215 ;
        RECT 263.845 44.020 264.125 44.390 ;
        RECT 263.915 43.175 264.055 44.020 ;
        RECT 264.835 43.175 264.975 45.915 ;
        RECT 265.235 45.575 265.495 45.895 ;
        RECT 263.855 42.855 264.115 43.175 ;
        RECT 264.775 42.855 265.035 43.175 ;
        RECT 263.395 42.175 263.655 42.495 ;
        RECT 253.735 42.065 253.995 42.155 ;
        RECT 260.175 42.065 260.435 42.155 ;
        RECT 253.335 41.925 253.995 42.065 ;
        RECT 253.735 41.835 253.995 41.925 ;
        RECT 259.775 41.925 260.435 42.065 ;
        RECT 248.675 40.135 248.935 40.455 ;
        RECT 248.735 39.775 248.875 40.135 ;
        RECT 248.675 39.630 248.935 39.775 ;
        RECT 248.215 39.115 248.475 39.435 ;
        RECT 248.665 39.260 248.945 39.630 ;
        RECT 248.275 38.075 248.415 39.115 ;
        RECT 248.215 37.755 248.475 38.075 ;
        RECT 249.195 32.635 249.335 41.835 ;
        RECT 254.655 41.495 254.915 41.815 ;
        RECT 256.035 41.495 256.295 41.815 ;
        RECT 249.595 40.475 249.855 40.795 ;
        RECT 249.655 38.075 249.795 40.475 ;
        RECT 253.275 39.455 253.535 39.775 ;
        RECT 249.595 37.755 249.855 38.075 ;
        RECT 253.335 35.355 253.475 39.455 ;
        RECT 253.275 35.035 253.535 35.355 ;
        RECT 249.135 32.315 249.395 32.635 ;
        RECT 245.455 31.295 245.715 31.615 ;
        RECT 254.715 31.275 254.855 41.495 ;
        RECT 256.095 38.075 256.235 41.495 ;
        RECT 258.795 40.475 259.055 40.795 ;
        RECT 258.335 39.685 258.595 39.775 ;
        RECT 258.855 39.685 258.995 40.475 ;
        RECT 259.775 39.775 259.915 41.925 ;
        RECT 260.175 41.835 260.435 41.925 ;
        RECT 264.835 41.815 264.975 42.855 ;
        RECT 265.295 42.495 265.435 45.575 ;
        RECT 266.215 45.555 266.355 47.275 ;
        RECT 266.155 45.235 266.415 45.555 ;
        RECT 267.135 42.835 267.275 51.015 ;
        RECT 268.055 50.995 268.195 53.395 ;
        RECT 270.755 53.055 271.015 53.375 ;
        RECT 267.995 50.675 268.255 50.995 ;
        RECT 269.375 50.335 269.635 50.655 ;
        RECT 267.995 49.995 268.255 50.315 ;
        RECT 267.535 47.615 267.795 47.935 ;
        RECT 267.595 46.235 267.735 47.615 ;
        RECT 267.535 45.915 267.795 46.235 ;
        RECT 268.055 45.555 268.195 49.995 ;
        RECT 269.435 48.955 269.575 50.335 ;
        RECT 269.375 48.635 269.635 48.955 ;
        RECT 269.375 47.275 269.635 47.595 ;
        RECT 268.455 45.915 268.715 46.235 ;
        RECT 267.995 45.235 268.255 45.555 ;
        RECT 267.075 42.745 267.335 42.835 ;
        RECT 266.675 42.605 267.335 42.745 ;
        RECT 265.235 42.175 265.495 42.495 ;
        RECT 264.775 41.495 265.035 41.815 ;
        RECT 260.945 40.960 262.485 41.330 ;
        RECT 265.295 40.795 265.435 42.175 ;
        RECT 265.235 40.475 265.495 40.795 ;
        RECT 260.175 39.795 260.435 40.115 ;
        RECT 258.335 39.545 258.995 39.685 ;
        RECT 258.335 39.455 258.595 39.545 ;
        RECT 259.715 39.455 259.975 39.775 ;
        RECT 256.955 39.115 257.215 39.435 ;
        RECT 256.035 37.755 256.295 38.075 ;
        RECT 256.095 31.955 256.235 37.755 ;
        RECT 257.015 35.015 257.155 39.115 ;
        RECT 257.645 38.240 259.185 38.610 ;
        RECT 257.415 36.735 257.675 37.055 ;
        RECT 257.475 35.015 257.615 36.735 ;
        RECT 256.955 34.695 257.215 35.015 ;
        RECT 257.415 34.695 257.675 35.015 ;
        RECT 257.475 34.335 257.615 34.695 ;
        RECT 257.415 34.015 257.675 34.335 ;
        RECT 259.775 33.655 259.915 39.455 ;
        RECT 260.235 38.075 260.375 39.795 ;
        RECT 260.175 37.755 260.435 38.075 ;
        RECT 259.715 33.335 259.975 33.655 ;
        RECT 257.645 32.800 259.185 33.170 ;
        RECT 260.235 32.635 260.375 37.755 ;
        RECT 266.675 37.395 266.815 42.605 ;
        RECT 267.075 42.515 267.335 42.605 ;
        RECT 268.515 42.155 268.655 45.915 ;
        RECT 268.915 45.465 269.175 45.555 ;
        RECT 269.435 45.465 269.575 47.275 ;
        RECT 268.915 45.325 269.575 45.465 ;
        RECT 268.915 45.235 269.175 45.325 ;
        RECT 269.435 43.515 269.575 45.325 ;
        RECT 270.815 44.875 270.955 53.055 ;
        RECT 276.795 51.335 276.935 56.115 ;
        RECT 279.555 53.375 279.695 64.275 ;
        RECT 280.015 62.555 280.155 64.275 ;
        RECT 280.935 63.915 281.075 74.475 ;
        RECT 281.795 68.695 282.055 69.015 ;
        RECT 281.855 67.995 281.995 68.695 ;
        RECT 281.795 67.675 282.055 67.995 ;
        RECT 280.875 63.595 281.135 63.915 ;
        RECT 281.795 63.255 282.055 63.575 ;
        RECT 279.955 62.235 280.215 62.555 ;
        RECT 280.015 59.155 280.155 62.235 ;
        RECT 281.855 62.215 281.995 63.255 ;
        RECT 281.795 61.895 282.055 62.215 ;
        RECT 282.315 61.390 282.455 90.455 ;
        RECT 283.695 83.975 283.835 94.875 ;
        RECT 284.615 94.515 284.755 95.895 ;
        RECT 284.555 94.195 284.815 94.515 ;
        RECT 284.095 93.175 284.355 93.495 ;
        RECT 284.155 86.015 284.295 93.175 ;
        RECT 284.615 91.455 284.755 94.195 ;
        RECT 284.555 91.135 284.815 91.455 ;
        RECT 284.095 85.695 284.355 86.015 ;
        RECT 283.635 83.655 283.895 83.975 ;
        RECT 284.155 81.255 284.295 85.695 ;
        RECT 284.095 80.935 284.355 81.255 ;
        RECT 282.715 80.595 282.975 80.915 ;
        RECT 283.175 80.595 283.435 80.915 ;
        RECT 282.775 76.155 282.915 80.595 ;
        RECT 282.715 75.835 282.975 76.155 ;
        RECT 283.235 72.415 283.375 80.595 ;
        RECT 284.095 79.915 284.355 80.235 ;
        RECT 283.635 77.875 283.895 78.195 ;
        RECT 283.695 73.095 283.835 77.875 ;
        RECT 283.635 72.775 283.895 73.095 ;
        RECT 283.175 72.095 283.435 72.415 ;
        RECT 283.235 66.975 283.375 72.095 ;
        RECT 283.695 69.355 283.835 72.775 ;
        RECT 283.635 69.035 283.895 69.355 ;
        RECT 284.155 67.995 284.295 79.915 ;
        RECT 284.555 72.775 284.815 73.095 ;
        RECT 284.615 72.415 284.755 72.775 ;
        RECT 284.555 72.095 284.815 72.415 ;
        RECT 284.095 67.675 284.355 67.995 ;
        RECT 283.175 66.655 283.435 66.975 ;
        RECT 284.155 63.575 284.295 67.675 ;
        RECT 285.075 63.995 285.215 95.895 ;
        RECT 285.535 90.630 285.675 96.380 ;
        RECT 285.465 90.260 285.745 90.630 ;
        RECT 285.475 88.755 285.735 89.075 ;
        RECT 285.535 80.145 285.675 88.755 ;
        RECT 285.995 83.830 286.135 99.895 ;
        RECT 286.455 97.915 286.595 102.615 ;
        RECT 286.395 97.595 286.655 97.915 ;
        RECT 286.855 96.915 287.115 97.235 ;
        RECT 286.915 94.515 287.055 96.915 ;
        RECT 286.855 94.195 287.115 94.515 ;
        RECT 286.915 89.755 287.055 94.195 ;
        RECT 287.375 93.915 287.515 105.335 ;
        RECT 288.295 100.635 288.435 109.225 ;
        RECT 289.155 108.815 289.415 109.135 ;
        RECT 289.215 107.435 289.355 108.815 ;
        RECT 289.155 107.115 289.415 107.435 ;
        RECT 289.215 105.395 289.355 107.115 ;
        RECT 289.155 105.075 289.415 105.395 ;
        RECT 288.695 104.735 288.955 105.055 ;
        RECT 288.755 102.675 288.895 104.735 ;
        RECT 290.595 104.375 290.735 109.225 ;
        RECT 292.375 108.475 292.635 108.795 ;
        RECT 292.435 105.395 292.575 108.475 ;
        RECT 292.895 107.095 293.035 109.225 ;
        RECT 292.835 106.775 293.095 107.095 ;
        RECT 292.375 105.075 292.635 105.395 ;
        RECT 294.215 105.075 294.475 105.395 ;
        RECT 291.915 104.395 292.175 104.715 ;
        RECT 290.535 104.055 290.795 104.375 ;
        RECT 291.975 103.355 292.115 104.395 ;
        RECT 291.915 103.035 292.175 103.355 ;
        RECT 288.695 102.355 288.955 102.675 ;
        RECT 290.075 101.675 290.335 101.995 ;
        RECT 290.535 101.675 290.795 101.995 ;
        RECT 288.235 100.315 288.495 100.635 ;
        RECT 288.235 99.635 288.495 99.955 ;
        RECT 287.775 95.895 288.035 96.215 ;
        RECT 287.835 94.855 287.975 95.895 ;
        RECT 288.295 95.195 288.435 99.635 ;
        RECT 290.135 97.915 290.275 101.675 ;
        RECT 290.595 100.295 290.735 101.675 ;
        RECT 290.535 99.975 290.795 100.295 ;
        RECT 290.075 97.595 290.335 97.915 ;
        RECT 290.595 96.555 290.735 99.975 ;
        RECT 291.455 99.635 291.715 99.955 ;
        RECT 290.535 96.235 290.795 96.555 ;
        RECT 288.235 94.875 288.495 95.195 ;
        RECT 287.775 94.535 288.035 94.855 ;
        RECT 288.695 94.595 288.955 94.855 ;
        RECT 288.295 94.535 288.955 94.595 ;
        RECT 288.295 94.455 288.895 94.535 ;
        RECT 288.295 93.915 288.435 94.455 ;
        RECT 287.375 93.775 288.435 93.915 ;
        RECT 287.315 91.475 287.575 91.795 ;
        RECT 286.855 89.435 287.115 89.755 ;
        RECT 287.375 88.735 287.515 91.475 ;
        RECT 287.315 88.415 287.575 88.735 ;
        RECT 286.395 85.695 286.655 86.015 ;
        RECT 285.925 83.460 286.205 83.830 ;
        RECT 286.455 83.635 286.595 85.695 ;
        RECT 288.295 85.335 288.435 93.775 ;
        RECT 290.075 91.815 290.335 92.135 ;
        RECT 288.685 90.940 288.965 91.310 ;
        RECT 288.755 89.075 288.895 90.940 ;
        RECT 288.695 88.755 288.955 89.075 ;
        RECT 290.135 85.675 290.275 91.815 ;
        RECT 290.535 90.795 290.795 91.115 ;
        RECT 290.595 89.755 290.735 90.795 ;
        RECT 290.535 89.435 290.795 89.755 ;
        RECT 290.075 85.355 290.335 85.675 ;
        RECT 288.235 85.015 288.495 85.335 ;
        RECT 286.395 83.315 286.655 83.635 ;
        RECT 286.455 80.915 286.595 83.315 ;
        RECT 286.395 80.595 286.655 80.915 ;
        RECT 285.935 80.145 286.195 80.235 ;
        RECT 285.535 80.005 286.195 80.145 ;
        RECT 285.935 79.915 286.195 80.005 ;
        RECT 285.995 78.535 286.135 79.915 ;
        RECT 285.935 78.215 286.195 78.535 ;
        RECT 285.475 75.495 285.735 75.815 ;
        RECT 285.535 74.455 285.675 75.495 ;
        RECT 285.475 74.135 285.735 74.455 ;
        RECT 285.475 70.055 285.735 70.375 ;
        RECT 284.615 63.855 285.215 63.995 ;
        RECT 284.095 63.255 284.355 63.575 ;
        RECT 284.155 62.070 284.295 63.255 ;
        RECT 284.085 61.700 284.365 62.070 ;
        RECT 282.245 61.020 282.525 61.390 ;
        RECT 283.635 60.535 283.895 60.855 ;
        RECT 279.955 58.835 280.215 59.155 ;
        RECT 280.015 53.715 280.155 58.835 ;
        RECT 283.695 58.815 283.835 60.535 ;
        RECT 284.615 59.350 284.755 63.855 ;
        RECT 285.015 63.255 285.275 63.575 ;
        RECT 284.545 58.980 284.825 59.350 ;
        RECT 285.075 59.155 285.215 63.255 ;
        RECT 283.635 58.495 283.895 58.815 ;
        RECT 282.255 57.815 282.515 58.135 ;
        RECT 282.315 56.775 282.455 57.815 ;
        RECT 283.695 56.775 283.835 58.495 ;
        RECT 282.255 56.455 282.515 56.775 ;
        RECT 283.635 56.455 283.895 56.775 ;
        RECT 283.695 56.095 283.835 56.455 ;
        RECT 283.635 55.775 283.895 56.095 ;
        RECT 279.955 53.395 280.215 53.715 ;
        RECT 279.495 53.055 279.755 53.375 ;
        RECT 278.575 52.715 278.835 53.035 ;
        RECT 276.735 51.015 276.995 51.335 ;
        RECT 277.195 49.655 277.455 49.975 ;
        RECT 277.655 49.655 277.915 49.975 ;
        RECT 277.255 48.275 277.395 49.655 ;
        RECT 277.195 47.955 277.455 48.275 ;
        RECT 277.715 47.595 277.855 49.655 ;
        RECT 278.635 48.955 278.775 52.715 ;
        RECT 280.415 52.375 280.675 52.695 ;
        RECT 280.475 51.335 280.615 52.375 ;
        RECT 283.695 51.675 283.835 55.775 ;
        RECT 284.615 52.695 284.755 58.980 ;
        RECT 285.015 58.835 285.275 59.155 ;
        RECT 285.535 58.475 285.675 70.055 ;
        RECT 285.475 58.155 285.735 58.475 ;
        RECT 285.995 55.415 286.135 78.215 ;
        RECT 286.455 72.755 286.595 80.595 ;
        RECT 290.535 80.255 290.795 80.575 ;
        RECT 291.515 80.430 291.655 99.635 ;
        RECT 291.975 96.215 292.115 103.035 ;
        RECT 293.295 102.355 293.555 102.675 ;
        RECT 293.355 97.235 293.495 102.355 ;
        RECT 294.275 101.655 294.415 105.075 ;
        RECT 295.195 103.015 295.335 109.225 ;
        RECT 297.495 106.075 297.635 109.225 ;
        RECT 297.435 105.755 297.695 106.075 ;
        RECT 299.275 105.415 299.535 105.735 ;
        RECT 296.055 104.735 296.315 105.055 ;
        RECT 296.115 103.355 296.255 104.735 ;
        RECT 297.645 103.520 299.185 103.890 ;
        RECT 295.595 103.035 295.855 103.355 ;
        RECT 296.055 103.035 296.315 103.355 ;
        RECT 295.135 102.695 295.395 103.015 ;
        RECT 295.655 102.755 295.795 103.035 ;
        RECT 295.655 102.615 297.635 102.755 ;
        RECT 296.515 102.015 296.775 102.335 ;
        RECT 294.215 101.335 294.475 101.655 ;
        RECT 294.675 99.975 294.935 100.295 ;
        RECT 292.375 96.915 292.635 97.235 ;
        RECT 293.295 96.915 293.555 97.235 ;
        RECT 291.915 95.895 292.175 96.215 ;
        RECT 291.975 91.455 292.115 95.895 ;
        RECT 292.435 91.455 292.575 96.915 ;
        RECT 293.355 94.175 293.495 96.915 ;
        RECT 294.735 96.895 294.875 99.975 ;
        RECT 294.675 96.805 294.935 96.895 ;
        RECT 294.675 96.665 295.335 96.805 ;
        RECT 294.675 96.575 294.935 96.665 ;
        RECT 295.195 94.175 295.335 96.665 ;
        RECT 293.295 93.855 293.555 94.175 ;
        RECT 295.135 93.855 295.395 94.175 ;
        RECT 291.915 91.135 292.175 91.455 ;
        RECT 292.375 91.135 292.635 91.455 ;
        RECT 294.675 91.365 294.935 91.455 ;
        RECT 295.195 91.365 295.335 93.855 ;
        RECT 294.675 91.225 295.335 91.365 ;
        RECT 294.675 91.135 294.935 91.225 ;
        RECT 291.915 90.455 292.175 90.775 ;
        RECT 292.375 90.455 292.635 90.775 ;
        RECT 291.975 88.395 292.115 90.455 ;
        RECT 292.435 89.075 292.575 90.455 ;
        RECT 292.375 88.755 292.635 89.075 ;
        RECT 295.195 88.735 295.335 91.225 ;
        RECT 295.135 88.415 295.395 88.735 ;
        RECT 291.915 88.075 292.175 88.395 ;
        RECT 291.975 87.035 292.115 88.075 ;
        RECT 291.915 86.715 292.175 87.035 ;
        RECT 295.195 86.355 295.335 88.415 ;
        RECT 296.575 87.035 296.715 102.015 ;
        RECT 296.975 101.675 297.235 101.995 ;
        RECT 297.035 98.935 297.175 101.675 ;
        RECT 297.495 101.655 297.635 102.615 ;
        RECT 297.435 101.335 297.695 101.655 ;
        RECT 297.895 101.335 298.155 101.655 ;
        RECT 297.955 99.615 298.095 101.335 ;
        RECT 298.355 100.315 298.615 100.635 ;
        RECT 298.415 99.615 298.555 100.315 ;
        RECT 297.895 99.295 298.155 99.615 ;
        RECT 298.355 99.295 298.615 99.615 ;
        RECT 296.975 98.615 297.235 98.935 ;
        RECT 297.645 98.080 299.185 98.450 ;
        RECT 299.335 96.215 299.475 105.415 ;
        RECT 299.795 101.395 299.935 109.225 ;
        RECT 302.095 107.515 302.235 109.225 ;
        RECT 302.095 107.375 303.155 107.515 ;
        RECT 300.945 106.240 302.485 106.610 ;
        RECT 299.795 101.255 300.395 101.395 ;
        RECT 299.735 100.315 299.995 100.635 ;
        RECT 299.275 96.125 299.535 96.215 ;
        RECT 298.875 95.985 299.535 96.125 ;
        RECT 298.875 95.195 299.015 95.985 ;
        RECT 299.275 95.895 299.535 95.985 ;
        RECT 298.815 94.875 299.075 95.195 ;
        RECT 299.275 94.875 299.535 95.195 ;
        RECT 298.875 93.495 299.015 94.875 ;
        RECT 298.815 93.175 299.075 93.495 ;
        RECT 297.645 92.640 299.185 93.010 ;
        RECT 297.645 87.200 299.185 87.570 ;
        RECT 296.515 86.715 296.775 87.035 ;
        RECT 295.135 86.035 295.395 86.355 ;
        RECT 296.055 86.035 296.315 86.355 ;
        RECT 296.115 83.295 296.255 86.035 ;
        RECT 296.975 85.355 297.235 85.675 ;
        RECT 294.215 82.975 294.475 83.295 ;
        RECT 296.055 82.975 296.315 83.295 ;
        RECT 294.275 80.575 294.415 82.975 ;
        RECT 286.855 77.875 287.115 78.195 ;
        RECT 286.915 74.795 287.055 77.875 ;
        RECT 290.595 77.855 290.735 80.255 ;
        RECT 291.445 80.060 291.725 80.430 ;
        RECT 294.215 80.255 294.475 80.575 ;
        RECT 290.535 77.535 290.795 77.855 ;
        RECT 286.855 74.475 287.115 74.795 ;
        RECT 290.595 73.435 290.735 77.535 ;
        RECT 290.995 75.155 291.255 75.475 ;
        RECT 290.535 73.115 290.795 73.435 ;
        RECT 290.075 72.835 290.335 73.095 ;
        RECT 288.755 72.775 290.335 72.835 ;
        RECT 288.755 72.755 290.275 72.775 ;
        RECT 286.395 72.435 286.655 72.755 ;
        RECT 288.695 72.695 290.275 72.755 ;
        RECT 288.695 72.435 288.955 72.695 ;
        RECT 288.755 70.375 288.895 72.435 ;
        RECT 290.595 72.415 290.735 73.115 ;
        RECT 290.535 72.095 290.795 72.415 ;
        RECT 290.075 71.415 290.335 71.735 ;
        RECT 288.695 70.055 288.955 70.375 ;
        RECT 290.135 67.995 290.275 71.415 ;
        RECT 290.595 70.035 290.735 72.095 ;
        RECT 291.055 70.715 291.195 75.155 ;
        RECT 290.995 70.395 291.255 70.715 ;
        RECT 290.535 69.715 290.795 70.035 ;
        RECT 291.515 69.945 291.655 80.060 ;
        RECT 295.595 79.915 295.855 80.235 ;
        RECT 295.655 76.155 295.795 79.915 ;
        RECT 295.595 75.835 295.855 76.155 ;
        RECT 296.115 75.475 296.255 82.975 ;
        RECT 297.035 82.615 297.175 85.355 ;
        RECT 297.895 85.015 298.155 85.335 ;
        RECT 297.955 84.315 298.095 85.015 ;
        RECT 297.895 83.995 298.155 84.315 ;
        RECT 296.975 82.295 297.235 82.615 ;
        RECT 297.035 79.895 297.175 82.295 ;
        RECT 297.645 81.760 299.185 82.130 ;
        RECT 296.975 79.575 297.235 79.895 ;
        RECT 296.515 76.855 296.775 77.175 ;
        RECT 296.055 75.155 296.315 75.475 ;
        RECT 296.575 74.875 296.715 76.855 ;
        RECT 297.645 76.320 299.185 76.690 ;
        RECT 299.335 75.555 299.475 94.875 ;
        RECT 296.975 75.155 297.235 75.475 ;
        RECT 298.875 75.415 299.475 75.555 ;
        RECT 296.115 74.735 296.715 74.875 ;
        RECT 291.915 74.135 292.175 74.455 ;
        RECT 291.975 73.095 292.115 74.135 ;
        RECT 291.915 72.775 292.175 73.095 ;
        RECT 294.675 70.395 294.935 70.715 ;
        RECT 291.055 69.805 291.655 69.945 ;
        RECT 290.075 67.675 290.335 67.995 ;
        RECT 287.765 64.420 288.045 64.790 ;
        RECT 287.835 63.575 287.975 64.420 ;
        RECT 289.615 63.935 289.875 64.255 ;
        RECT 288.235 63.595 288.495 63.915 ;
        RECT 287.775 63.255 288.035 63.575 ;
        RECT 288.295 62.555 288.435 63.595 ;
        RECT 288.235 62.235 288.495 62.555 ;
        RECT 287.315 61.555 287.575 61.875 ;
        RECT 287.375 58.475 287.515 61.555 ;
        RECT 286.395 58.155 286.655 58.475 ;
        RECT 287.315 58.155 287.575 58.475 ;
        RECT 285.935 55.095 286.195 55.415 ;
        RECT 284.555 52.375 284.815 52.695 ;
        RECT 283.635 51.355 283.895 51.675 ;
        RECT 280.415 51.015 280.675 51.335 ;
        RECT 286.455 50.655 286.595 58.155 ;
        RECT 289.675 56.775 289.815 63.935 ;
        RECT 291.055 63.915 291.195 69.805 ;
        RECT 291.455 69.035 291.715 69.355 ;
        RECT 291.515 67.995 291.655 69.035 ;
        RECT 293.295 68.870 293.555 69.015 ;
        RECT 293.285 68.500 293.565 68.870 ;
        RECT 293.355 67.995 293.495 68.500 ;
        RECT 291.455 67.675 291.715 67.995 ;
        RECT 293.295 67.675 293.555 67.995 ;
        RECT 294.735 66.975 294.875 70.395 ;
        RECT 293.755 66.830 294.015 66.975 ;
        RECT 293.745 66.460 294.025 66.830 ;
        RECT 294.675 66.655 294.935 66.975 ;
        RECT 295.135 66.315 295.395 66.635 ;
        RECT 290.995 63.595 291.255 63.915 ;
        RECT 291.055 61.535 291.195 63.595 ;
        RECT 292.375 63.255 292.635 63.575 ;
        RECT 290.995 61.215 291.255 61.535 ;
        RECT 292.435 59.495 292.575 63.255 ;
        RECT 295.195 61.535 295.335 66.315 ;
        RECT 295.595 63.595 295.855 63.915 ;
        RECT 295.135 61.215 295.395 61.535 ;
        RECT 295.655 61.195 295.795 63.595 ;
        RECT 296.115 62.555 296.255 74.735 ;
        RECT 297.035 72.415 297.175 75.155 ;
        RECT 298.875 73.395 299.015 75.415 ;
        RECT 298.875 73.255 299.475 73.395 ;
        RECT 296.975 72.095 297.235 72.415 ;
        RECT 296.505 69.860 296.785 70.230 ;
        RECT 296.575 67.995 296.715 69.860 ;
        RECT 296.515 67.675 296.775 67.995 ;
        RECT 296.575 62.555 296.715 67.675 ;
        RECT 297.035 67.315 297.175 72.095 ;
        RECT 297.645 70.880 299.185 71.250 ;
        RECT 296.975 66.995 297.235 67.315 ;
        RECT 299.335 66.715 299.475 73.255 ;
        RECT 299.795 68.190 299.935 100.315 ;
        RECT 300.255 93.915 300.395 101.255 ;
        RECT 300.945 100.800 302.485 101.170 ;
        RECT 303.015 100.635 303.155 107.375 ;
        RECT 303.415 107.115 303.675 107.435 ;
        RECT 303.475 104.375 303.615 107.115 ;
        RECT 303.875 104.735 304.135 105.055 ;
        RECT 303.415 104.055 303.675 104.375 ;
        RECT 303.475 102.335 303.615 104.055 ;
        RECT 303.415 102.015 303.675 102.335 ;
        RECT 302.955 100.315 303.215 100.635 ;
        RECT 302.955 99.635 303.215 99.955 ;
        RECT 300.945 95.360 302.485 95.730 ;
        RECT 303.015 95.105 303.155 99.635 ;
        RECT 302.555 94.965 303.155 95.105 ;
        RECT 300.255 93.775 301.315 93.915 ;
        RECT 300.195 93.175 300.455 93.495 ;
        RECT 300.255 89.415 300.395 93.175 ;
        RECT 301.175 92.475 301.315 93.775 ;
        RECT 301.575 93.175 301.835 93.495 ;
        RECT 301.115 92.155 301.375 92.475 ;
        RECT 301.635 91.455 301.775 93.175 ;
        RECT 301.575 91.135 301.835 91.455 ;
        RECT 302.555 91.115 302.695 94.965 ;
        RECT 303.935 93.495 304.075 104.735 ;
        RECT 304.395 100.635 304.535 109.225 ;
        RECT 304.795 108.135 305.055 108.455 ;
        RECT 304.855 101.995 304.995 108.135 ;
        RECT 304.795 101.675 305.055 101.995 ;
        RECT 304.335 100.315 304.595 100.635 ;
        RECT 302.955 93.175 303.215 93.495 ;
        RECT 303.875 93.175 304.135 93.495 ;
        RECT 303.015 92.135 303.155 93.175 ;
        RECT 302.955 91.815 303.215 92.135 ;
        RECT 302.495 90.795 302.755 91.115 ;
        RECT 303.015 90.775 303.155 91.815 ;
        RECT 303.865 91.620 304.145 91.990 ;
        RECT 303.935 91.455 304.075 91.620 ;
        RECT 303.875 91.135 304.135 91.455 ;
        RECT 302.955 90.455 303.215 90.775 ;
        RECT 300.945 89.920 302.485 90.290 ;
        RECT 303.935 89.755 304.075 91.135 ;
        RECT 304.335 90.795 304.595 91.115 ;
        RECT 303.875 89.435 304.135 89.755 ;
        RECT 300.195 89.095 300.455 89.415 ;
        RECT 304.395 89.155 304.535 90.795 ;
        RECT 300.255 88.055 300.395 89.095 ;
        RECT 302.955 88.755 303.215 89.075 ;
        RECT 303.935 89.015 304.535 89.155 ;
        RECT 300.195 87.735 300.455 88.055 ;
        RECT 300.255 86.015 300.395 87.735 ;
        RECT 300.195 85.695 300.455 86.015 ;
        RECT 300.195 85.015 300.455 85.335 ;
        RECT 300.255 71.735 300.395 85.015 ;
        RECT 300.945 84.480 302.485 84.850 ;
        RECT 303.015 83.975 303.155 88.755 ;
        RECT 302.955 83.715 303.215 83.975 ;
        RECT 303.935 83.715 304.075 89.015 ;
        RECT 304.335 88.415 304.595 88.735 ;
        RECT 304.395 87.035 304.535 88.415 ;
        RECT 304.335 86.715 304.595 87.035 ;
        RECT 304.855 86.355 304.995 101.675 ;
        RECT 306.175 101.335 306.435 101.655 ;
        RECT 305.715 99.635 305.975 99.955 ;
        RECT 305.255 99.295 305.515 99.615 ;
        RECT 304.795 86.035 305.055 86.355 ;
        RECT 304.795 83.830 305.055 83.975 ;
        RECT 302.555 83.655 303.215 83.715 ;
        RECT 302.555 83.575 303.155 83.655 ;
        RECT 303.475 83.575 304.075 83.715 ;
        RECT 302.555 80.235 302.695 83.575 ;
        RECT 302.955 82.635 303.215 82.955 ;
        RECT 302.495 79.915 302.755 80.235 ;
        RECT 300.945 79.040 302.485 79.410 ;
        RECT 300.945 73.600 302.485 73.970 ;
        RECT 303.015 73.435 303.155 82.635 ;
        RECT 302.955 73.115 303.215 73.435 ;
        RECT 301.115 72.775 301.375 73.095 ;
        RECT 301.175 71.735 301.315 72.775 ;
        RECT 303.475 72.075 303.615 83.575 ;
        RECT 304.785 83.460 305.065 83.830 ;
        RECT 303.875 79.915 304.135 80.235 ;
        RECT 304.795 79.915 305.055 80.235 ;
        RECT 303.935 74.455 304.075 79.915 ;
        RECT 304.855 76.155 304.995 79.915 ;
        RECT 304.795 75.835 305.055 76.155 ;
        RECT 304.335 74.475 304.595 74.795 ;
        RECT 303.875 74.135 304.135 74.455 ;
        RECT 303.415 71.755 303.675 72.075 ;
        RECT 300.195 71.415 300.455 71.735 ;
        RECT 301.115 71.415 301.375 71.735 ;
        RECT 300.255 69.695 300.395 71.415 ;
        RECT 300.195 69.375 300.455 69.695 ;
        RECT 301.175 69.355 301.315 71.415 ;
        RECT 303.475 69.695 303.615 71.755 ;
        RECT 303.935 71.735 304.075 74.135 ;
        RECT 303.875 71.415 304.135 71.735 ;
        RECT 304.395 70.715 304.535 74.475 ;
        RECT 304.335 70.395 304.595 70.715 ;
        RECT 303.875 69.715 304.135 70.035 ;
        RECT 303.415 69.375 303.675 69.695 ;
        RECT 301.115 69.035 301.375 69.355 ;
        RECT 299.725 68.075 300.005 68.190 ;
        RECT 300.945 68.160 302.485 68.530 ;
        RECT 299.725 67.935 300.395 68.075 ;
        RECT 299.725 67.820 300.005 67.935 ;
        RECT 300.255 67.395 300.395 67.935 ;
        RECT 300.255 67.255 300.855 67.395 ;
        RECT 303.415 67.335 303.675 67.655 ;
        RECT 299.335 66.575 299.935 66.715 ;
        RECT 300.195 66.655 300.455 66.975 ;
        RECT 299.275 65.975 299.535 66.295 ;
        RECT 297.645 65.440 299.185 65.810 ;
        RECT 298.815 63.595 299.075 63.915 ;
        RECT 296.055 62.235 296.315 62.555 ;
        RECT 296.515 62.235 296.775 62.555 ;
        RECT 298.875 61.275 299.015 63.595 ;
        RECT 299.335 62.555 299.475 65.975 ;
        RECT 299.275 62.235 299.535 62.555 ;
        RECT 295.595 60.875 295.855 61.195 ;
        RECT 298.875 61.135 299.475 61.275 ;
        RECT 297.645 60.000 299.185 60.370 ;
        RECT 292.375 59.175 292.635 59.495 ;
        RECT 299.335 59.155 299.475 61.135 ;
        RECT 299.795 59.915 299.935 66.575 ;
        RECT 300.255 62.555 300.395 66.655 ;
        RECT 300.715 65.275 300.855 67.255 ;
        RECT 300.655 64.955 300.915 65.275 ;
        RECT 302.955 64.955 303.215 65.275 ;
        RECT 300.945 62.720 302.485 63.090 ;
        RECT 300.195 62.235 300.455 62.555 ;
        RECT 303.015 62.215 303.155 64.955 ;
        RECT 302.955 61.895 303.215 62.215 ;
        RECT 302.035 60.535 302.295 60.855 ;
        RECT 299.795 59.775 300.395 59.915 ;
        RECT 299.275 58.835 299.535 59.155 ;
        RECT 299.735 58.835 299.995 59.155 ;
        RECT 299.335 57.115 299.475 58.835 ;
        RECT 299.275 56.795 299.535 57.115 ;
        RECT 289.615 56.455 289.875 56.775 ;
        RECT 287.315 55.775 287.575 56.095 ;
        RECT 287.375 53.375 287.515 55.775 ;
        RECT 297.645 54.560 299.185 54.930 ;
        RECT 299.335 54.395 299.475 56.795 ;
        RECT 299.795 56.435 299.935 58.835 ;
        RECT 299.735 56.115 299.995 56.435 ;
        RECT 299.275 54.075 299.535 54.395 ;
        RECT 290.535 53.735 290.795 54.055 ;
        RECT 287.315 53.055 287.575 53.375 ;
        RECT 283.635 50.335 283.895 50.655 ;
        RECT 286.395 50.335 286.655 50.655 ;
        RECT 278.575 48.635 278.835 48.955 ;
        RECT 277.655 47.275 277.915 47.595 ;
        RECT 274.435 46.935 274.695 47.255 ;
        RECT 274.495 46.235 274.635 46.935 ;
        RECT 274.435 45.915 274.695 46.235 ;
        RECT 278.635 45.895 278.775 48.635 ;
        RECT 283.695 47.595 283.835 50.335 ;
        RECT 287.375 48.275 287.515 53.055 ;
        RECT 287.775 52.375 288.035 52.695 ;
        RECT 287.835 50.655 287.975 52.375 ;
        RECT 287.775 50.335 288.035 50.655 ;
        RECT 287.315 47.955 287.575 48.275 ;
        RECT 289.615 47.955 289.875 48.275 ;
        RECT 283.635 47.275 283.895 47.595 ;
        RECT 285.935 47.275 286.195 47.595 ;
        RECT 285.995 46.235 286.135 47.275 ;
        RECT 285.935 45.915 286.195 46.235 ;
        RECT 278.575 45.575 278.835 45.895 ;
        RECT 272.135 45.235 272.395 45.555 ;
        RECT 270.755 44.555 271.015 44.875 ;
        RECT 271.675 44.390 271.935 44.535 ;
        RECT 271.665 44.020 271.945 44.390 ;
        RECT 272.195 43.515 272.335 45.235 ;
        RECT 289.155 44.215 289.415 44.535 ;
        RECT 269.375 43.195 269.635 43.515 ;
        RECT 272.135 43.195 272.395 43.515 ;
        RECT 267.075 41.835 267.335 42.155 ;
        RECT 268.455 42.065 268.715 42.155 ;
        RECT 268.455 41.925 269.115 42.065 ;
        RECT 268.455 41.835 268.715 41.925 ;
        RECT 263.855 37.075 264.115 37.395 ;
        RECT 266.615 37.075 266.875 37.395 ;
        RECT 260.945 35.520 262.485 35.890 ;
        RECT 263.915 35.355 264.055 37.075 ;
        RECT 267.135 36.715 267.275 41.835 ;
        RECT 267.535 39.455 267.795 39.775 ;
        RECT 264.775 36.395 265.035 36.715 ;
        RECT 267.075 36.395 267.335 36.715 ;
        RECT 263.855 35.035 264.115 35.355 ;
        RECT 260.635 33.335 260.895 33.655 ;
        RECT 260.175 32.315 260.435 32.635 ;
        RECT 256.035 31.635 256.295 31.955 ;
        RECT 260.695 31.615 260.835 33.335 ;
        RECT 264.835 32.295 264.975 36.395 ;
        RECT 265.235 36.055 265.495 36.375 ;
        RECT 265.295 34.675 265.435 36.055 ;
        RECT 265.235 34.355 265.495 34.675 ;
        RECT 267.595 34.335 267.735 39.455 ;
        RECT 268.455 37.755 268.715 38.075 ;
        RECT 268.515 34.675 268.655 37.755 ;
        RECT 268.975 36.715 269.115 41.925 ;
        RECT 269.435 40.455 269.575 43.195 ;
        RECT 280.415 42.855 280.675 43.175 ;
        RECT 272.135 42.515 272.395 42.835 ;
        RECT 269.375 40.135 269.635 40.455 ;
        RECT 270.295 40.135 270.555 40.455 ;
        RECT 269.835 39.115 270.095 39.435 ;
        RECT 269.895 38.075 270.035 39.115 ;
        RECT 269.835 37.755 270.095 38.075 ;
        RECT 270.355 37.055 270.495 40.135 ;
        RECT 272.195 40.115 272.335 42.515 ;
        RECT 280.475 42.495 280.615 42.855 ;
        RECT 289.215 42.835 289.355 44.215 ;
        RECT 289.155 42.515 289.415 42.835 ;
        RECT 273.975 42.175 274.235 42.495 ;
        RECT 277.655 42.175 277.915 42.495 ;
        RECT 280.415 42.175 280.675 42.495 ;
        RECT 281.335 42.175 281.595 42.495 ;
        RECT 284.555 42.175 284.815 42.495 ;
        RECT 274.035 40.115 274.175 42.175 ;
        RECT 272.135 39.795 272.395 40.115 ;
        RECT 273.975 39.795 274.235 40.115 ;
        RECT 272.135 38.775 272.395 39.095 ;
        RECT 272.195 37.395 272.335 38.775 ;
        RECT 272.135 37.075 272.395 37.395 ;
        RECT 277.715 37.055 277.855 42.175 ;
        RECT 279.495 41.495 279.755 41.815 ;
        RECT 279.555 40.455 279.695 41.495 ;
        RECT 279.495 40.135 279.755 40.455 ;
        RECT 281.395 39.775 281.535 42.175 ;
        RECT 283.635 40.475 283.895 40.795 ;
        RECT 278.565 39.260 278.845 39.630 ;
        RECT 281.335 39.455 281.595 39.775 ;
        RECT 278.635 38.075 278.775 39.260 ;
        RECT 281.395 38.075 281.535 39.455 ;
        RECT 283.695 39.435 283.835 40.475 ;
        RECT 283.635 39.115 283.895 39.435 ;
        RECT 278.575 37.755 278.835 38.075 ;
        RECT 281.335 37.755 281.595 38.075 ;
        RECT 284.615 37.735 284.755 42.175 ;
        RECT 289.675 40.795 289.815 47.955 ;
        RECT 290.595 47.595 290.735 53.735 ;
        RECT 299.335 51.335 299.475 54.075 ;
        RECT 300.255 53.035 300.395 59.775 ;
        RECT 302.095 58.475 302.235 60.535 ;
        RECT 302.035 58.155 302.295 58.475 ;
        RECT 300.945 57.280 302.485 57.650 ;
        RECT 303.475 53.375 303.615 67.335 ;
        RECT 303.935 61.195 304.075 69.715 ;
        RECT 304.855 69.695 304.995 75.835 ;
        RECT 305.315 73.395 305.455 99.295 ;
        RECT 305.775 80.235 305.915 99.635 ;
        RECT 306.235 96.635 306.375 101.335 ;
        RECT 306.695 100.635 306.835 109.225 ;
        RECT 308.015 107.795 308.275 108.115 ;
        RECT 307.095 106.775 307.355 107.095 ;
        RECT 307.155 104.715 307.295 106.775 ;
        RECT 308.075 105.395 308.215 107.795 ;
        RECT 308.015 105.075 308.275 105.395 ;
        RECT 307.095 104.395 307.355 104.715 ;
        RECT 306.635 100.315 306.895 100.635 ;
        RECT 308.075 97.915 308.215 105.075 ;
        RECT 308.995 102.075 309.135 109.225 ;
        RECT 309.855 105.415 310.115 105.735 ;
        RECT 308.535 101.935 309.135 102.075 ;
        RECT 308.015 97.595 308.275 97.915 ;
        RECT 307.555 96.915 307.815 97.235 ;
        RECT 306.625 96.635 306.905 96.750 ;
        RECT 306.235 96.495 306.905 96.635 ;
        RECT 306.625 96.380 306.905 96.495 ;
        RECT 306.635 96.235 306.895 96.380 ;
        RECT 307.095 94.195 307.355 94.515 ;
        RECT 306.175 91.135 306.435 91.455 ;
        RECT 306.235 86.015 306.375 91.135 ;
        RECT 306.175 85.695 306.435 86.015 ;
        RECT 306.635 83.655 306.895 83.975 ;
        RECT 306.175 82.975 306.435 83.295 ;
        RECT 305.715 79.915 305.975 80.235 ;
        RECT 306.235 77.175 306.375 82.975 ;
        RECT 306.175 76.855 306.435 77.175 ;
        RECT 306.695 73.435 306.835 83.655 ;
        RECT 305.315 73.255 306.375 73.395 ;
        RECT 305.255 70.055 305.515 70.375 ;
        RECT 304.795 69.375 305.055 69.695 ;
        RECT 305.315 62.555 305.455 70.055 ;
        RECT 305.255 62.235 305.515 62.555 ;
        RECT 306.235 61.875 306.375 73.255 ;
        RECT 306.635 73.115 306.895 73.435 ;
        RECT 306.635 72.435 306.895 72.755 ;
        RECT 304.795 61.555 305.055 61.875 ;
        RECT 306.175 61.555 306.435 61.875 ;
        RECT 303.875 60.875 304.135 61.195 ;
        RECT 304.855 59.835 304.995 61.555 ;
        RECT 304.795 59.515 305.055 59.835 ;
        RECT 303.415 53.055 303.675 53.375 ;
        RECT 305.715 53.055 305.975 53.375 ;
        RECT 300.195 52.715 300.455 53.035 ;
        RECT 300.945 51.840 302.485 52.210 ;
        RECT 299.275 51.015 299.535 51.335 ;
        RECT 297.645 49.120 299.185 49.490 ;
        RECT 303.475 47.595 303.615 53.055 ;
        RECT 305.775 52.550 305.915 53.055 ;
        RECT 305.705 52.180 305.985 52.550 ;
        RECT 305.715 50.335 305.975 50.655 ;
        RECT 290.535 47.275 290.795 47.595 ;
        RECT 297.435 47.275 297.695 47.595 ;
        RECT 303.415 47.275 303.675 47.595 ;
        RECT 297.495 45.895 297.635 47.275 ;
        RECT 298.815 46.935 299.075 47.255 ;
        RECT 298.875 45.895 299.015 46.935 ;
        RECT 300.945 46.400 302.485 46.770 ;
        RECT 297.435 45.575 297.695 45.895 ;
        RECT 298.815 45.575 299.075 45.895 ;
        RECT 297.645 43.680 299.185 44.050 ;
        RECT 300.945 40.960 302.485 41.330 ;
        RECT 303.475 40.795 303.615 47.275 ;
        RECT 305.775 45.215 305.915 50.335 ;
        RECT 306.695 49.715 306.835 72.435 ;
        RECT 307.155 67.995 307.295 94.195 ;
        RECT 307.615 91.795 307.755 96.915 ;
        RECT 308.535 95.195 308.675 101.935 ;
        RECT 308.925 101.140 309.205 101.510 ;
        RECT 308.995 95.195 309.135 101.140 ;
        RECT 308.475 94.875 308.735 95.195 ;
        RECT 308.935 94.875 309.195 95.195 ;
        RECT 307.555 91.475 307.815 91.795 ;
        RECT 307.615 86.355 307.755 91.475 ;
        RECT 307.555 86.035 307.815 86.355 ;
        RECT 309.395 85.695 309.655 86.015 ;
        RECT 307.555 85.015 307.815 85.335 ;
        RECT 309.455 85.190 309.595 85.695 ;
        RECT 307.095 67.675 307.355 67.995 ;
        RECT 307.095 52.375 307.355 52.695 ;
        RECT 307.155 50.655 307.295 52.375 ;
        RECT 307.095 50.335 307.355 50.655 ;
        RECT 306.695 49.575 307.295 49.715 ;
        RECT 305.715 44.895 305.975 45.215 ;
        RECT 289.615 40.475 289.875 40.795 ;
        RECT 303.415 40.475 303.675 40.795 ;
        RECT 286.395 40.135 286.655 40.455 ;
        RECT 286.455 39.095 286.595 40.135 ;
        RECT 289.675 39.685 289.815 40.475 ;
        RECT 302.955 40.195 303.215 40.455 ;
        RECT 303.475 40.195 303.615 40.475 ;
        RECT 302.955 40.135 303.615 40.195 ;
        RECT 303.015 40.055 303.615 40.135 ;
        RECT 290.075 39.685 290.335 39.775 ;
        RECT 289.675 39.545 290.335 39.685 ;
        RECT 290.075 39.455 290.335 39.545 ;
        RECT 286.395 38.775 286.655 39.095 ;
        RECT 297.645 38.240 299.185 38.610 ;
        RECT 284.555 37.415 284.815 37.735 ;
        RECT 270.295 36.735 270.555 37.055 ;
        RECT 277.655 36.735 277.915 37.055 ;
        RECT 281.795 36.735 282.055 37.055 ;
        RECT 268.915 36.395 269.175 36.715 ;
        RECT 281.855 35.355 281.995 36.735 ;
        RECT 300.945 35.520 302.485 35.890 ;
        RECT 281.795 35.035 282.055 35.355 ;
        RECT 303.475 35.015 303.615 40.055 ;
        RECT 305.775 39.095 305.915 44.895 ;
        RECT 306.175 42.175 306.435 42.495 ;
        RECT 305.715 38.775 305.975 39.095 ;
        RECT 304.795 36.735 305.055 37.055 ;
        RECT 304.855 36.230 304.995 36.735 ;
        RECT 304.785 35.860 305.065 36.230 ;
        RECT 305.775 35.015 305.915 38.775 ;
        RECT 306.235 38.075 306.375 42.175 ;
        RECT 307.155 41.815 307.295 49.575 ;
        RECT 307.095 41.495 307.355 41.815 ;
        RECT 307.155 40.115 307.295 41.495 ;
        RECT 307.095 39.795 307.355 40.115 ;
        RECT 306.635 38.775 306.895 39.095 ;
        RECT 306.175 37.755 306.435 38.075 ;
        RECT 306.695 37.395 306.835 38.775 ;
        RECT 306.635 37.075 306.895 37.395 ;
        RECT 307.155 36.795 307.295 39.795 ;
        RECT 307.615 39.775 307.755 85.015 ;
        RECT 309.385 84.820 309.665 85.190 ;
        RECT 309.385 68.500 309.665 68.870 ;
        RECT 309.455 67.315 309.595 68.500 ;
        RECT 309.395 66.995 309.655 67.315 ;
        RECT 308.475 66.315 308.735 66.635 ;
        RECT 308.535 56.095 308.675 66.315 ;
        RECT 309.915 63.575 310.055 105.415 ;
        RECT 309.855 63.255 310.115 63.575 ;
        RECT 308.475 55.775 308.735 56.095 ;
        RECT 308.935 55.095 309.195 55.415 ;
        RECT 308.995 53.715 309.135 55.095 ;
        RECT 308.935 53.395 309.195 53.715 ;
        RECT 307.555 39.455 307.815 39.775 ;
        RECT 306.695 36.655 307.295 36.795 ;
        RECT 306.695 36.375 306.835 36.655 ;
        RECT 306.635 36.055 306.895 36.375 ;
        RECT 307.095 36.055 307.355 36.375 ;
        RECT 303.415 34.695 303.675 35.015 ;
        RECT 305.715 34.695 305.975 35.015 ;
        RECT 268.455 34.355 268.715 34.675 ;
        RECT 307.155 34.335 307.295 36.055 ;
        RECT 316.555 35.745 318.485 36.545 ;
        RECT 267.535 34.015 267.795 34.335 ;
        RECT 307.095 34.015 307.355 34.335 ;
        RECT 297.645 32.800 299.185 33.170 ;
        RECT 264.775 31.975 265.035 32.295 ;
        RECT 260.635 31.295 260.895 31.615 ;
        RECT 237.635 30.955 237.895 31.275 ;
        RECT 241.775 30.955 242.035 31.275 ;
        RECT 254.655 30.955 254.915 31.275 ;
        RECT 235.795 30.615 236.055 30.935 ;
        RECT 235.855 29.915 235.995 30.615 ;
        RECT 260.945 30.080 262.485 30.450 ;
        RECT 300.945 30.080 302.485 30.450 ;
        RECT 235.795 29.595 236.055 29.915 ;
        RECT 189.335 28.915 189.595 29.235 ;
        RECT 205.895 28.915 206.155 29.235 ;
        RECT 234.875 28.915 235.135 29.235 ;
        RECT 304.325 28.380 304.605 28.750 ;
        RECT 217.645 27.360 219.185 27.730 ;
        RECT 257.645 27.360 259.185 27.730 ;
        RECT 297.645 27.360 299.185 27.730 ;
        RECT 187.955 26.875 188.215 27.195 ;
        RECT 79.810 25.165 127.975 26.265 ;
        RECT 180.135 26.195 180.395 26.515 ;
        RECT 183.355 26.195 183.615 26.515 ;
        RECT 10.170 23.510 74.550 25.010 ;
        RECT 79.810 23.665 127.975 24.765 ;
        RECT 180.945 24.640 182.485 25.010 ;
        RECT 220.945 24.640 222.485 25.010 ;
        RECT 260.945 24.640 262.485 25.010 ;
        RECT 300.945 24.640 302.485 25.010 ;
        RECT 10.170 21.510 74.550 23.010 ;
        RECT 79.810 22.165 127.975 23.265 ;
        RECT 177.645 21.920 179.185 22.290 ;
        RECT 217.645 21.920 219.185 22.290 ;
        RECT 257.645 21.920 259.185 22.290 ;
        RECT 297.645 21.920 299.185 22.290 ;
        RECT 79.810 20.665 127.975 21.765 ;
        RECT 10.170 18.105 74.550 20.485 ;
        RECT 79.810 19.165 127.975 20.265 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 304.395 19.910 304.535 28.380 ;
        RECT 180.945 19.200 182.485 19.570 ;
        RECT 220.945 19.200 222.485 19.570 ;
        RECT 260.945 19.200 262.485 19.570 ;
        RECT 300.945 19.200 302.485 19.570 ;
        RECT 304.325 19.540 304.605 19.910 ;
        RECT 10.170 15.580 74.550 17.080 ;
        RECT 177.645 16.480 179.185 16.850 ;
        RECT 217.645 16.480 219.185 16.850 ;
        RECT 257.645 16.480 259.185 16.850 ;
        RECT 297.645 16.480 299.185 16.850 ;
        RECT 10.170 13.580 74.550 15.080 ;
        RECT 180.945 13.760 182.485 14.130 ;
        RECT 220.945 13.760 222.485 14.130 ;
        RECT 260.945 13.760 262.485 14.130 ;
        RECT 300.945 13.760 302.485 14.130 ;
        RECT 10.170 11.580 74.550 13.080 ;
        RECT 10.170 9.555 74.550 10.555 ;
        RECT 80.745 9.665 82.345 10.465 ;
        RECT 7.065 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.965 5.690 130.565 8.890 ;
      LAYER met3 ;
        RECT 125.730 225.710 126.530 225.760 ;
        RECT 23.260 225.160 23.660 225.560 ;
        RECT 1.000 224.760 23.660 225.160 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.310 65.510 225.710 ;
        RECT 125.730 225.410 252.160 225.710 ;
        RECT 125.730 225.360 126.530 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 1.000 221.560 1.400 224.760 ;
        RECT 67.470 224.710 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 75.700 223.310 76.100 224.860 ;
        RECT 75.700 222.910 76.500 223.310 ;
        RECT 78.545 222.710 78.945 224.860 ;
        RECT 78.545 222.310 79.345 222.710 ;
        RECT 83.980 222.110 84.380 224.860 ;
        RECT 83.980 221.710 84.780 222.110 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 86.740 221.510 87.140 224.860 ;
        RECT 86.740 221.110 87.540 221.510 ;
        RECT 92.260 220.910 92.660 224.860 ;
        RECT 129.375 224.750 251.225 225.050 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 108.865 224.515 109.665 224.615 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.915 106.460 224.450 ;
        RECT 108.865 224.215 129.040 224.515 ;
        RECT 95.070 221.515 95.370 223.650 ;
        RECT 97.830 222.115 98.130 223.650 ;
        RECT 100.590 222.715 100.890 223.650 ;
        RECT 103.350 223.315 103.650 223.650 ;
        RECT 106.060 223.615 125.010 223.915 ;
        RECT 103.350 223.015 120.980 223.315 ;
        RECT 100.590 222.415 116.950 222.715 ;
        RECT 97.830 221.815 112.920 222.115 ;
        RECT 95.070 221.215 108.890 221.515 ;
        RECT 92.260 220.510 93.060 220.910 ;
        RECT 1.000 218.590 12.150 220.190 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.920 188.640 10.720 211.890 ;
        RECT 15.720 198.970 38.920 209.370 ;
        RECT 9.520 187.840 11.120 188.640 ;
        RECT 15.720 186.970 38.920 197.370 ;
        RECT 44.120 188.440 44.920 211.890 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.520 182.990 11.120 183.790 ;
        RECT 3.600 176.050 7.510 179.250 ;
        RECT 9.920 163.040 10.720 182.990 ;
        RECT 15.720 174.970 38.920 185.370 ;
        RECT 45.870 181.190 46.670 210.555 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 47.470 182.790 48.270 204.590 ;
        RECT 108.590 202.625 108.890 221.215 ;
        RECT 109.240 207.925 109.640 219.305 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 111.820 207.925 112.220 219.305 ;
        RECT 109.240 207.525 110.490 207.925 ;
        RECT 108.540 201.825 108.940 202.625 ;
        RECT 63.550 200.610 98.400 200.615 ;
        RECT 63.550 199.815 106.330 200.610 ;
        RECT 98.400 199.810 106.330 199.815 ;
        RECT 68.970 196.830 100.300 197.630 ;
        RECT 74.545 193.735 98.000 194.535 ;
        RECT 66.295 190.655 95.650 191.455 ;
        RECT 52.860 188.465 53.660 190.065 ;
        RECT 55.320 184.940 56.920 186.540 ;
        RECT 47.470 181.990 54.670 182.790 ;
        RECT 45.870 180.390 53.020 181.190 ;
        RECT 9.520 162.240 11.120 163.040 ;
        RECT 15.720 162.970 38.920 173.370 ;
        RECT 52.220 170.440 53.020 180.390 ;
        RECT 53.870 175.290 54.670 181.990 ;
        RECT 53.870 164.840 54.670 174.240 ;
        RECT 55.720 166.640 56.520 184.940 ;
        RECT 57.020 177.390 57.820 178.990 ;
        RECT 61.980 174.370 90.220 175.170 ;
        RECT 57.020 168.290 57.820 169.890 ;
        RECT 55.320 165.840 56.920 166.640 ;
        RECT 53.470 164.040 55.070 164.840 ;
        RECT 9.920 153.790 10.720 162.240 ;
        RECT 9.520 152.990 11.120 153.790 ;
        RECT 9.920 152.915 10.720 152.990 ;
        RECT 15.720 150.970 38.920 161.370 ;
        RECT 51.570 160.190 53.170 160.990 ;
        RECT 51.970 155.790 52.770 160.190 ;
        RECT 51.570 154.990 53.170 155.790 ;
        RECT 41.830 149.410 46.630 150.210 ;
        RECT 51.970 148.290 52.770 154.990 ;
        RECT 53.870 151.990 54.670 164.040 ;
        RECT 53.470 151.190 55.070 151.990 ;
        RECT 55.720 150.240 56.520 165.840 ;
        RECT 54.920 149.440 56.520 150.240 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 61.980 143.690 62.780 174.370 ;
        RECT 3.600 132.225 7.510 135.425 ;
        RECT 9.095 134.635 18.955 143.035 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 28.140 142.890 62.780 143.690 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 20.650 131.410 21.050 138.770 ;
        RECT 61.980 135.095 62.780 142.890 ;
        RECT 70.165 172.130 84.650 172.930 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 12.915 45.565 14.515 119.215 ;
        RECT 16.165 56.765 17.765 121.615 ;
        RECT 21.615 95.165 22.415 132.545 ;
        RECT 27.065 95.165 27.865 130.795 ;
        RECT 70.165 128.125 70.965 172.130 ;
        RECT 74.940 154.795 86.100 155.595 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 145.235 75.740 154.795 ;
        RECT 94.850 150.520 95.650 190.655 ;
        RECT 80.010 149.520 95.650 150.520 ;
        RECT 74.940 144.435 86.100 145.235 ;
        RECT 63.315 103.770 64.915 123.715 ;
        RECT 65.865 110.280 67.465 127.485 ;
        RECT 75.510 123.715 77.110 135.155 ;
        RECT 80.125 133.320 80.925 144.435 ;
        RECT 94.850 131.745 95.650 149.520 ;
        RECT 97.200 137.420 98.000 193.735 ;
        RECT 99.500 129.995 100.300 196.830 ;
        RECT 102.950 168.255 103.750 186.540 ;
        RECT 105.530 170.890 106.330 199.810 ;
        RECT 109.240 198.885 109.640 205.545 ;
        RECT 110.090 197.895 110.490 207.525 ;
        RECT 109.240 197.495 110.490 197.895 ;
        RECT 110.970 207.525 112.220 207.925 ;
        RECT 110.970 197.895 111.370 207.525 ;
        RECT 111.820 198.885 112.220 206.755 ;
        RECT 112.620 202.625 112.920 221.815 ;
        RECT 113.270 207.925 113.670 219.305 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 115.850 207.925 116.250 219.305 ;
        RECT 113.270 207.525 114.520 207.925 ;
        RECT 112.570 201.825 112.970 202.625 ;
        RECT 113.270 198.885 113.670 205.545 ;
        RECT 114.120 197.895 114.520 207.525 ;
        RECT 110.970 197.495 112.220 197.895 ;
        RECT 109.240 183.970 109.640 197.495 ;
        RECT 111.820 191.285 112.220 197.495 ;
        RECT 113.270 197.495 114.520 197.895 ;
        RECT 115.000 207.525 116.250 207.925 ;
        RECT 115.000 197.895 115.400 207.525 ;
        RECT 115.850 198.885 116.250 206.755 ;
        RECT 116.650 202.625 116.950 222.415 ;
        RECT 117.300 207.925 117.700 219.305 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 119.880 207.925 120.280 219.305 ;
        RECT 117.300 207.525 118.550 207.925 ;
        RECT 116.600 201.825 117.000 202.625 ;
        RECT 117.300 198.885 117.700 205.545 ;
        RECT 118.150 197.895 118.550 207.525 ;
        RECT 115.000 197.495 116.250 197.895 ;
        RECT 110.530 187.540 110.930 189.140 ;
        RECT 113.270 183.990 113.670 197.495 ;
        RECT 115.850 191.285 116.250 197.495 ;
        RECT 117.300 197.495 118.550 197.895 ;
        RECT 119.030 207.525 120.280 207.925 ;
        RECT 119.030 197.895 119.430 207.525 ;
        RECT 119.880 198.885 120.280 206.755 ;
        RECT 120.680 202.625 120.980 223.015 ;
        RECT 121.330 207.925 121.730 219.305 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 123.910 207.925 124.310 219.305 ;
        RECT 121.330 207.525 122.580 207.925 ;
        RECT 120.630 201.825 121.030 202.625 ;
        RECT 121.330 198.885 121.730 205.545 ;
        RECT 122.180 197.895 122.580 207.525 ;
        RECT 119.030 197.495 120.280 197.895 ;
        RECT 114.560 187.540 114.960 189.140 ;
        RECT 111.685 183.590 113.670 183.990 ;
        RECT 105.530 168.255 106.730 170.890 ;
        RECT 107.380 168.490 107.780 170.890 ;
        RECT 103.350 152.765 103.750 160.495 ;
        RECT 103.350 143.435 103.750 145.835 ;
        RECT 104.640 140.165 105.040 167.190 ;
        RECT 105.385 157.365 105.785 158.165 ;
        RECT 106.330 145.835 106.730 168.255 ;
        RECT 107.380 152.765 107.780 160.495 ;
        RECT 108.670 147.135 109.070 178.990 ;
        RECT 109.960 168.490 110.760 170.890 ;
        RECT 109.415 156.165 109.815 156.965 ;
        RECT 110.360 145.835 110.760 168.490 ;
        RECT 111.685 157.765 112.085 183.590 ;
        RECT 117.300 182.580 117.700 197.495 ;
        RECT 119.880 191.285 120.280 197.495 ;
        RECT 121.330 197.495 122.580 197.895 ;
        RECT 123.060 207.525 124.310 207.925 ;
        RECT 123.060 197.895 123.460 207.525 ;
        RECT 123.910 198.885 124.310 206.755 ;
        RECT 124.710 202.625 125.010 223.615 ;
        RECT 125.360 207.925 125.760 219.305 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 127.940 207.925 128.340 219.305 ;
        RECT 125.360 207.525 126.610 207.925 ;
        RECT 124.660 201.825 125.060 202.625 ;
        RECT 125.360 198.885 125.760 205.545 ;
        RECT 126.210 197.895 126.610 207.525 ;
        RECT 123.060 197.495 124.310 197.895 ;
        RECT 118.590 187.540 118.990 189.140 ;
        RECT 113.085 182.180 117.700 182.580 ;
        RECT 113.085 156.165 113.485 182.180 ;
        RECT 121.330 181.545 121.730 197.495 ;
        RECT 123.910 191.285 124.310 197.495 ;
        RECT 125.360 197.495 126.610 197.895 ;
        RECT 127.090 207.525 128.340 207.925 ;
        RECT 127.090 197.895 127.490 207.525 ;
        RECT 127.940 198.885 128.340 206.755 ;
        RECT 128.740 202.625 129.040 224.215 ;
        RECT 132.720 220.715 133.120 221.515 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 129.390 207.925 129.790 219.305 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 131.970 207.925 132.370 219.305 ;
        RECT 129.390 207.525 130.640 207.925 ;
        RECT 128.690 201.825 129.090 202.625 ;
        RECT 129.390 198.885 129.790 205.545 ;
        RECT 130.240 197.895 130.640 207.525 ;
        RECT 127.090 197.495 128.340 197.895 ;
        RECT 122.620 187.540 123.020 189.140 ;
        RECT 116.415 181.145 121.730 181.545 ;
        RECT 116.415 176.215 116.815 181.145 ;
        RECT 125.360 180.565 125.760 197.495 ;
        RECT 127.940 191.285 128.340 197.495 ;
        RECT 129.390 197.495 130.640 197.895 ;
        RECT 131.120 207.525 132.370 207.925 ;
        RECT 131.120 197.895 131.520 207.525 ;
        RECT 131.970 198.885 132.370 206.755 ;
        RECT 132.770 202.625 133.070 220.715 ;
        RECT 133.420 207.925 133.820 219.305 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 136.000 207.925 136.400 219.305 ;
        RECT 133.420 207.525 134.670 207.925 ;
        RECT 132.720 201.825 133.120 202.625 ;
        RECT 133.420 198.885 133.820 205.545 ;
        RECT 134.270 197.895 134.670 207.525 ;
        RECT 131.120 197.495 132.370 197.895 ;
        RECT 126.650 187.540 127.050 189.140 ;
        RECT 121.035 180.165 125.760 180.565 ;
        RECT 121.035 176.215 121.435 180.165 ;
        RECT 129.390 179.490 129.790 197.495 ;
        RECT 131.970 191.285 132.370 197.495 ;
        RECT 133.420 197.495 134.670 197.895 ;
        RECT 135.150 207.525 136.400 207.925 ;
        RECT 135.150 197.895 135.550 207.525 ;
        RECT 136.000 198.885 136.400 206.755 ;
        RECT 136.800 202.625 137.100 220.715 ;
        RECT 137.450 207.925 137.850 219.305 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 140.030 207.925 140.430 219.305 ;
        RECT 137.450 207.525 138.700 207.925 ;
        RECT 136.750 201.825 137.150 202.625 ;
        RECT 137.450 198.885 137.850 205.545 ;
        RECT 138.300 197.895 138.700 207.525 ;
        RECT 135.150 197.495 136.400 197.895 ;
        RECT 130.680 187.540 131.080 189.140 ;
        RECT 125.660 179.090 129.790 179.490 ;
        RECT 125.660 176.215 126.060 179.090 ;
        RECT 133.420 178.920 133.820 197.495 ;
        RECT 136.000 191.285 136.400 197.495 ;
        RECT 137.450 197.495 138.700 197.895 ;
        RECT 139.180 207.525 140.430 207.925 ;
        RECT 139.180 197.895 139.580 207.525 ;
        RECT 140.030 198.885 140.430 206.755 ;
        RECT 140.830 202.625 141.130 220.715 ;
        RECT 141.480 207.925 141.880 219.305 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 144.060 207.925 144.460 219.305 ;
        RECT 141.480 207.525 142.730 207.925 ;
        RECT 140.780 201.825 141.180 202.625 ;
        RECT 141.480 198.885 141.880 205.545 ;
        RECT 142.330 197.895 142.730 207.525 ;
        RECT 139.180 197.495 140.430 197.895 ;
        RECT 134.710 187.540 135.110 189.140 ;
        RECT 137.450 178.920 137.850 197.495 ;
        RECT 140.030 191.285 140.430 197.495 ;
        RECT 141.480 197.495 142.730 197.895 ;
        RECT 143.210 207.525 144.460 207.925 ;
        RECT 143.210 197.895 143.610 207.525 ;
        RECT 144.060 198.885 144.460 206.755 ;
        RECT 144.860 202.625 145.160 220.715 ;
        RECT 145.510 207.925 145.910 219.305 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 148.090 207.925 148.490 219.305 ;
        RECT 145.510 207.525 146.760 207.925 ;
        RECT 144.810 201.825 145.210 202.625 ;
        RECT 145.510 198.885 145.910 205.545 ;
        RECT 146.360 197.895 146.760 207.525 ;
        RECT 143.210 197.495 144.460 197.895 ;
        RECT 138.740 187.540 139.140 189.140 ;
        RECT 141.480 178.920 141.880 197.495 ;
        RECT 144.060 191.285 144.460 197.495 ;
        RECT 145.510 197.495 146.760 197.895 ;
        RECT 147.240 207.525 148.490 207.925 ;
        RECT 147.240 197.895 147.640 207.525 ;
        RECT 148.090 198.885 148.490 206.755 ;
        RECT 148.890 202.625 149.190 220.715 ;
        RECT 162.100 220.260 162.500 220.910 ;
        RECT 163.100 220.860 163.500 221.510 ;
        RECT 164.100 221.460 164.500 222.110 ;
        RECT 164.100 221.160 250.220 221.460 ;
        RECT 163.100 220.560 249.370 220.860 ;
        RECT 162.100 219.960 248.285 220.260 ;
        RECT 149.540 207.925 149.940 219.305 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 152.120 207.925 152.520 219.305 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 180.915 212.210 222.515 213.810 ;
        RECT 177.615 209.640 219.215 211.240 ;
        RECT 149.540 207.525 150.790 207.925 ;
        RECT 148.840 201.825 149.240 202.625 ;
        RECT 149.540 198.885 149.940 205.545 ;
        RECT 150.390 197.895 150.790 207.525 ;
        RECT 147.240 197.495 148.490 197.895 ;
        RECT 142.770 187.540 143.170 189.140 ;
        RECT 145.510 178.920 145.910 197.495 ;
        RECT 148.090 191.285 148.490 197.495 ;
        RECT 149.540 197.495 150.790 197.895 ;
        RECT 151.270 207.525 152.520 207.925 ;
        RECT 151.270 197.895 151.670 207.525 ;
        RECT 152.120 198.885 152.520 206.755 ;
        RECT 177.625 201.325 179.205 201.655 ;
        RECT 217.625 201.325 219.205 201.655 ;
        RECT 180.925 198.605 182.505 198.935 ;
        RECT 220.925 198.605 222.505 198.935 ;
        RECT 159.335 197.900 161.335 198.050 ;
        RECT 164.000 197.900 164.330 197.915 ;
        RECT 151.270 197.495 152.520 197.895 ;
        RECT 146.800 187.540 147.200 189.140 ;
        RECT 149.540 178.920 149.940 197.495 ;
        RECT 152.120 191.285 152.520 197.495 ;
        RECT 157.560 197.600 164.330 197.900 ;
        RECT 150.830 187.540 151.230 189.140 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 130.275 178.520 133.820 178.920 ;
        RECT 134.895 178.520 137.850 178.920 ;
        RECT 139.510 178.520 141.880 178.920 ;
        RECT 144.135 178.520 145.910 178.920 ;
        RECT 148.755 178.520 149.940 178.920 ;
        RECT 130.275 176.215 130.675 178.520 ;
        RECT 134.895 176.215 135.295 178.520 ;
        RECT 139.510 176.215 139.910 178.520 ;
        RECT 144.135 176.215 144.535 178.520 ;
        RECT 148.755 176.215 149.155 178.520 ;
        RECT 116.215 175.815 117.015 176.215 ;
        RECT 120.835 175.815 121.635 176.215 ;
        RECT 125.455 175.815 126.255 176.215 ;
        RECT 130.075 175.815 130.875 176.215 ;
        RECT 134.695 175.815 135.495 176.215 ;
        RECT 139.315 175.815 140.115 176.215 ;
        RECT 143.935 175.815 144.735 176.215 ;
        RECT 148.555 175.815 149.355 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 115.815 173.070 117.415 173.870 ;
        RECT 120.435 173.070 122.035 173.870 ;
        RECT 125.055 173.070 126.655 173.870 ;
        RECT 129.675 173.070 131.275 173.870 ;
        RECT 134.295 173.070 135.895 173.870 ;
        RECT 138.915 173.070 140.515 173.870 ;
        RECT 143.535 173.070 145.135 173.870 ;
        RECT 148.155 173.070 149.755 173.870 ;
        RECT 105.930 143.435 106.730 145.835 ;
        RECT 104.640 139.365 105.440 140.165 ;
        RECT 107.380 136.325 107.780 145.835 ;
        RECT 109.960 143.435 110.760 145.835 ;
        RECT 116.310 144.730 116.910 173.070 ;
        RECT 120.930 147.530 121.530 173.070 ;
        RECT 125.550 148.690 126.150 173.070 ;
        RECT 130.175 149.890 130.775 173.070 ;
        RECT 134.795 160.260 135.395 173.070 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 133.275 152.100 134.875 152.200 ;
        RECT 136.875 152.100 137.475 161.650 ;
        RECT 133.275 151.500 137.475 152.100 ;
        RECT 133.275 151.400 134.875 151.500 ;
        RECT 133.275 150.930 134.875 151.030 ;
        RECT 139.410 150.930 140.010 173.070 ;
        RECT 144.035 162.450 144.635 173.070 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 148.655 161.210 149.255 173.070 ;
        RECT 133.275 150.330 140.010 150.930 ;
        RECT 141.715 160.610 149.255 161.210 ;
        RECT 133.275 150.230 134.875 150.330 ;
        RECT 130.175 149.290 136.695 149.890 ;
        RECT 125.550 148.090 133.635 148.690 ;
        RECT 130.615 147.530 132.215 147.630 ;
        RECT 120.930 146.930 132.215 147.530 ;
        RECT 130.615 146.830 132.215 146.930 ;
        RECT 122.645 144.730 124.245 144.830 ;
        RECT 116.310 144.130 124.245 144.730 ;
        RECT 122.645 144.030 124.245 144.130 ;
        RECT 133.035 144.520 133.635 148.090 ;
        RECT 136.095 148.010 136.695 149.290 ;
        RECT 138.525 148.010 140.125 148.110 ;
        RECT 136.095 147.410 140.125 148.010 ;
        RECT 138.525 147.310 140.125 147.410 ;
        RECT 138.525 144.520 140.125 144.620 ;
        RECT 133.035 143.920 140.125 144.520 ;
        RECT 141.715 144.040 142.315 160.610 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 138.525 143.820 140.125 143.920 ;
        RECT 109.960 138.220 110.360 143.435 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 142.690 142.815 142.790 ;
        RECT 145.625 142.690 146.225 159.460 ;
        RECT 141.215 142.090 146.225 142.690 ;
        RECT 141.215 141.990 142.815 142.090 ;
        RECT 109.560 137.420 110.760 138.220 ;
        RECT 107.380 135.525 108.180 136.325 ;
        RECT 72.765 103.865 74.365 122.215 ;
        RECT 75.510 114.215 77.115 123.715 ;
        RECT 75.515 100.215 77.115 114.215 ;
        RECT 21.215 51.675 22.815 95.165 ;
        RECT 26.665 61.465 28.265 95.165 ;
        RECT 97.165 93.265 98.765 119.215 ;
        RECT 100.515 117.715 101.315 128.925 ;
        RECT 100.115 96.415 101.715 117.715 ;
        RECT 103.315 111.365 104.915 123.165 ;
        RECT 116.915 121.965 118.515 122.765 ;
        RECT 105.965 103.965 107.565 120.665 ;
        RECT 109.865 108.365 111.465 119.215 ;
        RECT 117.115 108.365 118.715 118.265 ;
        RECT 121.565 113.015 123.165 127.485 ;
        RECT 116.965 104.015 118.565 104.815 ;
        RECT 42.740 71.190 53.140 83.050 ;
        RECT 55.740 71.190 66.140 83.050 ;
        RECT 68.740 71.190 79.140 83.050 ;
        RECT 81.740 71.190 92.140 83.050 ;
        RECT 94.740 71.190 105.140 83.050 ;
        RECT 42.740 57.830 53.140 69.690 ;
        RECT 55.740 57.830 66.140 69.690 ;
        RECT 68.740 57.830 79.140 69.690 ;
        RECT 81.740 57.830 92.140 69.690 ;
        RECT 94.740 57.830 105.140 69.690 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 3.600 36.430 8.665 39.630 ;
        RECT 3.600 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 34.940 ;
        RECT 65.765 15.915 67.365 44.215 ;
        RECT 68.865 11.965 70.465 41.615 ;
        RECT 72.095 9.665 73.695 38.865 ;
        RECT 80.745 9.665 82.345 37.635 ;
        RECT 84.015 22.315 85.615 41.615 ;
        RECT 87.165 26.815 88.765 44.215 ;
        RECT 90.715 19.315 92.315 47.165 ;
        RECT 116.115 42.615 117.715 90.815 ;
        RECT 119.215 40.015 120.815 84.315 ;
        RECT 123.215 23.815 124.815 94.865 ;
        RECT 126.165 25.365 127.765 98.015 ;
        RECT 128.965 5.690 130.565 8.890 ;
        RECT 2.705 1.285 98.380 2.085 ;
        RECT 131.665 1.800 132.465 136.325 ;
        RECT 133.265 111.795 134.065 130.795 ;
        RECT 134.865 110.315 135.665 132.545 ;
        RECT 136.465 114.770 137.265 134.120 ;
        RECT 137.945 133.410 138.745 133.810 ;
        RECT 137.945 131.410 138.345 133.410 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.970 125.690 142.100 127.290 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 133.525 109.515 138.400 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 136.495 29.375 138.195 94.305 ;
        RECT 139.355 30.545 141.055 114.150 ;
        RECT 141.900 110.315 142.700 117.170 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 141.495 20.015 143.195 110.315 ;
        RECT 143.640 32.885 145.340 114.150 ;
        RECT 146.950 110.315 147.750 138.220 ;
        RECT 149.945 116.370 150.745 170.845 ;
        RECT 146.490 104.255 148.190 110.315 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 151.560 1.800 152.360 140.165 ;
        RECT 153.945 129.145 154.345 184.370 ;
        RECT 157.560 28.035 157.860 197.600 ;
        RECT 159.335 197.450 161.335 197.600 ;
        RECT 164.000 197.585 164.330 197.600 ;
        RECT 177.625 195.885 179.205 196.215 ;
        RECT 217.625 195.885 219.205 196.215 ;
        RECT 180.925 193.165 182.505 193.495 ;
        RECT 220.925 193.165 222.505 193.495 ;
        RECT 177.625 190.445 179.205 190.775 ;
        RECT 217.625 190.445 219.205 190.775 ;
        RECT 177.340 189.740 177.670 189.755 ;
        RECT 185.160 189.740 185.490 189.755 ;
        RECT 186.540 189.750 186.870 189.755 ;
        RECT 186.285 189.740 186.870 189.750 ;
        RECT 177.340 189.440 185.490 189.740 ;
        RECT 186.085 189.440 186.870 189.740 ;
        RECT 177.340 189.425 177.670 189.440 ;
        RECT 185.160 189.425 185.490 189.440 ;
        RECT 186.285 189.430 186.870 189.440 ;
        RECT 186.540 189.425 186.870 189.430 ;
        RECT 202.640 189.740 202.970 189.755 ;
        RECT 207.445 189.740 207.825 189.750 ;
        RECT 202.640 189.440 207.825 189.740 ;
        RECT 202.640 189.425 202.970 189.440 ;
        RECT 207.445 189.430 207.825 189.440 ;
        RECT 174.580 189.060 174.910 189.075 ;
        RECT 188.840 189.060 189.170 189.075 ;
        RECT 174.580 188.760 189.170 189.060 ;
        RECT 174.580 188.745 174.910 188.760 ;
        RECT 188.840 188.745 189.170 188.760 ;
        RECT 159.335 188.380 161.335 188.530 ;
        RECT 163.540 188.380 163.870 188.395 ;
        RECT 169.980 188.380 170.310 188.395 ;
        RECT 176.880 188.380 177.210 188.395 ;
        RECT 179.180 188.380 179.510 188.395 ;
        RECT 158.335 188.080 164.390 188.380 ;
        RECT 169.980 188.080 179.510 188.380 ;
        RECT 158.335 60.675 158.635 188.080 ;
        RECT 159.335 187.930 161.335 188.080 ;
        RECT 163.540 188.065 163.870 188.080 ;
        RECT 169.980 188.065 170.310 188.080 ;
        RECT 176.880 188.065 177.210 188.080 ;
        RECT 179.180 188.065 179.510 188.080 ;
        RECT 180.925 187.725 182.505 188.055 ;
        RECT 220.925 187.725 222.505 188.055 ;
        RECT 169.520 187.700 169.850 187.715 ;
        RECT 170.900 187.700 171.230 187.715 ;
        RECT 169.520 187.400 171.230 187.700 ;
        RECT 169.520 187.385 169.850 187.400 ;
        RECT 170.900 187.385 171.230 187.400 ;
        RECT 186.080 187.700 186.410 187.715 ;
        RECT 189.300 187.700 189.630 187.715 ;
        RECT 186.080 187.400 189.630 187.700 ;
        RECT 186.080 187.385 186.410 187.400 ;
        RECT 189.300 187.385 189.630 187.400 ;
        RECT 181.020 187.020 181.350 187.035 ;
        RECT 192.520 187.020 192.850 187.035 ;
        RECT 181.020 186.720 192.850 187.020 ;
        RECT 181.020 186.705 181.350 186.720 ;
        RECT 192.520 186.705 192.850 186.720 ;
        RECT 208.160 187.020 208.490 187.035 ;
        RECT 224.720 187.020 225.050 187.035 ;
        RECT 208.160 186.720 225.050 187.020 ;
        RECT 208.160 186.705 208.490 186.720 ;
        RECT 224.720 186.705 225.050 186.720 ;
        RECT 176.880 186.340 177.210 186.355 ;
        RECT 214.600 186.340 214.930 186.355 ;
        RECT 176.880 186.040 214.930 186.340 ;
        RECT 176.880 186.025 177.210 186.040 ;
        RECT 214.600 186.025 214.930 186.040 ;
        RECT 209.285 185.660 209.665 185.670 ;
        RECT 210.460 185.660 210.790 185.675 ;
        RECT 209.285 185.360 210.790 185.660 ;
        RECT 209.285 185.350 209.665 185.360 ;
        RECT 210.460 185.345 210.790 185.360 ;
        RECT 177.625 185.005 179.205 185.335 ;
        RECT 217.625 185.005 219.205 185.335 ;
        RECT 207.700 184.980 208.030 184.995 ;
        RECT 208.620 184.980 208.950 184.995 ;
        RECT 207.700 184.680 208.950 184.980 ;
        RECT 207.700 184.665 208.030 184.680 ;
        RECT 208.620 184.665 208.950 184.680 ;
        RECT 171.360 184.300 171.690 184.315 ;
        RECT 175.500 184.300 175.830 184.315 ;
        RECT 171.360 184.000 175.830 184.300 ;
        RECT 171.360 183.985 171.690 184.000 ;
        RECT 175.500 183.985 175.830 184.000 ;
        RECT 188.840 184.300 189.170 184.315 ;
        RECT 192.520 184.300 192.850 184.315 ;
        RECT 195.280 184.300 195.610 184.315 ;
        RECT 231.160 184.300 231.490 184.315 ;
        RECT 188.840 184.000 195.610 184.300 ;
        RECT 188.840 183.985 189.170 184.000 ;
        RECT 192.520 183.985 192.850 184.000 ;
        RECT 195.280 183.985 195.610 184.000 ;
        RECT 206.565 184.000 231.490 184.300 ;
        RECT 181.480 183.620 181.810 183.635 ;
        RECT 195.280 183.620 195.610 183.635 ;
        RECT 181.480 183.320 195.610 183.620 ;
        RECT 181.480 183.305 181.810 183.320 ;
        RECT 195.280 183.305 195.610 183.320 ;
        RECT 172.740 182.940 173.070 182.955 ;
        RECT 177.340 182.940 177.670 182.955 ;
        RECT 172.740 182.640 177.670 182.940 ;
        RECT 172.740 182.625 173.070 182.640 ;
        RECT 177.340 182.625 177.670 182.640 ;
        RECT 192.520 182.940 192.850 182.955 ;
        RECT 206.565 182.940 206.865 184.000 ;
        RECT 231.160 183.985 231.490 184.000 ;
        RECT 208.160 183.620 208.490 183.635 ;
        RECT 209.080 183.620 209.410 183.635 ;
        RECT 208.160 183.320 209.410 183.620 ;
        RECT 208.160 183.305 208.490 183.320 ;
        RECT 209.080 183.305 209.410 183.320 ;
        RECT 210.460 183.620 210.790 183.635 ;
        RECT 228.860 183.620 229.190 183.635 ;
        RECT 210.460 183.320 229.190 183.620 ;
        RECT 210.460 183.305 210.790 183.320 ;
        RECT 228.860 183.305 229.190 183.320 ;
        RECT 192.520 182.640 206.865 182.940 ;
        RECT 207.240 182.940 207.570 182.955 ;
        RECT 220.120 182.940 220.450 182.955 ;
        RECT 207.240 182.640 220.450 182.940 ;
        RECT 192.520 182.625 192.850 182.640 ;
        RECT 207.240 182.625 207.570 182.640 ;
        RECT 220.120 182.625 220.450 182.640 ;
        RECT 180.925 182.285 182.505 182.615 ;
        RECT 220.925 182.285 222.505 182.615 ;
        RECT 169.060 182.260 169.390 182.275 ;
        RECT 169.980 182.260 170.310 182.275 ;
        RECT 169.060 181.960 170.310 182.260 ;
        RECT 169.060 181.945 169.390 181.960 ;
        RECT 169.980 181.945 170.310 181.960 ;
        RECT 170.900 182.260 171.230 182.275 ;
        RECT 175.500 182.260 175.830 182.275 ;
        RECT 213.680 182.260 214.010 182.275 ;
        RECT 170.900 181.960 175.830 182.260 ;
        RECT 170.900 181.945 171.230 181.960 ;
        RECT 175.500 181.945 175.830 181.960 ;
        RECT 211.165 181.960 214.010 182.260 ;
        RECT 164.920 181.580 165.250 181.595 ;
        RECT 172.740 181.580 173.070 181.595 ;
        RECT 164.920 181.280 173.070 181.580 ;
        RECT 164.920 181.265 165.250 181.280 ;
        RECT 172.740 181.265 173.070 181.280 ;
        RECT 181.940 181.580 182.270 181.595 ;
        RECT 191.600 181.580 191.930 181.595 ;
        RECT 181.940 181.280 191.930 181.580 ;
        RECT 181.940 181.265 182.270 181.280 ;
        RECT 191.600 181.265 191.930 181.280 ;
        RECT 171.820 180.900 172.150 180.915 ;
        RECT 211.165 180.900 211.465 181.960 ;
        RECT 213.680 181.945 214.010 181.960 ;
        RECT 211.840 181.580 212.170 181.595 ;
        RECT 232.540 181.580 232.870 181.595 ;
        RECT 211.840 181.280 232.870 181.580 ;
        RECT 211.840 181.265 212.170 181.280 ;
        RECT 232.540 181.265 232.870 181.280 ;
        RECT 171.820 180.600 211.465 180.900 ;
        RECT 215.980 180.900 216.310 180.915 ;
        RECT 217.360 180.900 217.690 180.915 ;
        RECT 215.980 180.600 217.690 180.900 ;
        RECT 171.820 180.585 172.150 180.600 ;
        RECT 215.980 180.585 216.310 180.600 ;
        RECT 217.360 180.585 217.690 180.600 ;
        RECT 218.740 180.900 219.070 180.915 ;
        RECT 231.160 180.900 231.490 180.915 ;
        RECT 218.740 180.600 231.490 180.900 ;
        RECT 218.740 180.585 219.070 180.600 ;
        RECT 231.160 180.585 231.490 180.600 ;
        RECT 189.760 180.220 190.090 180.235 ;
        RECT 190.680 180.220 191.010 180.235 ;
        RECT 189.760 179.920 191.010 180.220 ;
        RECT 189.760 179.905 190.090 179.920 ;
        RECT 190.680 179.905 191.010 179.920 ;
        RECT 208.620 180.220 208.950 180.235 ;
        RECT 209.285 180.220 209.665 180.230 ;
        RECT 208.620 179.920 209.665 180.220 ;
        RECT 208.620 179.905 208.950 179.920 ;
        RECT 209.285 179.910 209.665 179.920 ;
        RECT 220.120 180.220 220.450 180.235 ;
        RECT 222.880 180.220 223.210 180.235 ;
        RECT 220.120 179.920 223.210 180.220 ;
        RECT 220.120 179.905 220.450 179.920 ;
        RECT 222.880 179.905 223.210 179.920 ;
        RECT 227.020 180.220 227.350 180.235 ;
        RECT 230.700 180.220 231.030 180.235 ;
        RECT 227.020 179.920 231.030 180.220 ;
        RECT 227.020 179.905 227.350 179.920 ;
        RECT 230.700 179.905 231.030 179.920 ;
        RECT 177.625 179.565 179.205 179.895 ;
        RECT 217.625 179.565 219.205 179.895 ;
        RECT 210.460 179.540 210.790 179.555 ;
        RECT 214.600 179.540 214.930 179.555 ;
        RECT 223.340 179.550 223.670 179.555 ;
        RECT 223.085 179.540 223.670 179.550 ;
        RECT 210.460 179.240 214.930 179.540 ;
        RECT 222.885 179.240 223.670 179.540 ;
        RECT 210.460 179.225 210.790 179.240 ;
        RECT 214.600 179.225 214.930 179.240 ;
        RECT 223.085 179.230 223.670 179.240 ;
        RECT 223.340 179.225 223.670 179.230 ;
        RECT 224.260 179.540 224.590 179.555 ;
        RECT 233.460 179.540 233.790 179.555 ;
        RECT 224.260 179.240 233.790 179.540 ;
        RECT 224.260 179.225 224.590 179.240 ;
        RECT 233.460 179.225 233.790 179.240 ;
        RECT 159.335 178.860 161.335 179.010 ;
        RECT 163.540 178.860 163.870 178.875 ;
        RECT 159.185 178.560 163.870 178.860 ;
        RECT 159.185 178.410 161.335 178.560 ;
        RECT 163.540 178.545 163.870 178.560 ;
        RECT 168.600 178.860 168.930 178.875 ;
        RECT 175.960 178.860 176.290 178.875 ;
        RECT 168.600 178.560 176.290 178.860 ;
        RECT 168.600 178.545 168.930 178.560 ;
        RECT 175.960 178.545 176.290 178.560 ;
        RECT 186.540 178.860 186.870 178.875 ;
        RECT 191.600 178.860 191.930 178.875 ;
        RECT 186.540 178.560 191.930 178.860 ;
        RECT 186.540 178.545 186.870 178.560 ;
        RECT 191.600 178.545 191.930 178.560 ;
        RECT 209.080 178.860 209.410 178.875 ;
        RECT 229.780 178.860 230.110 178.875 ;
        RECT 209.080 178.560 230.110 178.860 ;
        RECT 209.080 178.545 209.410 178.560 ;
        RECT 229.780 178.545 230.110 178.560 ;
        RECT 159.185 93.465 159.485 178.410 ;
        RECT 165.380 178.180 165.710 178.195 ;
        RECT 173.660 178.180 173.990 178.195 ;
        RECT 191.140 178.180 191.470 178.195 ;
        RECT 165.380 177.880 173.990 178.180 ;
        RECT 165.380 177.865 165.710 177.880 ;
        RECT 173.660 177.865 173.990 177.880 ;
        RECT 174.365 177.880 191.470 178.180 ;
        RECT 164.000 177.500 164.330 177.515 ;
        RECT 170.900 177.500 171.230 177.515 ;
        RECT 164.000 177.200 171.230 177.500 ;
        RECT 164.000 177.185 164.330 177.200 ;
        RECT 170.900 177.185 171.230 177.200 ;
        RECT 172.280 177.500 172.610 177.515 ;
        RECT 174.365 177.500 174.665 177.880 ;
        RECT 191.140 177.865 191.470 177.880 ;
        RECT 214.140 178.180 214.470 178.195 ;
        RECT 215.980 178.180 216.310 178.195 ;
        RECT 214.140 177.880 216.310 178.180 ;
        RECT 214.140 177.865 214.470 177.880 ;
        RECT 215.980 177.865 216.310 177.880 ;
        RECT 219.660 178.180 219.990 178.195 ;
        RECT 227.940 178.180 228.270 178.195 ;
        RECT 219.660 177.880 228.270 178.180 ;
        RECT 219.660 177.865 219.990 177.880 ;
        RECT 227.940 177.865 228.270 177.880 ;
        RECT 172.280 177.200 174.665 177.500 ;
        RECT 210.920 177.500 211.250 177.515 ;
        RECT 220.120 177.500 220.450 177.515 ;
        RECT 210.920 177.200 220.450 177.500 ;
        RECT 172.280 177.185 172.610 177.200 ;
        RECT 210.920 177.185 211.250 177.200 ;
        RECT 220.120 177.185 220.450 177.200 ;
        RECT 180.925 176.845 182.505 177.175 ;
        RECT 220.925 176.845 222.505 177.175 ;
        RECT 169.520 176.820 169.850 176.835 ;
        RECT 179.180 176.820 179.510 176.835 ;
        RECT 169.520 176.520 179.510 176.820 ;
        RECT 169.520 176.505 169.850 176.520 ;
        RECT 179.180 176.505 179.510 176.520 ;
        RECT 182.860 176.820 183.190 176.835 ;
        RECT 184.240 176.820 184.570 176.835 ;
        RECT 182.860 176.520 184.570 176.820 ;
        RECT 182.860 176.505 183.190 176.520 ;
        RECT 184.240 176.505 184.570 176.520 ;
        RECT 222.880 176.820 223.210 176.835 ;
        RECT 234.380 176.820 234.710 176.835 ;
        RECT 222.880 176.520 234.710 176.820 ;
        RECT 222.880 176.505 223.210 176.520 ;
        RECT 234.380 176.505 234.710 176.520 ;
        RECT 182.400 176.140 182.730 176.155 ;
        RECT 183.320 176.140 183.650 176.155 ;
        RECT 182.400 175.840 183.650 176.140 ;
        RECT 182.400 175.825 182.730 175.840 ;
        RECT 183.320 175.825 183.650 175.840 ;
        RECT 221.960 176.140 222.290 176.155 ;
        RECT 230.240 176.140 230.570 176.155 ;
        RECT 221.960 175.840 230.570 176.140 ;
        RECT 221.960 175.825 222.290 175.840 ;
        RECT 230.240 175.825 230.570 175.840 ;
        RECT 186.285 175.460 186.665 175.470 ;
        RECT 223.085 175.460 223.465 175.470 ;
        RECT 186.285 175.160 223.465 175.460 ;
        RECT 186.285 175.150 186.665 175.160 ;
        RECT 223.085 175.150 223.465 175.160 ;
        RECT 207.445 174.780 207.825 174.790 ;
        RECT 233.000 174.780 233.330 174.795 ;
        RECT 207.445 174.480 233.330 174.780 ;
        RECT 207.445 174.470 207.825 174.480 ;
        RECT 233.000 174.465 233.330 174.480 ;
        RECT 246.665 152.705 246.965 217.650 ;
        RECT 247.985 153.875 248.285 219.960 ;
        RECT 249.070 154.925 249.370 220.560 ;
        RECT 249.920 155.950 250.220 221.160 ;
        RECT 250.925 157.080 251.225 224.750 ;
        RECT 251.860 158.175 252.160 225.410 ;
        RECT 251.860 157.875 318.785 158.175 ;
        RECT 250.925 156.780 317.675 157.080 ;
        RECT 249.920 155.650 316.845 155.950 ;
        RECT 249.070 154.625 316.145 154.925 ;
        RECT 247.985 153.575 315.370 153.875 ;
        RECT 246.665 152.405 314.635 152.705 ;
        RECT 180.915 121.980 302.515 123.580 ;
        RECT 177.615 119.175 299.215 120.775 ;
        RECT 180.925 106.260 182.505 106.590 ;
        RECT 220.925 106.260 222.505 106.590 ;
        RECT 260.925 106.260 262.505 106.590 ;
        RECT 300.925 106.260 302.505 106.590 ;
        RECT 247.260 104.195 247.590 104.210 ;
        RECT 256.000 104.195 256.330 104.210 ;
        RECT 247.260 103.895 256.330 104.195 ;
        RECT 247.260 103.880 247.590 103.895 ;
        RECT 256.000 103.880 256.330 103.895 ;
        RECT 177.625 103.540 179.205 103.870 ;
        RECT 217.625 103.540 219.205 103.870 ;
        RECT 257.625 103.540 259.205 103.870 ;
        RECT 297.625 103.540 299.205 103.870 ;
        RECT 314.335 101.625 314.635 152.405 ;
        RECT 308.900 101.475 309.230 101.490 ;
        RECT 312.335 101.475 314.635 101.625 ;
        RECT 308.900 101.175 314.635 101.475 ;
        RECT 308.900 101.160 309.230 101.175 ;
        RECT 180.925 100.820 182.505 101.150 ;
        RECT 220.925 100.820 222.505 101.150 ;
        RECT 260.925 100.820 262.505 101.150 ;
        RECT 300.925 100.820 302.505 101.150 ;
        RECT 312.335 101.025 314.635 101.175 ;
        RECT 207.700 100.115 208.030 100.130 ;
        RECT 221.040 100.115 221.370 100.130 ;
        RECT 223.800 100.115 224.130 100.130 ;
        RECT 207.700 99.815 224.130 100.115 ;
        RECT 207.700 99.800 208.030 99.815 ;
        RECT 221.040 99.800 221.370 99.815 ;
        RECT 223.800 99.800 224.130 99.815 ;
        RECT 229.320 100.115 229.650 100.130 ;
        RECT 260.600 100.115 260.930 100.130 ;
        RECT 229.320 99.815 260.930 100.115 ;
        RECT 229.320 99.800 229.650 99.815 ;
        RECT 260.600 99.800 260.930 99.815 ;
        RECT 173.660 99.435 173.990 99.450 ;
        RECT 175.960 99.435 176.290 99.450 ;
        RECT 228.400 99.435 228.730 99.450 ;
        RECT 173.660 99.135 228.730 99.435 ;
        RECT 173.660 99.120 173.990 99.135 ;
        RECT 175.960 99.120 176.290 99.135 ;
        RECT 228.400 99.120 228.730 99.135 ;
        RECT 230.240 99.435 230.570 99.450 ;
        RECT 250.020 99.435 250.350 99.450 ;
        RECT 230.240 99.135 250.350 99.435 ;
        RECT 230.240 99.120 230.570 99.135 ;
        RECT 250.020 99.120 250.350 99.135 ;
        RECT 232.540 98.755 232.870 98.770 ;
        RECT 250.940 98.755 251.270 98.770 ;
        RECT 232.540 98.455 251.270 98.755 ;
        RECT 232.540 98.440 232.870 98.455 ;
        RECT 250.940 98.440 251.270 98.455 ;
        RECT 177.625 98.100 179.205 98.430 ;
        RECT 217.625 98.100 219.205 98.430 ;
        RECT 257.625 98.100 259.205 98.430 ;
        RECT 297.625 98.100 299.205 98.430 ;
        RECT 221.500 98.075 221.830 98.090 ;
        RECT 221.500 97.775 256.085 98.075 ;
        RECT 221.500 97.760 221.830 97.775 ;
        RECT 203.560 97.395 203.890 97.410 ;
        RECT 243.120 97.395 243.450 97.410 ;
        RECT 203.560 97.095 243.450 97.395 ;
        RECT 255.785 97.395 256.085 97.775 ;
        RECT 257.380 97.395 257.710 97.410 ;
        RECT 278.080 97.395 278.410 97.410 ;
        RECT 255.785 97.095 278.410 97.395 ;
        RECT 203.560 97.080 203.890 97.095 ;
        RECT 243.120 97.080 243.450 97.095 ;
        RECT 257.380 97.080 257.710 97.095 ;
        RECT 278.080 97.080 278.410 97.095 ;
        RECT 182.400 96.715 182.730 96.730 ;
        RECT 187.000 96.715 187.330 96.730 ;
        RECT 193.440 96.715 193.770 96.730 ;
        RECT 182.400 96.415 193.770 96.715 ;
        RECT 182.400 96.400 182.730 96.415 ;
        RECT 187.000 96.400 187.330 96.415 ;
        RECT 193.440 96.400 193.770 96.415 ;
        RECT 196.660 96.715 196.990 96.730 ;
        RECT 222.880 96.715 223.210 96.730 ;
        RECT 260.140 96.715 260.470 96.730 ;
        RECT 278.540 96.715 278.870 96.730 ;
        RECT 196.660 96.415 278.870 96.715 ;
        RECT 196.660 96.400 196.990 96.415 ;
        RECT 222.880 96.400 223.210 96.415 ;
        RECT 260.140 96.400 260.470 96.415 ;
        RECT 278.540 96.400 278.870 96.415 ;
        RECT 285.440 96.715 285.770 96.730 ;
        RECT 306.600 96.715 306.930 96.730 ;
        RECT 285.440 96.415 306.930 96.715 ;
        RECT 285.440 96.400 285.770 96.415 ;
        RECT 306.600 96.400 306.930 96.415 ;
        RECT 247.720 96.035 248.050 96.050 ;
        RECT 253.240 96.035 253.570 96.050 ;
        RECT 247.720 95.735 253.570 96.035 ;
        RECT 247.720 95.720 248.050 95.735 ;
        RECT 253.240 95.720 253.570 95.735 ;
        RECT 180.925 95.380 182.505 95.710 ;
        RECT 220.925 95.380 222.505 95.710 ;
        RECT 260.925 95.380 262.505 95.710 ;
        RECT 300.925 95.380 302.505 95.710 ;
        RECT 195.280 94.675 195.610 94.690 ;
        RECT 242.660 94.675 242.990 94.690 ;
        RECT 195.280 94.375 242.990 94.675 ;
        RECT 195.280 94.360 195.610 94.375 ;
        RECT 242.660 94.360 242.990 94.375 ;
        RECT 256.205 94.675 256.585 94.685 ;
        RECT 257.380 94.675 257.710 94.690 ;
        RECT 276.700 94.675 277.030 94.690 ;
        RECT 256.205 94.375 277.030 94.675 ;
        RECT 256.205 94.365 256.585 94.375 ;
        RECT 257.380 94.360 257.710 94.375 ;
        RECT 276.700 94.360 277.030 94.375 ;
        RECT 193.900 93.995 194.230 94.010 ;
        RECT 260.140 93.995 260.470 94.010 ;
        RECT 193.900 93.695 260.470 93.995 ;
        RECT 193.900 93.680 194.230 93.695 ;
        RECT 260.140 93.680 260.470 93.695 ;
        RECT 159.185 93.315 161.335 93.465 ;
        RECT 164.000 93.315 164.330 93.330 ;
        RECT 159.185 93.015 164.330 93.315 ;
        RECT 159.185 92.865 161.335 93.015 ;
        RECT 164.000 93.000 164.330 93.015 ;
        RECT 177.625 92.660 179.205 92.990 ;
        RECT 217.625 92.660 219.205 92.990 ;
        RECT 257.625 92.660 259.205 92.990 ;
        RECT 297.625 92.660 299.205 92.990 ;
        RECT 263.820 92.645 264.150 92.650 ;
        RECT 263.565 92.635 264.150 92.645 ;
        RECT 263.365 92.335 264.150 92.635 ;
        RECT 263.565 92.325 264.150 92.335 ;
        RECT 263.820 92.320 264.150 92.325 ;
        RECT 211.380 91.955 211.710 91.970 ;
        RECT 248.180 91.955 248.510 91.970 ;
        RECT 211.380 91.655 248.510 91.955 ;
        RECT 211.380 91.640 211.710 91.655 ;
        RECT 248.180 91.640 248.510 91.655 ;
        RECT 250.940 91.955 251.270 91.970 ;
        RECT 303.840 91.955 304.170 91.970 ;
        RECT 250.940 91.655 304.170 91.955 ;
        RECT 250.940 91.640 251.270 91.655 ;
        RECT 303.840 91.640 304.170 91.655 ;
        RECT 200.800 91.275 201.130 91.290 ;
        RECT 231.160 91.275 231.490 91.290 ;
        RECT 200.800 90.975 231.490 91.275 ;
        RECT 200.800 90.960 201.130 90.975 ;
        RECT 231.160 90.960 231.490 90.975 ;
        RECT 242.660 91.275 242.990 91.290 ;
        RECT 245.880 91.275 246.210 91.290 ;
        RECT 247.260 91.275 247.590 91.290 ;
        RECT 242.660 90.975 247.590 91.275 ;
        RECT 242.660 90.960 242.990 90.975 ;
        RECT 245.880 90.960 246.210 90.975 ;
        RECT 247.260 90.960 247.590 90.975 ;
        RECT 258.300 91.275 258.630 91.290 ;
        RECT 265.200 91.275 265.530 91.290 ;
        RECT 288.660 91.275 288.990 91.290 ;
        RECT 258.300 90.975 264.825 91.275 ;
        RECT 258.300 90.960 258.630 90.975 ;
        RECT 264.525 90.595 264.825 90.975 ;
        RECT 265.200 90.975 288.990 91.275 ;
        RECT 265.200 90.960 265.530 90.975 ;
        RECT 288.660 90.960 288.990 90.975 ;
        RECT 285.440 90.595 285.770 90.610 ;
        RECT 264.525 90.295 285.770 90.595 ;
        RECT 285.440 90.280 285.770 90.295 ;
        RECT 180.925 89.940 182.505 90.270 ;
        RECT 220.925 89.940 222.505 90.270 ;
        RECT 260.925 89.940 262.505 90.270 ;
        RECT 300.925 89.940 302.505 90.270 ;
        RECT 259.680 89.915 260.010 89.930 ;
        RECT 225.885 89.615 260.010 89.915 ;
        RECT 183.780 89.235 184.110 89.250 ;
        RECT 225.885 89.235 226.185 89.615 ;
        RECT 259.680 89.600 260.010 89.615 ;
        RECT 183.780 88.935 226.185 89.235 ;
        RECT 226.560 89.235 226.890 89.250 ;
        RECT 277.620 89.235 277.950 89.250 ;
        RECT 226.560 88.935 277.950 89.235 ;
        RECT 183.780 88.920 184.110 88.935 ;
        RECT 226.560 88.920 226.890 88.935 ;
        RECT 277.620 88.920 277.950 88.935 ;
        RECT 213.220 88.555 213.550 88.570 ;
        RECT 268.880 88.555 269.210 88.570 ;
        RECT 213.220 88.255 269.210 88.555 ;
        RECT 213.220 88.240 213.550 88.255 ;
        RECT 268.880 88.240 269.210 88.255 ;
        RECT 244.500 87.875 244.830 87.890 ;
        RECT 253.700 87.875 254.030 87.890 ;
        RECT 256.920 87.875 257.250 87.890 ;
        RECT 244.500 87.575 257.250 87.875 ;
        RECT 244.500 87.560 244.830 87.575 ;
        RECT 253.700 87.560 254.030 87.575 ;
        RECT 256.920 87.560 257.250 87.575 ;
        RECT 177.625 87.220 179.205 87.550 ;
        RECT 217.625 87.220 219.205 87.550 ;
        RECT 257.625 87.220 259.205 87.550 ;
        RECT 297.625 87.220 299.205 87.550 ;
        RECT 259.680 87.205 260.010 87.210 ;
        RECT 259.680 87.195 260.265 87.205 ;
        RECT 259.680 86.895 260.465 87.195 ;
        RECT 259.680 86.885 260.265 86.895 ;
        RECT 259.680 86.880 260.010 86.885 ;
        RECT 211.840 86.515 212.170 86.530 ;
        RECT 234.380 86.515 234.710 86.530 ;
        RECT 211.840 86.215 234.710 86.515 ;
        RECT 211.840 86.200 212.170 86.215 ;
        RECT 234.380 86.200 234.710 86.215 ;
        RECT 309.360 85.155 309.690 85.170 ;
        RECT 312.335 85.155 314.335 85.305 ;
        RECT 309.360 85.145 314.335 85.155 ;
        RECT 315.070 85.145 315.370 153.575 ;
        RECT 309.360 84.855 315.370 85.145 ;
        RECT 309.360 84.840 309.690 84.855 ;
        RECT 312.335 84.845 315.370 84.855 ;
        RECT 180.925 84.500 182.505 84.830 ;
        RECT 220.925 84.500 222.505 84.830 ;
        RECT 260.925 84.500 262.505 84.830 ;
        RECT 300.925 84.500 302.505 84.830 ;
        RECT 312.335 84.705 314.335 84.845 ;
        RECT 216.440 83.795 216.770 83.810 ;
        RECT 228.400 83.795 228.730 83.810 ;
        RECT 216.440 83.495 228.730 83.795 ;
        RECT 216.440 83.480 216.770 83.495 ;
        RECT 228.400 83.480 228.730 83.495 ;
        RECT 238.060 83.795 238.390 83.810 ;
        RECT 244.960 83.795 245.290 83.810 ;
        RECT 285.900 83.795 286.230 83.810 ;
        RECT 304.760 83.795 305.090 83.810 ;
        RECT 238.060 83.495 305.090 83.795 ;
        RECT 238.060 83.480 238.390 83.495 ;
        RECT 244.960 83.480 245.290 83.495 ;
        RECT 285.900 83.480 286.230 83.495 ;
        RECT 304.760 83.480 305.090 83.495 ;
        RECT 197.580 83.115 197.910 83.130 ;
        RECT 269.340 83.115 269.670 83.130 ;
        RECT 197.580 82.815 269.670 83.115 ;
        RECT 197.580 82.800 197.910 82.815 ;
        RECT 269.340 82.800 269.670 82.815 ;
        RECT 241.740 82.435 242.070 82.450 ;
        RECT 252.780 82.435 253.110 82.450 ;
        RECT 241.740 82.135 253.110 82.435 ;
        RECT 241.740 82.120 242.070 82.135 ;
        RECT 252.780 82.120 253.110 82.135 ;
        RECT 177.625 81.780 179.205 82.110 ;
        RECT 217.625 81.780 219.205 82.110 ;
        RECT 257.625 81.780 259.205 82.110 ;
        RECT 297.625 81.780 299.205 82.110 ;
        RECT 229.320 81.755 229.650 81.770 ;
        RECT 247.260 81.755 247.590 81.770 ;
        RECT 229.320 81.455 247.590 81.755 ;
        RECT 229.320 81.440 229.650 81.455 ;
        RECT 247.260 81.440 247.590 81.455 ;
        RECT 261.980 81.755 262.310 81.770 ;
        RECT 263.820 81.755 264.150 81.770 ;
        RECT 267.960 81.755 268.290 81.770 ;
        RECT 261.980 81.455 268.290 81.755 ;
        RECT 261.980 81.440 262.310 81.455 ;
        RECT 263.820 81.440 264.150 81.455 ;
        RECT 267.960 81.440 268.290 81.455 ;
        RECT 212.300 81.075 212.630 81.090 ;
        RECT 241.740 81.075 242.070 81.090 ;
        RECT 249.560 81.075 249.890 81.090 ;
        RECT 212.300 80.775 222.505 81.075 ;
        RECT 212.300 80.760 212.630 80.775 ;
        RECT 212.760 80.395 213.090 80.410 ;
        RECT 217.360 80.395 217.690 80.410 ;
        RECT 212.760 80.095 217.690 80.395 ;
        RECT 222.205 80.395 222.505 80.775 ;
        RECT 241.740 80.775 249.890 81.075 ;
        RECT 241.740 80.760 242.070 80.775 ;
        RECT 249.560 80.760 249.890 80.775 ;
        RECT 261.520 81.075 261.850 81.090 ;
        RECT 262.900 81.075 263.230 81.090 ;
        RECT 265.200 81.075 265.530 81.090 ;
        RECT 261.520 80.775 265.530 81.075 ;
        RECT 261.520 80.760 261.850 80.775 ;
        RECT 262.900 80.760 263.230 80.775 ;
        RECT 265.200 80.760 265.530 80.775 ;
        RECT 229.780 80.395 230.110 80.410 ;
        RECT 222.205 80.095 230.110 80.395 ;
        RECT 212.760 80.080 213.090 80.095 ;
        RECT 217.360 80.080 217.690 80.095 ;
        RECT 229.780 80.080 230.110 80.095 ;
        RECT 248.640 80.405 248.970 80.410 ;
        RECT 248.640 80.395 249.225 80.405 ;
        RECT 264.280 80.395 264.610 80.410 ;
        RECT 269.340 80.395 269.670 80.410 ;
        RECT 291.420 80.395 291.750 80.410 ;
        RECT 248.640 80.095 249.425 80.395 ;
        RECT 264.280 80.095 291.750 80.395 ;
        RECT 248.640 80.085 249.225 80.095 ;
        RECT 248.640 80.080 248.970 80.085 ;
        RECT 264.280 80.080 264.610 80.095 ;
        RECT 269.340 80.080 269.670 80.095 ;
        RECT 291.420 80.080 291.750 80.095 ;
        RECT 227.020 79.715 227.350 79.730 ;
        RECT 246.800 79.715 247.130 79.730 ;
        RECT 249.560 79.715 249.890 79.730 ;
        RECT 227.020 79.415 249.890 79.715 ;
        RECT 227.020 79.400 227.350 79.415 ;
        RECT 246.800 79.400 247.130 79.415 ;
        RECT 249.560 79.400 249.890 79.415 ;
        RECT 180.925 79.060 182.505 79.390 ;
        RECT 220.925 79.060 222.505 79.390 ;
        RECT 260.925 79.060 262.505 79.390 ;
        RECT 300.925 79.060 302.505 79.390 ;
        RECT 213.680 79.035 214.010 79.050 ;
        RECT 217.820 79.035 218.150 79.050 ;
        RECT 213.680 78.735 218.150 79.035 ;
        RECT 213.680 78.720 214.010 78.735 ;
        RECT 217.820 78.720 218.150 78.735 ;
        RECT 230.700 79.035 231.030 79.050 ;
        RECT 248.180 79.035 248.510 79.050 ;
        RECT 230.700 78.735 248.510 79.035 ;
        RECT 230.700 78.720 231.030 78.735 ;
        RECT 248.180 78.720 248.510 78.735 ;
        RECT 179.640 78.355 179.970 78.370 ;
        RECT 256.460 78.355 256.790 78.370 ;
        RECT 179.640 78.055 256.790 78.355 ;
        RECT 179.640 78.040 179.970 78.055 ;
        RECT 256.460 78.040 256.790 78.055 ;
        RECT 258.300 78.355 258.630 78.370 ;
        RECT 259.885 78.355 260.265 78.365 ;
        RECT 266.580 78.355 266.910 78.370 ;
        RECT 258.300 78.055 266.910 78.355 ;
        RECT 258.300 78.040 258.630 78.055 ;
        RECT 259.885 78.045 260.265 78.055 ;
        RECT 266.580 78.040 266.910 78.055 ;
        RECT 185.620 77.675 185.950 77.690 ;
        RECT 259.220 77.675 259.550 77.690 ;
        RECT 259.885 77.675 260.265 77.685 ;
        RECT 185.620 77.375 260.265 77.675 ;
        RECT 185.620 77.360 185.950 77.375 ;
        RECT 259.220 77.360 259.550 77.375 ;
        RECT 259.885 77.365 260.265 77.375 ;
        RECT 260.600 77.675 260.930 77.690 ;
        RECT 263.820 77.675 264.150 77.690 ;
        RECT 260.600 77.375 264.150 77.675 ;
        RECT 260.600 77.360 260.930 77.375 ;
        RECT 263.820 77.360 264.150 77.375 ;
        RECT 177.625 76.340 179.205 76.670 ;
        RECT 217.625 76.340 219.205 76.670 ;
        RECT 257.625 76.340 259.205 76.670 ;
        RECT 297.625 76.340 299.205 76.670 ;
        RECT 259.680 76.000 260.010 76.330 ;
        RECT 261.980 76.315 262.310 76.330 ;
        RECT 264.280 76.315 264.610 76.330 ;
        RECT 261.980 76.015 264.610 76.315 ;
        RECT 261.980 76.000 262.310 76.015 ;
        RECT 264.280 76.000 264.610 76.015 ;
        RECT 184.240 75.635 184.570 75.650 ;
        RECT 186.080 75.635 186.410 75.650 ;
        RECT 184.240 75.335 186.410 75.635 ;
        RECT 184.240 75.320 184.570 75.335 ;
        RECT 186.080 75.320 186.410 75.335 ;
        RECT 214.140 75.635 214.470 75.650 ;
        RECT 259.695 75.635 259.995 76.000 ;
        RECT 261.520 75.635 261.850 75.650 ;
        RECT 214.140 75.335 261.850 75.635 ;
        RECT 214.140 75.320 214.470 75.335 ;
        RECT 261.520 75.320 261.850 75.335 ;
        RECT 212.300 74.955 212.630 74.970 ;
        RECT 253.700 74.955 254.030 74.970 ;
        RECT 212.300 74.655 254.030 74.955 ;
        RECT 212.300 74.640 212.630 74.655 ;
        RECT 253.700 74.640 254.030 74.655 ;
        RECT 255.080 74.955 255.410 74.970 ;
        RECT 265.200 74.955 265.530 74.970 ;
        RECT 255.080 74.655 265.530 74.955 ;
        RECT 255.080 74.640 255.410 74.655 ;
        RECT 265.200 74.640 265.530 74.655 ;
        RECT 257.840 74.275 258.170 74.290 ;
        RECT 259.680 74.275 260.010 74.290 ;
        RECT 257.840 73.975 260.010 74.275 ;
        RECT 257.840 73.960 258.170 73.975 ;
        RECT 259.680 73.960 260.010 73.975 ;
        RECT 180.925 73.620 182.505 73.950 ;
        RECT 220.925 73.620 222.505 73.950 ;
        RECT 260.925 73.620 262.505 73.950 ;
        RECT 300.925 73.620 302.505 73.950 ;
        RECT 172.740 73.595 173.070 73.610 ;
        RECT 175.040 73.595 175.370 73.610 ;
        RECT 172.740 73.295 175.370 73.595 ;
        RECT 172.740 73.280 173.070 73.295 ;
        RECT 175.040 73.280 175.370 73.295 ;
        RECT 182.860 73.595 183.190 73.610 ;
        RECT 203.100 73.595 203.430 73.610 ;
        RECT 182.860 73.295 203.430 73.595 ;
        RECT 182.860 73.280 183.190 73.295 ;
        RECT 203.100 73.280 203.430 73.295 ;
        RECT 257.380 73.595 257.710 73.610 ;
        RECT 259.885 73.595 260.265 73.605 ;
        RECT 257.380 73.295 260.265 73.595 ;
        RECT 257.380 73.280 257.710 73.295 ;
        RECT 259.885 73.285 260.265 73.295 ;
        RECT 184.700 72.915 185.030 72.930 ;
        RECT 216.440 72.915 216.770 72.930 ;
        RECT 220.120 72.915 220.450 72.930 ;
        RECT 184.700 72.615 220.450 72.915 ;
        RECT 184.700 72.600 185.030 72.615 ;
        RECT 216.440 72.600 216.770 72.615 ;
        RECT 220.120 72.600 220.450 72.615 ;
        RECT 256.205 72.915 256.585 72.925 ;
        RECT 261.520 72.915 261.850 72.930 ;
        RECT 256.205 72.615 261.850 72.915 ;
        RECT 256.205 72.605 256.585 72.615 ;
        RECT 261.520 72.600 261.850 72.615 ;
        RECT 262.440 72.915 262.770 72.930 ;
        RECT 268.880 72.915 269.210 72.930 ;
        RECT 262.440 72.615 269.210 72.915 ;
        RECT 262.440 72.600 262.770 72.615 ;
        RECT 268.880 72.600 269.210 72.615 ;
        RECT 227.940 72.235 228.270 72.250 ;
        RECT 262.455 72.235 262.755 72.600 ;
        RECT 227.940 71.935 262.755 72.235 ;
        RECT 227.940 71.920 228.270 71.935 ;
        RECT 177.625 70.900 179.205 71.230 ;
        RECT 217.625 70.900 219.205 71.230 ;
        RECT 257.625 70.900 259.205 71.230 ;
        RECT 297.625 70.900 299.205 71.230 ;
        RECT 179.640 70.875 179.970 70.890 ;
        RECT 234.380 70.875 234.710 70.890 ;
        RECT 256.205 70.875 256.585 70.885 ;
        RECT 256.920 70.875 257.250 70.890 ;
        RECT 179.640 70.560 180.185 70.875 ;
        RECT 234.380 70.575 248.265 70.875 ;
        RECT 234.380 70.560 234.710 70.575 ;
        RECT 179.885 70.195 180.185 70.560 ;
        RECT 242.660 70.195 242.990 70.210 ;
        RECT 246.800 70.195 247.130 70.210 ;
        RECT 179.885 69.895 247.130 70.195 ;
        RECT 247.965 70.195 248.265 70.575 ;
        RECT 256.205 70.575 257.250 70.875 ;
        RECT 256.205 70.565 256.585 70.575 ;
        RECT 256.920 70.560 257.250 70.575 ;
        RECT 261.520 70.875 261.850 70.890 ;
        RECT 263.565 70.875 263.945 70.885 ;
        RECT 261.520 70.575 263.945 70.875 ;
        RECT 261.520 70.560 261.850 70.575 ;
        RECT 263.565 70.565 263.945 70.575 ;
        RECT 296.480 70.195 296.810 70.210 ;
        RECT 247.965 69.895 296.810 70.195 ;
        RECT 242.660 69.880 242.990 69.895 ;
        RECT 246.800 69.880 247.130 69.895 ;
        RECT 296.480 69.880 296.810 69.895 ;
        RECT 175.960 69.515 176.290 69.530 ;
        RECT 207.700 69.515 208.030 69.530 ;
        RECT 247.720 69.515 248.050 69.530 ;
        RECT 250.940 69.515 251.270 69.530 ;
        RECT 175.960 69.215 203.415 69.515 ;
        RECT 175.960 69.200 176.290 69.215 ;
        RECT 203.115 68.850 203.415 69.215 ;
        RECT 207.700 69.215 247.345 69.515 ;
        RECT 207.700 69.200 208.030 69.215 ;
        RECT 203.100 68.835 203.430 68.850 ;
        RECT 219.660 68.835 219.990 68.850 ;
        RECT 203.100 68.535 219.990 68.835 ;
        RECT 247.045 68.835 247.345 69.215 ;
        RECT 247.720 69.215 263.905 69.515 ;
        RECT 247.720 69.200 248.050 69.215 ;
        RECT 250.940 69.200 251.270 69.215 ;
        RECT 250.020 68.835 250.350 68.850 ;
        RECT 247.045 68.535 250.350 68.835 ;
        RECT 263.605 68.835 263.905 69.215 ;
        RECT 279.000 68.835 279.330 68.850 ;
        RECT 293.260 68.835 293.590 68.850 ;
        RECT 263.605 68.535 293.590 68.835 ;
        RECT 203.100 68.520 203.430 68.535 ;
        RECT 219.660 68.520 219.990 68.535 ;
        RECT 250.020 68.520 250.350 68.535 ;
        RECT 279.000 68.520 279.330 68.535 ;
        RECT 293.260 68.520 293.590 68.535 ;
        RECT 309.360 68.835 309.690 68.850 ;
        RECT 312.335 68.835 314.335 68.985 ;
        RECT 309.360 68.820 314.335 68.835 ;
        RECT 315.845 68.820 316.145 154.625 ;
        RECT 309.360 68.535 316.145 68.820 ;
        RECT 309.360 68.520 309.690 68.535 ;
        RECT 312.335 68.520 316.145 68.535 ;
        RECT 180.925 68.180 182.505 68.510 ;
        RECT 220.925 68.180 222.505 68.510 ;
        RECT 260.925 68.180 262.505 68.510 ;
        RECT 300.925 68.180 302.505 68.510 ;
        RECT 312.335 68.385 314.335 68.520 ;
        RECT 192.520 68.155 192.850 68.170 ;
        RECT 206.320 68.155 206.650 68.170 ;
        RECT 192.520 67.855 206.650 68.155 ;
        RECT 192.520 67.840 192.850 67.855 ;
        RECT 206.320 67.840 206.650 67.855 ;
        RECT 212.760 68.155 213.090 68.170 ;
        RECT 217.820 68.155 218.150 68.170 ;
        RECT 212.760 67.855 218.150 68.155 ;
        RECT 212.760 67.840 213.090 67.855 ;
        RECT 217.820 67.840 218.150 67.855 ;
        RECT 240.360 68.155 240.690 68.170 ;
        RECT 299.700 68.155 300.030 68.170 ;
        RECT 240.360 67.855 260.225 68.155 ;
        RECT 240.360 67.840 240.690 67.855 ;
        RECT 172.280 67.475 172.610 67.490 ;
        RECT 207.700 67.475 208.030 67.490 ;
        RECT 218.280 67.475 218.610 67.490 ;
        RECT 259.220 67.475 259.550 67.490 ;
        RECT 172.280 67.175 218.610 67.475 ;
        RECT 172.280 67.160 172.610 67.175 ;
        RECT 207.700 67.160 208.030 67.175 ;
        RECT 218.280 67.160 218.610 67.175 ;
        RECT 221.285 67.175 259.550 67.475 ;
        RECT 259.925 67.475 260.225 67.855 ;
        RECT 269.585 67.855 300.030 68.155 ;
        RECT 269.585 67.475 269.885 67.855 ;
        RECT 299.700 67.840 300.030 67.855 ;
        RECT 259.925 67.175 269.885 67.475 ;
        RECT 199.880 66.795 200.210 66.810 ;
        RECT 204.480 66.795 204.810 66.810 ;
        RECT 221.285 66.795 221.585 67.175 ;
        RECT 259.220 67.160 259.550 67.175 ;
        RECT 199.880 66.495 221.585 66.795 ;
        RECT 248.640 66.805 248.970 66.810 ;
        RECT 248.640 66.795 249.225 66.805 ;
        RECT 257.840 66.795 258.170 66.810 ;
        RECT 264.280 66.795 264.610 66.810 ;
        RECT 248.640 66.495 249.425 66.795 ;
        RECT 257.840 66.495 264.610 66.795 ;
        RECT 199.880 66.480 200.210 66.495 ;
        RECT 204.480 66.480 204.810 66.495 ;
        RECT 248.640 66.485 249.225 66.495 ;
        RECT 248.640 66.480 248.970 66.485 ;
        RECT 257.840 66.480 258.170 66.495 ;
        RECT 264.280 66.480 264.610 66.495 ;
        RECT 279.460 66.795 279.790 66.810 ;
        RECT 293.720 66.795 294.050 66.810 ;
        RECT 279.460 66.495 294.050 66.795 ;
        RECT 279.460 66.480 279.790 66.495 ;
        RECT 293.720 66.480 294.050 66.495 ;
        RECT 177.625 65.460 179.205 65.790 ;
        RECT 217.625 65.460 219.205 65.790 ;
        RECT 257.625 65.460 259.205 65.790 ;
        RECT 297.625 65.460 299.205 65.790 ;
        RECT 208.160 65.435 208.490 65.450 ;
        RECT 215.520 65.435 215.850 65.450 ;
        RECT 208.160 65.135 215.850 65.435 ;
        RECT 208.160 65.120 208.490 65.135 ;
        RECT 215.520 65.120 215.850 65.135 ;
        RECT 243.580 65.435 243.910 65.450 ;
        RECT 243.580 65.135 256.085 65.435 ;
        RECT 243.580 65.120 243.910 65.135 ;
        RECT 192.520 64.755 192.850 64.770 ;
        RECT 196.200 64.755 196.530 64.770 ;
        RECT 245.420 64.755 245.750 64.770 ;
        RECT 192.520 64.455 245.750 64.755 ;
        RECT 255.785 64.755 256.085 65.135 ;
        RECT 287.740 64.755 288.070 64.770 ;
        RECT 255.785 64.455 288.070 64.755 ;
        RECT 192.520 64.440 192.850 64.455 ;
        RECT 196.200 64.440 196.530 64.455 ;
        RECT 245.420 64.440 245.750 64.455 ;
        RECT 287.740 64.440 288.070 64.455 ;
        RECT 179.640 64.075 179.970 64.090 ;
        RECT 187.000 64.075 187.330 64.090 ;
        RECT 179.640 63.775 187.330 64.075 ;
        RECT 179.640 63.760 179.970 63.775 ;
        RECT 187.000 63.760 187.330 63.775 ;
        RECT 193.900 64.075 194.230 64.090 ;
        RECT 197.120 64.075 197.450 64.090 ;
        RECT 259.220 64.075 259.550 64.090 ;
        RECT 193.900 63.775 259.550 64.075 ;
        RECT 193.900 63.760 194.230 63.775 ;
        RECT 197.120 63.760 197.450 63.775 ;
        RECT 259.220 63.760 259.550 63.775 ;
        RECT 213.680 63.395 214.010 63.410 ;
        RECT 217.360 63.395 217.690 63.410 ;
        RECT 213.680 63.095 217.690 63.395 ;
        RECT 213.680 63.080 214.010 63.095 ;
        RECT 217.360 63.080 217.690 63.095 ;
        RECT 180.925 62.740 182.505 63.070 ;
        RECT 220.925 62.740 222.505 63.070 ;
        RECT 260.925 62.740 262.505 63.070 ;
        RECT 300.925 62.740 302.505 63.070 ;
        RECT 211.380 62.035 211.710 62.050 ;
        RECT 248.640 62.035 248.970 62.050 ;
        RECT 211.380 61.735 248.970 62.035 ;
        RECT 211.380 61.720 211.710 61.735 ;
        RECT 248.640 61.720 248.970 61.735 ;
        RECT 253.700 62.035 254.030 62.050 ;
        RECT 284.060 62.035 284.390 62.050 ;
        RECT 253.700 61.735 284.390 62.035 ;
        RECT 253.700 61.720 254.030 61.735 ;
        RECT 284.060 61.720 284.390 61.735 ;
        RECT 193.440 61.355 193.770 61.370 ;
        RECT 255.540 61.355 255.870 61.370 ;
        RECT 193.440 61.055 255.870 61.355 ;
        RECT 193.440 61.040 193.770 61.055 ;
        RECT 255.540 61.040 255.870 61.055 ;
        RECT 262.440 61.355 262.770 61.370 ;
        RECT 282.220 61.355 282.550 61.370 ;
        RECT 262.440 61.055 282.550 61.355 ;
        RECT 262.440 61.040 262.770 61.055 ;
        RECT 282.220 61.040 282.550 61.055 ;
        RECT 159.335 60.675 161.335 60.825 ;
        RECT 164.000 60.675 164.330 60.690 ;
        RECT 158.335 60.375 164.330 60.675 ;
        RECT 159.335 60.225 161.335 60.375 ;
        RECT 164.000 60.360 164.330 60.375 ;
        RECT 177.625 60.020 179.205 60.350 ;
        RECT 217.625 60.020 219.205 60.350 ;
        RECT 257.625 60.020 259.205 60.350 ;
        RECT 297.625 60.020 299.205 60.350 ;
        RECT 244.040 59.315 244.370 59.330 ;
        RECT 247.925 59.315 248.305 59.325 ;
        RECT 284.520 59.315 284.850 59.330 ;
        RECT 244.040 59.015 284.850 59.315 ;
        RECT 244.040 59.000 244.370 59.015 ;
        RECT 247.925 59.005 248.305 59.015 ;
        RECT 284.520 59.000 284.850 59.015 ;
        RECT 182.400 58.635 182.730 58.650 ;
        RECT 203.560 58.635 203.890 58.650 ;
        RECT 182.400 58.335 203.890 58.635 ;
        RECT 182.400 58.320 182.730 58.335 ;
        RECT 203.560 58.320 203.890 58.335 ;
        RECT 249.560 58.635 249.890 58.650 ;
        RECT 279.000 58.635 279.330 58.650 ;
        RECT 249.560 58.335 279.330 58.635 ;
        RECT 249.560 58.320 249.890 58.335 ;
        RECT 279.000 58.320 279.330 58.335 ;
        RECT 248.180 57.955 248.510 57.970 ;
        RECT 254.620 57.955 254.950 57.970 ;
        RECT 248.180 57.655 254.950 57.955 ;
        RECT 248.180 57.640 248.510 57.655 ;
        RECT 254.620 57.640 254.950 57.655 ;
        RECT 180.925 57.300 182.505 57.630 ;
        RECT 220.925 57.300 222.505 57.630 ;
        RECT 260.925 57.300 262.505 57.630 ;
        RECT 300.925 57.300 302.505 57.630 ;
        RECT 184.700 57.275 185.030 57.290 ;
        RECT 197.120 57.275 197.450 57.290 ;
        RECT 184.700 56.975 197.450 57.275 ;
        RECT 184.700 56.960 185.030 56.975 ;
        RECT 197.120 56.960 197.450 56.975 ;
        RECT 226.100 57.275 226.430 57.290 ;
        RECT 245.420 57.275 245.750 57.290 ;
        RECT 256.000 57.275 256.330 57.290 ;
        RECT 226.100 56.975 256.330 57.275 ;
        RECT 226.100 56.960 226.430 56.975 ;
        RECT 245.420 56.960 245.750 56.975 ;
        RECT 256.000 56.960 256.330 56.975 ;
        RECT 181.480 56.595 181.810 56.610 ;
        RECT 204.940 56.595 205.270 56.610 ;
        RECT 181.480 56.295 205.270 56.595 ;
        RECT 181.480 56.280 181.810 56.295 ;
        RECT 204.940 56.280 205.270 56.295 ;
        RECT 183.320 55.915 183.650 55.930 ;
        RECT 194.360 55.915 194.690 55.930 ;
        RECT 183.320 55.615 194.690 55.915 ;
        RECT 183.320 55.600 183.650 55.615 ;
        RECT 194.360 55.600 194.690 55.615 ;
        RECT 224.260 55.235 224.590 55.250 ;
        RECT 234.380 55.235 234.710 55.250 ;
        RECT 224.260 54.935 234.710 55.235 ;
        RECT 224.260 54.920 224.590 54.935 ;
        RECT 234.380 54.920 234.710 54.935 ;
        RECT 177.625 54.580 179.205 54.910 ;
        RECT 217.625 54.580 219.205 54.910 ;
        RECT 257.625 54.580 259.205 54.910 ;
        RECT 297.625 54.580 299.205 54.910 ;
        RECT 231.620 54.555 231.950 54.570 ;
        RECT 233.460 54.555 233.790 54.570 ;
        RECT 231.620 54.255 233.790 54.555 ;
        RECT 231.620 54.240 231.950 54.255 ;
        RECT 233.460 54.240 233.790 54.255 ;
        RECT 185.160 52.515 185.490 52.530 ;
        RECT 191.600 52.515 191.930 52.530 ;
        RECT 185.160 52.215 191.930 52.515 ;
        RECT 185.160 52.200 185.490 52.215 ;
        RECT 191.600 52.200 191.930 52.215 ;
        RECT 252.320 52.515 252.650 52.530 ;
        RECT 255.080 52.515 255.410 52.530 ;
        RECT 252.320 52.215 255.410 52.515 ;
        RECT 252.320 52.200 252.650 52.215 ;
        RECT 255.080 52.200 255.410 52.215 ;
        RECT 305.680 52.515 306.010 52.530 ;
        RECT 312.335 52.515 314.335 52.665 ;
        RECT 305.680 52.505 314.335 52.515 ;
        RECT 316.545 52.505 316.845 155.650 ;
        RECT 305.680 52.215 316.845 52.505 ;
        RECT 305.680 52.200 306.010 52.215 ;
        RECT 312.335 52.205 316.845 52.215 ;
        RECT 180.925 51.860 182.505 52.190 ;
        RECT 220.925 51.860 222.505 52.190 ;
        RECT 260.925 51.860 262.505 52.190 ;
        RECT 300.925 51.860 302.505 52.190 ;
        RECT 312.335 52.065 314.335 52.205 ;
        RECT 210.920 51.155 211.250 51.170 ;
        RECT 253.700 51.155 254.030 51.170 ;
        RECT 210.920 50.855 254.030 51.155 ;
        RECT 210.920 50.840 211.250 50.855 ;
        RECT 253.700 50.840 254.030 50.855 ;
        RECT 175.960 50.475 176.290 50.490 ;
        RECT 247.260 50.475 247.590 50.490 ;
        RECT 175.960 50.175 247.590 50.475 ;
        RECT 175.960 50.160 176.290 50.175 ;
        RECT 247.260 50.160 247.590 50.175 ;
        RECT 242.200 49.795 242.530 49.810 ;
        RECT 249.560 49.795 249.890 49.810 ;
        RECT 242.200 49.495 249.890 49.795 ;
        RECT 242.200 49.480 242.530 49.495 ;
        RECT 249.560 49.480 249.890 49.495 ;
        RECT 177.625 49.140 179.205 49.470 ;
        RECT 217.625 49.140 219.205 49.470 ;
        RECT 257.625 49.140 259.205 49.470 ;
        RECT 297.625 49.140 299.205 49.470 ;
        RECT 233.000 47.075 233.330 47.090 ;
        RECT 241.740 47.075 242.070 47.090 ;
        RECT 233.000 46.775 242.070 47.075 ;
        RECT 233.000 46.760 233.330 46.775 ;
        RECT 241.740 46.760 242.070 46.775 ;
        RECT 180.925 46.420 182.505 46.750 ;
        RECT 220.925 46.420 222.505 46.750 ;
        RECT 260.925 46.420 262.505 46.750 ;
        RECT 300.925 46.420 302.505 46.750 ;
        RECT 227.020 45.715 227.350 45.730 ;
        RECT 236.220 45.715 236.550 45.730 ;
        RECT 242.660 45.715 242.990 45.730 ;
        RECT 227.020 45.415 242.990 45.715 ;
        RECT 227.020 45.400 227.350 45.415 ;
        RECT 236.220 45.400 236.550 45.415 ;
        RECT 240.605 44.370 240.905 45.415 ;
        RECT 242.660 45.400 242.990 45.415 ;
        RECT 240.360 44.055 240.905 44.370 ;
        RECT 263.820 44.355 264.150 44.370 ;
        RECT 271.640 44.355 271.970 44.370 ;
        RECT 263.820 44.055 271.970 44.355 ;
        RECT 240.360 44.040 240.690 44.055 ;
        RECT 263.820 44.040 264.150 44.055 ;
        RECT 271.640 44.040 271.970 44.055 ;
        RECT 177.625 43.700 179.205 44.030 ;
        RECT 217.625 43.700 219.205 44.030 ;
        RECT 257.625 43.700 259.205 44.030 ;
        RECT 297.625 43.700 299.205 44.030 ;
        RECT 180.925 40.980 182.505 41.310 ;
        RECT 220.925 40.980 222.505 41.310 ;
        RECT 260.925 40.980 262.505 41.310 ;
        RECT 300.925 40.980 302.505 41.310 ;
        RECT 248.640 39.595 248.970 39.610 ;
        RECT 278.540 39.595 278.870 39.610 ;
        RECT 248.640 39.295 278.870 39.595 ;
        RECT 248.640 39.280 248.970 39.295 ;
        RECT 278.540 39.280 278.870 39.295 ;
        RECT 177.625 38.260 179.205 38.590 ;
        RECT 217.625 38.260 219.205 38.590 ;
        RECT 257.625 38.260 259.205 38.590 ;
        RECT 297.625 38.260 299.205 38.590 ;
        RECT 316.555 36.345 316.955 36.545 ;
        RECT 304.760 36.195 305.090 36.210 ;
        RECT 312.335 36.195 316.955 36.345 ;
        RECT 304.760 35.895 316.955 36.195 ;
        RECT 304.760 35.880 305.090 35.895 ;
        RECT 180.925 35.540 182.505 35.870 ;
        RECT 220.925 35.540 222.505 35.870 ;
        RECT 260.925 35.540 262.505 35.870 ;
        RECT 300.925 35.540 302.505 35.870 ;
        RECT 312.335 35.745 316.955 35.895 ;
        RECT 177.625 32.820 179.205 33.150 ;
        RECT 217.625 32.820 219.205 33.150 ;
        RECT 257.625 32.820 259.205 33.150 ;
        RECT 297.625 32.820 299.205 33.150 ;
        RECT 180.925 30.100 182.505 30.430 ;
        RECT 220.925 30.100 222.505 30.430 ;
        RECT 260.925 30.100 262.505 30.430 ;
        RECT 300.925 30.100 302.505 30.430 ;
        RECT 248.845 28.715 249.225 28.725 ;
        RECT 304.300 28.715 304.630 28.730 ;
        RECT 248.845 28.415 304.630 28.715 ;
        RECT 248.845 28.405 249.225 28.415 ;
        RECT 304.300 28.400 304.630 28.415 ;
        RECT 159.335 28.035 161.335 28.185 ;
        RECT 164.000 28.035 164.330 28.050 ;
        RECT 157.560 27.735 164.330 28.035 ;
        RECT 159.335 27.585 161.335 27.735 ;
        RECT 164.000 27.720 164.330 27.735 ;
        RECT 177.625 27.380 179.205 27.710 ;
        RECT 217.625 27.380 219.205 27.710 ;
        RECT 257.625 27.380 259.205 27.710 ;
        RECT 297.625 27.380 299.205 27.710 ;
        RECT 180.925 24.660 182.505 24.990 ;
        RECT 220.925 24.660 222.505 24.990 ;
        RECT 260.925 24.660 262.505 24.990 ;
        RECT 300.925 24.660 302.505 24.990 ;
        RECT 177.625 21.940 179.205 22.270 ;
        RECT 217.625 21.940 219.205 22.270 ;
        RECT 257.625 21.940 259.205 22.270 ;
        RECT 297.625 21.940 299.205 22.270 ;
        RECT 304.300 19.875 304.630 19.890 ;
        RECT 312.335 19.875 314.335 20.025 ;
        RECT 304.300 19.845 314.335 19.875 ;
        RECT 317.375 19.845 317.675 156.780 ;
        RECT 318.485 36.545 318.785 157.875 ;
        RECT 318.085 35.745 318.785 36.545 ;
        RECT 304.300 19.575 317.675 19.845 ;
        RECT 304.300 19.560 304.630 19.575 ;
        RECT 180.925 19.220 182.505 19.550 ;
        RECT 220.925 19.220 222.505 19.550 ;
        RECT 260.925 19.220 262.505 19.550 ;
        RECT 300.925 19.220 302.505 19.550 ;
        RECT 312.335 19.545 317.675 19.575 ;
        RECT 312.335 19.425 314.335 19.545 ;
        RECT 177.625 16.500 179.205 16.830 ;
        RECT 217.625 16.500 219.205 16.830 ;
        RECT 257.625 16.500 259.205 16.830 ;
        RECT 297.625 16.500 299.205 16.830 ;
        RECT 180.925 13.780 182.505 14.110 ;
        RECT 220.925 13.780 222.505 14.110 ;
        RECT 260.925 13.780 262.505 14.110 ;
        RECT 300.925 13.780 302.505 14.110 ;
        RECT 174.515 5.690 302.515 7.290 ;
        RECT 177.615 2.590 299.215 4.190 ;
      LAYER met4 ;
        RECT 23.260 224.760 23.310 225.560 ;
        RECT 23.610 224.760 23.660 225.560 ;
        RECT 45.340 224.760 45.390 225.560 ;
        RECT 45.690 224.760 45.740 225.560 ;
        RECT 65.010 225.310 65.510 225.710 ;
        RECT 125.730 225.360 126.530 225.760 ;
        RECT 59.490 224.760 59.990 225.160 ;
        RECT 67.770 224.760 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 75.700 224.760 75.750 224.860 ;
        RECT 76.050 224.760 76.100 224.860 ;
        RECT 78.810 224.760 78.945 224.860 ;
        RECT 15.030 224.460 15.330 224.760 ;
        RECT 17.790 224.460 18.090 224.760 ;
        RECT 20.550 224.460 20.850 224.760 ;
        RECT 26.070 224.460 26.370 224.760 ;
        RECT 28.830 224.460 29.130 224.760 ;
        RECT 31.590 224.460 31.890 224.760 ;
        RECT 34.350 224.460 34.650 224.760 ;
        RECT 37.110 224.460 37.410 224.760 ;
        RECT 39.870 224.460 40.170 224.760 ;
        RECT 42.630 224.460 42.930 224.760 ;
        RECT 48.150 224.460 48.450 224.760 ;
        RECT 50.910 224.460 51.210 224.760 ;
        RECT 53.670 224.460 53.970 224.760 ;
        RECT 56.430 224.460 56.730 224.760 ;
        RECT 3.600 224.060 56.730 224.460 ;
        RECT 61.950 224.560 62.250 224.760 ;
        RECT 67.470 224.710 68.270 224.760 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.510 70.530 224.760 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 3.600 220.760 5.200 224.060 ;
        RECT 72.990 223.910 73.290 224.760 ;
        RECT 75.700 224.060 76.100 224.760 ;
        RECT 78.510 224.060 78.945 224.760 ;
        RECT 83.980 224.760 84.030 224.860 ;
        RECT 84.330 224.760 84.380 224.860 ;
        RECT 83.980 224.060 84.380 224.760 ;
        RECT 86.740 224.760 86.790 224.860 ;
        RECT 87.090 224.760 87.140 224.860 ;
        RECT 86.740 224.060 87.140 224.760 ;
        RECT 92.260 224.760 92.310 224.860 ;
        RECT 92.610 224.760 92.660 224.860 ;
        RECT 128.490 224.760 130.195 225.050 ;
        RECT 92.260 224.060 92.660 224.760 ;
        RECT 95.070 224.450 95.370 224.760 ;
        RECT 97.830 224.450 98.130 224.760 ;
        RECT 100.590 224.450 100.890 224.760 ;
        RECT 103.350 224.450 103.650 224.760 ;
        RECT 106.110 224.450 106.410 224.760 ;
        RECT 108.870 224.615 109.170 224.760 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.650 106.460 224.450 ;
        RECT 108.865 224.215 109.665 224.615 ;
        RECT 6.200 221.180 109.540 222.780 ;
        RECT 111.630 221.515 111.930 224.760 ;
        RECT 114.390 222.115 114.690 224.760 ;
        RECT 117.150 222.715 117.450 224.760 ;
        RECT 119.910 223.315 120.210 224.760 ;
        RECT 122.670 223.915 122.970 224.760 ;
        RECT 128.190 224.750 130.195 224.760 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 122.670 223.615 149.190 223.915 ;
        RECT 119.910 223.015 145.160 223.315 ;
        RECT 117.150 222.415 141.130 222.715 ;
        RECT 114.390 221.815 137.100 222.115 ;
        RECT 136.800 221.515 137.100 221.815 ;
        RECT 140.830 221.515 141.130 222.415 ;
        RECT 144.860 221.515 145.160 223.015 ;
        RECT 148.890 221.515 149.190 223.615 ;
      LAYER met4 ;
        RECT 255.465 221.585 317.065 223.185 ;
      LAYER met4 ;
        RECT 111.630 221.215 133.120 221.515 ;
        RECT 6.200 220.760 7.800 221.180 ;
        RECT 10.550 218.590 105.040 220.190 ;
        RECT 7.800 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 103.440 211.240 105.040 218.590 ;
        RECT 106.340 219.305 109.540 221.180 ;
        RECT 132.720 220.715 133.120 221.215 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 106.340 217.705 151.230 219.305 ;
        RECT 106.340 217.515 109.540 217.705 ;
        RECT 106.415 211.240 108.015 213.740 ;
        RECT 27.080 209.940 53.660 210.740 ;
        RECT 27.080 209.640 27.570 209.940 ;
        RECT 16.115 199.365 25.725 208.975 ;
        RECT 16.115 196.975 16.715 199.365 ;
        RECT 16.115 187.365 25.725 196.975 ;
        RECT 16.115 184.975 16.715 187.365 ;
        RECT 16.115 175.365 25.725 184.975 ;
        RECT 16.115 172.975 16.715 175.365 ;
        RECT 16.115 163.365 25.725 172.975 ;
        RECT 16.115 160.975 16.715 163.365 ;
        RECT 16.115 151.365 25.725 160.975 ;
        RECT 16.115 150.210 16.715 151.365 ;
        RECT 27.080 150.970 27.565 209.640 ;
        RECT 28.915 199.365 38.525 208.975 ;
        RECT 37.925 196.975 38.525 199.365 ;
        RECT 28.915 187.365 38.525 196.975 ;
        RECT 52.860 188.465 53.660 209.940 ;
        RECT 103.440 209.640 177.615 211.240 ;
      LAYER met4 ;
        RECT 255.465 207.185 257.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 219.185 271.465 221.585 ;
      LAYER met4 ;
        RECT 271.465 219.585 277.065 221.585 ;
      LAYER met4 ;
        RECT 277.065 219.585 279.465 221.585 ;
      LAYER met4 ;
        RECT 279.465 219.585 285.065 221.585 ;
      LAYER met4 ;
        RECT 285.065 219.585 289.465 221.585 ;
      LAYER met4 ;
        RECT 289.465 219.585 293.065 221.585 ;
      LAYER met4 ;
        RECT 293.065 219.585 297.465 221.585 ;
      LAYER met4 ;
        RECT 297.465 219.585 301.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 209.585 259.465 219.185 ;
      LAYER met4 ;
        RECT 259.465 217.585 269.065 219.185 ;
        RECT 259.465 211.185 261.065 217.585 ;
      LAYER met4 ;
        RECT 261.065 211.185 267.465 217.585 ;
      LAYER met4 ;
        RECT 267.465 211.185 269.065 217.585 ;
        RECT 259.465 209.585 269.065 211.185 ;
      LAYER met4 ;
        RECT 269.065 209.585 271.465 219.185 ;
      LAYER met4 ;
        RECT 271.465 215.185 273.065 219.585 ;
      LAYER met4 ;
        RECT 273.065 217.185 279.465 219.585 ;
      LAYER met4 ;
        RECT 279.465 217.185 283.065 219.585 ;
      LAYER met4 ;
        RECT 283.065 217.185 289.465 219.585 ;
      LAYER met4 ;
        RECT 289.465 217.185 291.065 219.585 ;
      LAYER met4 ;
        RECT 291.065 219.185 299.465 219.585 ;
        RECT 291.065 217.585 295.465 219.185 ;
      LAYER met4 ;
        RECT 295.465 217.585 297.065 219.185 ;
      LAYER met4 ;
        RECT 297.065 217.585 299.465 219.185 ;
        RECT 291.065 217.185 299.465 217.585 ;
        RECT 273.065 215.585 275.465 217.185 ;
      LAYER met4 ;
        RECT 275.465 215.585 291.065 217.185 ;
      LAYER met4 ;
        RECT 291.065 215.585 293.465 217.185 ;
      LAYER met4 ;
        RECT 293.465 215.585 295.065 217.185 ;
      LAYER met4 ;
        RECT 295.065 215.585 299.465 217.185 ;
        RECT 273.065 215.185 277.465 215.585 ;
      LAYER met4 ;
        RECT 271.465 213.585 275.065 215.185 ;
      LAYER met4 ;
        RECT 275.065 213.585 277.465 215.185 ;
      LAYER met4 ;
        RECT 277.465 213.585 281.065 215.585 ;
      LAYER met4 ;
        RECT 281.065 213.585 285.465 215.585 ;
      LAYER met4 ;
        RECT 285.465 213.585 287.065 215.585 ;
      LAYER met4 ;
        RECT 287.065 213.585 289.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 215.185 291.065 215.585 ;
      LAYER met4 ;
        RECT 291.065 215.185 299.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 213.585 293.065 215.185 ;
      LAYER met4 ;
        RECT 293.065 213.585 299.465 215.185 ;
        RECT 257.065 207.185 271.465 209.585 ;
      LAYER met4 ;
        RECT 271.465 207.185 273.065 213.585 ;
      LAYER met4 ;
        RECT 273.065 211.185 279.465 213.585 ;
      LAYER met4 ;
        RECT 255.465 205.585 273.065 207.185 ;
      LAYER met4 ;
        RECT 273.065 205.585 275.465 211.185 ;
      LAYER met4 ;
        RECT 255.465 199.185 257.065 205.585 ;
      LAYER met4 ;
        RECT 257.065 201.585 261.465 205.585 ;
      LAYER met4 ;
        RECT 261.465 203.185 263.065 205.585 ;
      LAYER met4 ;
        RECT 263.065 203.185 265.465 205.585 ;
      LAYER met4 ;
        RECT 265.465 203.585 269.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 205.185 275.465 205.585 ;
      LAYER met4 ;
        RECT 275.465 205.185 277.065 211.185 ;
      LAYER met4 ;
        RECT 277.065 207.585 279.465 211.185 ;
      LAYER met4 ;
        RECT 279.465 207.585 281.065 213.585 ;
      LAYER met4 ;
        RECT 281.065 213.185 299.465 213.585 ;
      LAYER met4 ;
        RECT 299.465 213.185 301.065 219.585 ;
      LAYER met4 ;
        RECT 301.065 219.185 315.465 221.585 ;
        RECT 281.065 207.585 283.465 213.185 ;
      LAYER met4 ;
        RECT 283.465 211.185 285.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.585 295.465 213.185 ;
      LAYER met4 ;
        RECT 295.465 211.585 301.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.185 297.465 211.585 ;
      LAYER met4 ;
        RECT 283.465 209.585 287.065 211.185 ;
      LAYER met4 ;
        RECT 287.065 209.585 289.465 211.185 ;
      LAYER met4 ;
        RECT 289.465 209.585 295.065 211.185 ;
      LAYER met4 ;
        RECT 295.065 209.585 297.465 211.185 ;
      LAYER met4 ;
        RECT 297.465 209.585 301.065 211.585 ;
      LAYER met4 ;
        RECT 301.065 209.585 303.465 219.185 ;
      LAYER met4 ;
        RECT 303.465 217.585 313.065 219.185 ;
        RECT 303.465 211.185 305.065 217.585 ;
      LAYER met4 ;
        RECT 305.065 211.185 311.465 217.585 ;
      LAYER met4 ;
        RECT 311.465 211.185 313.065 217.585 ;
        RECT 303.465 209.585 313.065 211.185 ;
      LAYER met4 ;
        RECT 313.065 209.585 315.465 219.185 ;
      LAYER met4 ;
        RECT 283.465 207.585 285.065 209.585 ;
      LAYER met4 ;
        RECT 285.065 209.185 291.465 209.585 ;
        RECT 285.065 207.585 287.465 209.185 ;
        RECT 277.065 207.185 287.465 207.585 ;
      LAYER met4 ;
        RECT 287.465 207.185 289.065 209.185 ;
      LAYER met4 ;
        RECT 289.065 207.585 291.465 209.185 ;
      LAYER met4 ;
        RECT 291.465 207.585 293.065 209.585 ;
      LAYER met4 ;
        RECT 293.065 209.185 299.465 209.585 ;
        RECT 293.065 207.585 295.465 209.185 ;
        RECT 277.065 205.585 281.465 207.185 ;
      LAYER met4 ;
        RECT 281.465 205.585 283.065 207.185 ;
      LAYER met4 ;
        RECT 283.065 205.585 285.465 207.185 ;
      LAYER met4 ;
        RECT 285.465 205.585 289.065 207.185 ;
      LAYER met4 ;
        RECT 289.065 205.585 295.465 207.585 ;
      LAYER met4 ;
        RECT 295.465 205.585 297.065 209.185 ;
      LAYER met4 ;
        RECT 297.065 205.585 299.465 209.185 ;
      LAYER met4 ;
        RECT 299.465 207.185 301.065 209.585 ;
      LAYER met4 ;
        RECT 301.065 207.185 315.465 209.585 ;
      LAYER met4 ;
        RECT 315.465 207.185 317.065 221.585 ;
        RECT 299.465 205.585 317.065 207.185 ;
      LAYER met4 ;
        RECT 277.065 205.185 287.465 205.585 ;
      LAYER met4 ;
        RECT 287.465 205.185 289.065 205.585 ;
      LAYER met4 ;
        RECT 289.065 205.185 299.465 205.585 ;
      LAYER met4 ;
        RECT 299.465 205.185 301.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 203.585 273.465 205.185 ;
      LAYER met4 ;
        RECT 273.465 203.585 279.065 205.185 ;
      LAYER met4 ;
        RECT 279.065 203.585 283.465 205.185 ;
      LAYER met4 ;
        RECT 283.465 203.585 285.065 205.185 ;
      LAYER met4 ;
        RECT 285.065 203.585 287.465 205.185 ;
      LAYER met4 ;
        RECT 287.465 203.585 295.065 205.185 ;
      LAYER met4 ;
        RECT 295.065 203.585 297.465 205.185 ;
      LAYER met4 ;
        RECT 297.465 203.585 301.065 205.185 ;
      LAYER met4 ;
        RECT 301.065 203.585 307.465 205.585 ;
      LAYER met4 ;
        RECT 307.465 203.585 309.065 205.585 ;
      LAYER met4 ;
        RECT 309.065 203.585 313.465 205.585 ;
      LAYER met4 ;
        RECT 313.465 203.585 317.065 205.585 ;
        RECT 265.465 203.185 267.065 203.585 ;
      LAYER met4 ;
        RECT 267.065 203.185 277.465 203.585 ;
      LAYER met4 ;
        RECT 261.465 201.585 267.065 203.185 ;
      LAYER met4 ;
        RECT 267.065 201.585 269.465 203.185 ;
      LAYER met4 ;
        RECT 269.465 201.585 271.065 203.185 ;
      LAYER met4 ;
        RECT 271.065 201.585 277.465 203.185 ;
        RECT 257.065 201.185 277.465 201.585 ;
      LAYER met4 ;
        RECT 277.465 201.185 279.065 203.585 ;
      LAYER met4 ;
        RECT 279.065 203.185 287.465 203.585 ;
      LAYER met4 ;
        RECT 287.465 203.185 289.065 203.585 ;
      LAYER met4 ;
        RECT 289.065 203.185 297.465 203.585 ;
      LAYER met4 ;
        RECT 297.465 203.185 299.065 203.585 ;
      LAYER met4 ;
        RECT 299.065 203.185 315.465 203.585 ;
        RECT 279.065 201.585 285.465 203.185 ;
      LAYER met4 ;
        RECT 285.465 201.585 289.065 203.185 ;
      LAYER met4 ;
        RECT 289.065 201.585 295.465 203.185 ;
      LAYER met4 ;
        RECT 295.465 201.585 299.065 203.185 ;
      LAYER met4 ;
        RECT 299.065 201.585 303.465 203.185 ;
      LAYER met4 ;
        RECT 303.465 201.585 307.065 203.185 ;
      LAYER met4 ;
        RECT 257.065 199.185 271.465 201.185 ;
      LAYER met4 ;
        RECT 271.465 199.185 273.065 201.185 ;
      LAYER met4 ;
        RECT 273.065 199.585 275.465 201.185 ;
      LAYER met4 ;
        RECT 275.465 199.585 279.065 201.185 ;
      LAYER met4 ;
        RECT 279.065 199.585 287.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 201.185 289.065 201.585 ;
      LAYER met4 ;
        RECT 289.065 201.185 305.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 199.585 291.065 201.185 ;
      LAYER met4 ;
        RECT 291.065 199.585 299.465 201.185 ;
      LAYER met4 ;
        RECT 299.465 199.585 301.065 201.185 ;
      LAYER met4 ;
        RECT 301.065 199.585 305.465 201.185 ;
        RECT 273.065 199.185 287.465 199.585 ;
      LAYER met4 ;
        RECT 287.465 199.185 289.065 199.585 ;
      LAYER met4 ;
        RECT 289.065 199.185 305.465 199.585 ;
      LAYER met4 ;
        RECT 305.465 199.185 307.065 201.585 ;
      LAYER met4 ;
        RECT 307.065 201.185 315.465 203.185 ;
      LAYER met4 ;
        RECT 315.465 201.185 317.065 203.585 ;
      LAYER met4 ;
        RECT 307.065 199.185 313.465 201.185 ;
      LAYER met4 ;
        RECT 255.465 195.185 259.065 199.185 ;
      LAYER met4 ;
        RECT 259.065 197.585 261.465 199.185 ;
        POLYGON 261.465 199.185 261.770 199.185 261.465 198.880 ;
      LAYER met4 ;
        RECT 261.770 198.880 273.065 199.185 ;
        RECT 261.465 197.585 273.065 198.880 ;
      LAYER met4 ;
        RECT 273.065 197.585 285.465 199.185 ;
      LAYER met4 ;
        RECT 285.465 197.585 289.065 199.185 ;
      LAYER met4 ;
        RECT 289.065 197.585 291.465 199.185 ;
      LAYER met4 ;
        RECT 291.465 197.585 293.065 199.185 ;
      LAYER met4 ;
        RECT 293.065 197.585 301.465 199.185 ;
      LAYER met4 ;
        RECT 301.465 197.585 309.065 199.185 ;
      LAYER met4 ;
        RECT 309.065 197.585 313.465 199.185 ;
      LAYER met4 ;
        RECT 313.465 197.585 317.065 201.185 ;
      LAYER met4 ;
        RECT 259.065 195.585 265.465 197.585 ;
      LAYER met4 ;
        RECT 265.465 195.585 267.065 197.585 ;
      LAYER met4 ;
        RECT 267.065 197.185 287.465 197.585 ;
      LAYER met4 ;
        RECT 287.465 197.185 289.065 197.585 ;
      LAYER met4 ;
        RECT 289.065 197.185 303.465 197.585 ;
        RECT 267.065 195.585 275.465 197.185 ;
        RECT 259.065 195.185 275.465 195.585 ;
      LAYER met4 ;
        RECT 275.465 195.185 277.065 197.185 ;
      LAYER met4 ;
        RECT 277.065 195.185 281.465 197.185 ;
      LAYER met4 ;
        RECT 281.465 195.585 285.065 197.185 ;
      LAYER met4 ;
        RECT 285.065 195.585 287.465 197.185 ;
      LAYER met4 ;
        RECT 255.465 193.585 263.065 195.185 ;
      LAYER met4 ;
        RECT 263.065 193.585 269.465 195.185 ;
      LAYER met4 ;
        RECT 269.465 193.585 273.065 195.185 ;
      LAYER met4 ;
        RECT 273.065 193.585 275.465 195.185 ;
      LAYER met4 ;
        RECT 255.465 191.585 259.065 193.585 ;
      LAYER met4 ;
        RECT 259.065 193.185 275.465 193.585 ;
        RECT 259.065 191.585 263.465 193.185 ;
      LAYER met4 ;
        RECT 263.465 191.585 269.065 193.185 ;
      LAYER met4 ;
        RECT 269.065 191.585 275.465 193.185 ;
        RECT 186.310 189.425 186.640 189.755 ;
        RECT 207.470 189.425 207.800 189.755 ;
        RECT 110.530 187.540 156.765 189.140 ;
        RECT 37.925 184.975 38.525 187.365 ;
        RECT 28.915 175.365 38.525 184.975 ;
        RECT 37.925 172.975 38.525 175.365 ;
        RECT 28.915 163.365 38.525 172.975 ;
        RECT 51.950 184.940 103.750 186.540 ;
        RECT 51.950 169.890 53.550 184.940 ;
        RECT 57.020 177.390 109.070 178.990 ;
        RECT 153.565 178.210 156.765 187.540 ;
        RECT 151.155 175.010 156.765 178.210 ;
        RECT 186.325 175.475 186.625 189.425 ;
        RECT 186.310 175.145 186.640 175.475 ;
        RECT 51.950 168.290 58.420 169.890 ;
        RECT 37.925 160.975 38.525 163.365 ;
        RECT 28.915 151.365 38.525 160.975 ;
        RECT 111.685 158.165 112.085 158.565 ;
        RECT 105.385 157.765 112.085 158.165 ;
        RECT 105.385 157.365 105.785 157.765 ;
        RECT 109.415 156.565 109.815 156.965 ;
        RECT 113.085 156.565 113.485 156.965 ;
        RECT 109.415 156.165 113.485 156.565 ;
        RECT 37.925 150.210 38.525 151.365 ;
        RECT 16.115 149.410 46.630 150.210 ;
        RECT 51.575 145.090 73.495 148.290 ;
        RECT 9.490 135.030 17.100 142.640 ;
        RECT 18.455 142.175 20.750 142.975 ;
        RECT 13.385 130.025 14.185 135.030 ;
        RECT 18.455 134.695 18.935 142.175 ;
        RECT 20.350 141.375 20.750 142.175 ;
        RECT 61.980 135.495 62.780 135.895 ;
        RECT 61.980 135.095 140.370 135.495 ;
        RECT 22.615 133.320 80.925 134.120 ;
        RECT 20.650 131.810 21.050 132.210 ;
        RECT 137.945 131.810 138.345 132.210 ;
        RECT 20.650 131.410 138.345 131.810 ;
        RECT 139.120 130.025 139.520 132.990 ;
        RECT 13.385 129.625 139.520 130.025 ;
        RECT 16.805 128.710 139.520 129.110 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 128.710 ;
        RECT 139.970 125.690 140.370 135.095 ;
        RECT 140.940 131.390 142.100 132.990 ;
        RECT 140.940 125.060 141.340 131.390 ;
        RECT 131.145 124.660 141.340 125.060 ;
        RECT 103.315 121.565 118.965 123.165 ;
        RECT 109.865 107.965 118.715 109.565 ;
        RECT 63.315 103.465 74.365 105.065 ;
        RECT 105.965 103.615 118.565 105.215 ;
        RECT 131.145 98.015 131.545 124.660 ;
        RECT 153.565 124.090 156.765 175.010 ;
        RECT 207.485 174.795 207.785 189.425 ;
      LAYER met4 ;
        RECT 255.465 189.185 257.065 191.585 ;
      LAYER met4 ;
        RECT 257.065 191.185 263.465 191.585 ;
        RECT 257.065 189.585 259.465 191.185 ;
      LAYER met4 ;
        RECT 259.465 189.585 261.065 191.185 ;
      LAYER met4 ;
        RECT 261.065 189.585 263.465 191.185 ;
      LAYER met4 ;
        RECT 263.465 189.585 267.065 191.585 ;
      LAYER met4 ;
        RECT 267.065 191.185 275.465 191.585 ;
      LAYER met4 ;
        RECT 275.465 191.185 279.065 195.185 ;
      LAYER met4 ;
        RECT 267.065 189.585 269.465 191.185 ;
      LAYER met4 ;
        RECT 269.465 189.585 271.065 191.185 ;
      LAYER met4 ;
        RECT 271.065 189.585 273.465 191.185 ;
      LAYER met4 ;
        RECT 273.465 189.585 279.065 191.185 ;
      LAYER met4 ;
        RECT 279.065 189.585 281.465 195.185 ;
      LAYER met4 ;
        RECT 281.465 191.185 283.065 195.585 ;
      LAYER met4 ;
        RECT 283.065 191.585 287.465 195.585 ;
      LAYER met4 ;
        RECT 287.465 191.585 291.065 197.185 ;
      LAYER met4 ;
        RECT 291.065 191.585 293.465 197.185 ;
      LAYER met4 ;
        RECT 293.465 193.185 295.065 197.185 ;
      LAYER met4 ;
        RECT 295.065 195.185 303.465 197.185 ;
      LAYER met4 ;
        RECT 303.465 195.185 307.065 197.585 ;
      LAYER met4 ;
        RECT 307.065 197.185 315.465 197.585 ;
        RECT 295.065 193.185 299.465 195.185 ;
      LAYER met4 ;
        RECT 299.465 193.585 307.065 195.185 ;
        RECT 299.465 193.185 301.065 193.585 ;
        RECT 293.465 191.585 301.065 193.185 ;
      LAYER met4 ;
        RECT 301.065 191.585 303.465 193.585 ;
      LAYER met4 ;
        RECT 303.465 191.585 307.065 193.585 ;
      LAYER met4 ;
        RECT 307.065 191.585 309.465 197.185 ;
      LAYER met4 ;
        RECT 309.465 195.185 311.065 197.185 ;
      LAYER met4 ;
        RECT 311.065 195.185 315.465 197.185 ;
      LAYER met4 ;
        RECT 315.465 195.185 317.065 197.585 ;
        RECT 309.465 193.585 317.065 195.185 ;
      LAYER met4 ;
        RECT 283.065 191.185 297.465 191.585 ;
      LAYER met4 ;
        RECT 281.465 189.585 287.065 191.185 ;
      LAYER met4 ;
        RECT 257.065 189.185 263.465 189.585 ;
      LAYER met4 ;
        RECT 263.465 189.185 265.065 189.585 ;
      LAYER met4 ;
        RECT 265.065 189.185 273.465 189.585 ;
        RECT 209.310 185.345 209.640 185.675 ;
      LAYER met4 ;
        RECT 255.465 185.585 259.065 189.185 ;
      LAYER met4 ;
        RECT 259.065 185.585 261.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 187.890 265.065 189.185 ;
        RECT 261.465 187.585 264.760 187.890 ;
        POLYGON 264.760 187.890 265.065 187.890 264.760 187.585 ;
      LAYER met4 ;
        RECT 265.065 187.585 267.465 189.185 ;
      LAYER met4 ;
        RECT 267.465 187.585 269.065 189.185 ;
      LAYER met4 ;
        RECT 269.065 187.585 273.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 185.585 263.065 187.585 ;
      LAYER met4 ;
        RECT 263.065 187.185 273.465 187.585 ;
      LAYER met4 ;
        RECT 273.465 187.185 275.065 189.585 ;
      LAYER met4 ;
        RECT 275.065 187.585 277.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 189.185 279.065 189.585 ;
      LAYER met4 ;
        RECT 279.065 189.185 285.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 187.585 281.065 189.185 ;
      LAYER met4 ;
        RECT 281.065 187.585 285.465 189.185 ;
      LAYER met4 ;
        RECT 285.465 187.585 287.065 189.585 ;
      LAYER met4 ;
        RECT 287.065 189.185 297.465 191.185 ;
        RECT 287.065 187.585 289.465 189.185 ;
        RECT 263.065 185.585 269.465 187.185 ;
      LAYER met4 ;
        RECT 269.465 185.585 275.065 187.185 ;
      LAYER met4 ;
        RECT 275.065 185.585 279.465 187.585 ;
      LAYER met4 ;
        RECT 279.465 185.585 281.065 187.585 ;
      LAYER met4 ;
        RECT 281.065 187.185 289.465 187.585 ;
      LAYER met4 ;
        RECT 289.465 187.185 291.065 189.185 ;
      LAYER met4 ;
        RECT 291.065 187.585 293.465 189.185 ;
      LAYER met4 ;
        RECT 293.465 187.585 295.065 189.185 ;
      LAYER met4 ;
        RECT 295.065 187.585 297.465 189.185 ;
        RECT 291.065 187.185 297.465 187.585 ;
      LAYER met4 ;
        RECT 297.465 187.185 299.065 191.585 ;
      LAYER met4 ;
        RECT 299.065 189.185 303.465 191.585 ;
      LAYER met4 ;
        RECT 303.465 189.185 305.065 191.585 ;
      LAYER met4 ;
        RECT 305.065 191.185 309.465 191.585 ;
      LAYER met4 ;
        RECT 309.465 191.185 311.065 193.585 ;
      LAYER met4 ;
        RECT 311.065 191.185 315.465 193.585 ;
      LAYER met4 ;
        RECT 315.465 191.185 317.065 193.585 ;
      LAYER met4 ;
        RECT 305.065 189.585 307.465 191.185 ;
      LAYER met4 ;
        RECT 307.465 189.585 317.065 191.185 ;
      LAYER met4 ;
        RECT 305.065 189.185 309.465 189.585 ;
        RECT 299.065 187.585 301.465 189.185 ;
      LAYER met4 ;
        RECT 301.465 187.585 307.065 189.185 ;
      LAYER met4 ;
        RECT 307.065 187.585 309.465 189.185 ;
      LAYER met4 ;
        RECT 309.465 187.585 313.065 189.585 ;
      LAYER met4 ;
        RECT 313.065 187.585 315.465 189.585 ;
        RECT 281.065 185.585 287.465 187.185 ;
      LAYER met4 ;
        RECT 287.465 185.585 293.065 187.185 ;
      LAYER met4 ;
        RECT 293.065 185.585 295.465 187.185 ;
        RECT 209.325 180.235 209.625 185.345 ;
      LAYER met4 ;
        RECT 255.465 183.185 257.065 185.585 ;
      LAYER met4 ;
        RECT 257.065 185.185 273.465 185.585 ;
      LAYER met4 ;
        RECT 273.465 185.185 275.065 185.585 ;
      LAYER met4 ;
        RECT 275.065 185.185 287.465 185.585 ;
        RECT 257.065 183.185 259.465 185.185 ;
      LAYER met4 ;
        RECT 259.465 183.185 261.065 185.185 ;
      LAYER met4 ;
        RECT 261.065 183.185 263.465 185.185 ;
      LAYER met4 ;
        RECT 263.465 183.185 265.065 185.185 ;
      LAYER met4 ;
        RECT 265.065 183.185 273.465 185.185 ;
      LAYER met4 ;
        RECT 273.465 183.585 277.065 185.185 ;
      LAYER met4 ;
        RECT 277.065 183.585 283.465 185.185 ;
      LAYER met4 ;
        RECT 255.465 181.585 265.065 183.185 ;
      LAYER met4 ;
        RECT 265.065 181.585 267.465 183.185 ;
      LAYER met4 ;
        RECT 267.465 181.585 271.065 183.185 ;
      LAYER met4 ;
        RECT 271.065 181.585 273.465 183.185 ;
        RECT 209.310 179.905 209.640 180.235 ;
        RECT 223.110 179.225 223.440 179.555 ;
        RECT 223.125 175.475 223.425 179.225 ;
      LAYER met4 ;
        RECT 255.465 179.185 257.065 181.585 ;
      LAYER met4 ;
        RECT 257.065 179.185 259.465 181.585 ;
      LAYER met4 ;
        RECT 259.465 179.185 265.065 181.585 ;
      LAYER met4 ;
        RECT 265.065 181.185 273.465 181.585 ;
      LAYER met4 ;
        RECT 273.465 181.185 275.065 183.585 ;
      LAYER met4 ;
        RECT 275.065 183.185 283.465 183.585 ;
        RECT 275.065 181.185 279.465 183.185 ;
      LAYER met4 ;
        RECT 279.465 181.185 281.065 183.185 ;
      LAYER met4 ;
        RECT 281.065 181.185 283.465 183.185 ;
      LAYER met4 ;
        RECT 283.465 181.185 285.065 185.185 ;
      LAYER met4 ;
        RECT 285.065 183.585 287.465 185.185 ;
      LAYER met4 ;
        RECT 287.465 183.585 289.065 185.585 ;
      LAYER met4 ;
        RECT 289.065 183.585 295.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 185.185 299.065 187.185 ;
      LAYER met4 ;
        RECT 299.065 185.585 303.465 187.585 ;
      LAYER met4 ;
        RECT 303.465 185.585 307.065 187.585 ;
      LAYER met4 ;
        RECT 307.065 185.585 315.465 187.585 ;
        RECT 299.065 185.185 315.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 183.585 303.065 185.185 ;
      LAYER met4 ;
        RECT 303.065 183.585 307.465 185.185 ;
        RECT 285.065 183.185 299.465 183.585 ;
        RECT 285.065 181.585 293.465 183.185 ;
      LAYER met4 ;
        RECT 293.465 181.585 295.065 183.185 ;
      LAYER met4 ;
        RECT 295.065 181.585 299.465 183.185 ;
      LAYER met4 ;
        RECT 299.465 181.585 301.065 183.585 ;
      LAYER met4 ;
        RECT 301.065 183.185 307.465 183.585 ;
      LAYER met4 ;
        RECT 307.465 183.185 311.065 185.185 ;
      LAYER met4 ;
        RECT 311.065 183.185 315.465 185.185 ;
      LAYER met4 ;
        RECT 315.465 183.185 317.065 189.585 ;
      LAYER met4 ;
        RECT 301.065 181.585 303.465 183.185 ;
      LAYER met4 ;
        RECT 303.465 181.585 305.065 183.185 ;
      LAYER met4 ;
        RECT 305.065 181.585 307.465 183.185 ;
      LAYER met4 ;
        RECT 307.465 181.585 317.065 183.185 ;
      LAYER met4 ;
        RECT 285.065 181.185 307.465 181.585 ;
        RECT 265.065 179.185 271.465 181.185 ;
      LAYER met4 ;
        RECT 271.465 179.585 275.065 181.185 ;
      LAYER met4 ;
        RECT 275.065 179.585 277.465 181.185 ;
      LAYER met4 ;
        RECT 277.465 179.890 293.065 181.185 ;
      LAYER met4 ;
        POLYGON 277.465 179.890 277.770 179.585 277.465 179.585 ;
      LAYER met4 ;
        RECT 277.770 179.585 293.065 179.890 ;
        RECT 271.465 179.185 273.065 179.585 ;
        RECT 255.465 177.585 273.065 179.185 ;
      LAYER met4 ;
        RECT 223.110 175.145 223.440 175.475 ;
        RECT 207.470 174.465 207.800 174.795 ;
      LAYER met4 ;
        RECT 255.465 163.185 257.065 177.585 ;
      LAYER met4 ;
        RECT 257.065 175.185 271.465 177.585 ;
      LAYER met4 ;
        RECT 271.465 175.185 273.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 177.185 281.465 179.585 ;
      LAYER met4 ;
        RECT 281.465 177.185 285.065 179.585 ;
      LAYER met4 ;
        RECT 285.065 177.185 287.465 179.585 ;
      LAYER met4 ;
        RECT 287.465 179.185 293.065 179.585 ;
      LAYER met4 ;
        RECT 293.065 179.185 307.465 181.185 ;
      LAYER met4 ;
        RECT 287.465 177.585 295.065 179.185 ;
        RECT 287.465 177.185 289.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 175.585 277.465 177.185 ;
      LAYER met4 ;
        RECT 277.465 175.585 289.065 177.185 ;
      LAYER met4 ;
        RECT 289.065 175.585 293.465 177.585 ;
      LAYER met4 ;
        RECT 293.465 177.185 295.065 177.585 ;
      LAYER met4 ;
        RECT 295.065 177.185 299.465 179.185 ;
      LAYER met4 ;
        RECT 299.465 177.585 305.065 179.185 ;
      LAYER met4 ;
        RECT 305.065 177.585 307.465 179.185 ;
      LAYER met4 ;
        RECT 307.465 177.585 309.065 181.585 ;
      LAYER met4 ;
        RECT 309.065 177.585 315.465 181.585 ;
      LAYER met4 ;
        RECT 293.465 175.585 297.065 177.185 ;
      LAYER met4 ;
        RECT 273.065 175.185 279.465 175.585 ;
        RECT 257.065 165.585 259.465 175.185 ;
      LAYER met4 ;
        RECT 259.465 173.585 269.065 175.185 ;
        RECT 259.465 167.185 261.065 173.585 ;
      LAYER met4 ;
        RECT 261.065 167.185 267.465 173.585 ;
      LAYER met4 ;
        RECT 267.465 167.185 269.065 173.585 ;
        RECT 259.465 165.585 269.065 167.185 ;
      LAYER met4 ;
        RECT 269.065 165.585 271.465 175.185 ;
      LAYER met4 ;
        RECT 271.465 173.585 277.065 175.185 ;
      LAYER met4 ;
        RECT 277.065 173.585 279.465 175.185 ;
      LAYER met4 ;
        RECT 279.465 173.585 285.065 175.585 ;
      LAYER met4 ;
        RECT 285.065 175.185 295.465 175.585 ;
      LAYER met4 ;
        RECT 271.465 171.585 275.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 173.185 279.465 173.585 ;
      LAYER met4 ;
        RECT 279.465 173.185 281.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 171.585 277.465 173.185 ;
      LAYER met4 ;
        RECT 277.465 171.585 281.065 173.185 ;
      LAYER met4 ;
        RECT 281.065 171.585 283.465 173.585 ;
      LAYER met4 ;
        RECT 283.465 173.185 285.065 173.585 ;
      LAYER met4 ;
        RECT 285.065 173.185 289.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.585 293.065 175.185 ;
      LAYER met4 ;
        RECT 293.065 173.585 295.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.185 291.065 173.585 ;
      LAYER met4 ;
        RECT 291.065 173.185 295.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 173.185 297.065 175.585 ;
      LAYER met4 ;
        RECT 297.065 173.585 299.465 177.185 ;
      LAYER met4 ;
        RECT 299.465 175.185 301.065 177.585 ;
      LAYER met4 ;
        RECT 301.065 175.185 303.465 177.585 ;
      LAYER met4 ;
        RECT 303.465 175.185 305.065 177.585 ;
      LAYER met4 ;
        RECT 305.065 177.185 315.465 177.585 ;
      LAYER met4 ;
        RECT 315.465 177.185 317.065 181.585 ;
      LAYER met4 ;
        RECT 305.065 175.585 309.465 177.185 ;
      LAYER met4 ;
        RECT 309.465 175.585 311.065 177.185 ;
      LAYER met4 ;
        RECT 311.065 175.585 313.465 177.185 ;
        RECT 305.065 175.185 313.465 175.585 ;
      LAYER met4 ;
        RECT 313.465 175.185 317.065 177.185 ;
        RECT 299.465 173.585 305.065 175.185 ;
      LAYER met4 ;
        RECT 305.065 173.585 307.465 175.185 ;
      LAYER met4 ;
        RECT 283.465 171.585 291.065 173.185 ;
      LAYER met4 ;
        RECT 291.065 171.585 293.465 173.185 ;
      LAYER met4 ;
        RECT 293.465 171.890 297.065 173.185 ;
      LAYER met4 ;
        POLYGON 293.465 171.890 293.770 171.585 293.465 171.585 ;
      LAYER met4 ;
        RECT 293.770 171.585 297.065 171.890 ;
        RECT 271.465 169.185 273.065 171.585 ;
      LAYER met4 ;
        RECT 273.065 171.185 283.465 171.585 ;
        RECT 273.065 169.585 275.465 171.185 ;
      LAYER met4 ;
        RECT 275.465 169.585 277.065 171.185 ;
      LAYER met4 ;
        RECT 277.065 169.585 283.465 171.185 ;
        RECT 273.065 169.185 283.465 169.585 ;
      LAYER met4 ;
        RECT 271.465 167.585 275.065 169.185 ;
      LAYER met4 ;
        RECT 275.065 167.585 279.465 169.185 ;
        RECT 257.065 163.185 271.465 165.585 ;
      LAYER met4 ;
        RECT 271.465 163.185 273.065 167.585 ;
      LAYER met4 ;
        RECT 273.065 167.185 279.465 167.585 ;
      LAYER met4 ;
        RECT 279.465 167.185 281.065 169.185 ;
      LAYER met4 ;
        RECT 281.065 167.585 283.465 169.185 ;
      LAYER met4 ;
        RECT 283.465 167.585 289.065 171.585 ;
      LAYER met4 ;
        RECT 289.065 169.585 295.465 171.585 ;
      LAYER met4 ;
        RECT 295.465 171.185 297.065 171.585 ;
      LAYER met4 ;
        RECT 297.065 171.185 307.465 173.585 ;
      LAYER met4 ;
        RECT 307.465 173.185 309.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.585 311.465 175.185 ;
      LAYER met4 ;
        RECT 311.465 173.585 317.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.185 315.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 169.585 301.065 171.185 ;
      LAYER met4 ;
        RECT 301.065 169.585 307.465 171.185 ;
      LAYER met4 ;
        RECT 307.465 169.585 311.065 173.185 ;
      LAYER met4 ;
        RECT 311.065 171.185 315.465 173.185 ;
      LAYER met4 ;
        RECT 315.465 171.185 317.065 173.585 ;
      LAYER met4 ;
        RECT 311.065 169.585 313.465 171.185 ;
      LAYER met4 ;
        RECT 313.465 169.585 317.065 171.185 ;
      LAYER met4 ;
        RECT 289.065 169.185 297.465 169.585 ;
        RECT 289.065 167.585 293.465 169.185 ;
        RECT 273.065 165.585 275.465 167.185 ;
      LAYER met4 ;
        RECT 275.465 165.585 281.065 167.185 ;
      LAYER met4 ;
        RECT 281.065 165.585 293.465 167.585 ;
      LAYER met4 ;
        RECT 293.465 167.185 295.065 169.185 ;
      LAYER met4 ;
        RECT 295.065 167.585 297.465 169.185 ;
      LAYER met4 ;
        RECT 297.465 167.585 299.065 169.585 ;
      LAYER met4 ;
        RECT 299.065 169.185 315.465 169.585 ;
        RECT 299.065 167.585 301.465 169.185 ;
        RECT 295.065 167.185 301.465 167.585 ;
        RECT 273.065 163.185 277.465 165.585 ;
      LAYER met4 ;
        RECT 277.465 163.185 279.065 165.585 ;
      LAYER met4 ;
        RECT 279.065 165.185 293.465 165.585 ;
        RECT 279.065 163.185 281.465 165.185 ;
      LAYER met4 ;
        RECT 281.465 163.185 283.065 165.185 ;
      LAYER met4 ;
        RECT 283.065 163.185 287.465 165.185 ;
      LAYER met4 ;
        RECT 287.465 163.185 289.065 165.185 ;
      LAYER met4 ;
        RECT 289.065 163.185 293.465 165.185 ;
      LAYER met4 ;
        RECT 293.465 163.185 297.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.585 301.465 167.185 ;
      LAYER met4 ;
        RECT 301.465 165.585 305.065 169.185 ;
      LAYER met4 ;
        RECT 305.065 167.585 311.465 169.185 ;
      LAYER met4 ;
        RECT 311.465 167.585 313.065 169.185 ;
      LAYER met4 ;
        RECT 313.065 167.585 315.465 169.185 ;
        RECT 305.065 167.185 315.465 167.585 ;
      LAYER met4 ;
        RECT 315.465 167.185 317.065 169.585 ;
      LAYER met4 ;
        RECT 305.065 165.585 307.465 167.185 ;
      LAYER met4 ;
        RECT 307.465 165.585 311.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.185 309.465 165.585 ;
        RECT 297.065 163.185 305.465 165.185 ;
      LAYER met4 ;
        RECT 305.465 163.185 307.065 165.185 ;
      LAYER met4 ;
        RECT 307.065 163.185 309.465 165.185 ;
      LAYER met4 ;
        RECT 309.465 163.185 311.065 165.585 ;
      LAYER met4 ;
        RECT 311.065 163.185 313.465 167.185 ;
      LAYER met4 ;
        RECT 313.465 163.185 317.065 167.185 ;
        RECT 255.465 161.585 317.065 163.185 ;
      LAYER met4 ;
        RECT 142.760 122.490 156.765 124.090 ;
        RECT 153.565 114.150 156.765 122.490 ;
        RECT 139.355 113.350 156.765 114.150 ;
        RECT 100.115 96.415 132.145 98.015 ;
        RECT 97.165 93.265 124.815 94.865 ;
        RECT 43.135 78.605 52.745 82.655 ;
        RECT 56.135 78.605 65.745 82.655 ;
        RECT 69.135 78.605 78.745 82.655 ;
        RECT 82.135 78.605 91.745 82.655 ;
        RECT 95.135 78.605 104.745 82.655 ;
        RECT 130.545 78.605 132.145 96.415 ;
        RECT 38.470 77.005 132.145 78.605 ;
        RECT 38.470 63.590 39.745 77.005 ;
        RECT 43.135 73.045 52.745 77.005 ;
        RECT 56.135 73.045 65.745 77.005 ;
        RECT 69.135 73.045 78.745 77.005 ;
        RECT 82.135 73.045 91.745 77.005 ;
        RECT 95.135 73.045 104.745 77.005 ;
        RECT 42.800 71.180 108.800 71.690 ;
        RECT 133.525 71.180 135.125 110.315 ;
        RECT 42.800 69.580 135.125 71.180 ;
        RECT 42.800 69.190 108.800 69.580 ;
        RECT 43.135 63.590 52.745 67.835 ;
        RECT 56.135 63.590 65.745 67.835 ;
        RECT 69.135 63.590 78.745 67.835 ;
        RECT 82.135 63.590 91.745 67.835 ;
        RECT 95.135 63.590 104.745 67.835 ;
        RECT 38.470 61.990 104.745 63.590 ;
        RECT 43.135 58.225 52.745 61.990 ;
        RECT 56.135 58.225 65.745 61.990 ;
        RECT 69.135 58.225 78.745 61.990 ;
        RECT 82.135 58.225 91.745 61.990 ;
        RECT 95.135 58.225 104.745 61.990 ;
        RECT 12.915 45.565 92.315 47.165 ;
        RECT 65.765 42.615 117.715 44.215 ;
        RECT 68.865 40.015 120.815 41.615 ;
        RECT 72.095 9.265 82.535 10.865 ;
        RECT 153.565 8.890 156.765 113.350 ;
        RECT 256.230 94.360 256.560 94.690 ;
        RECT 248.870 80.080 249.200 80.410 ;
        RECT 248.885 73.475 249.185 80.080 ;
        RECT 247.965 73.175 249.185 73.475 ;
        RECT 247.965 59.330 248.265 73.175 ;
        RECT 256.245 72.930 256.545 94.360 ;
        RECT 256.230 72.600 256.560 72.930 ;
        RECT 256.245 70.890 256.545 72.600 ;
        RECT 256.230 70.560 256.560 70.890 ;
        RECT 248.870 66.480 249.200 66.810 ;
        RECT 247.950 59.000 248.280 59.330 ;
        RECT 248.885 28.730 249.185 66.480 ;
        RECT 248.870 28.400 249.200 28.730 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.160 7.290 156.765 8.890 ;
        RECT 128.160 5.690 176.115 7.290 ;
        RECT 97.530 1.000 98.430 2.125 ;
        RECT 116.850 1.750 132.465 2.650 ;
        RECT 136.170 1.750 152.360 2.650 ;
        RECT 257.615 2.590 259.215 120.775 ;
        RECT 259.910 86.880 260.240 87.210 ;
        RECT 259.925 78.370 260.225 86.880 ;
        RECT 259.910 78.040 260.240 78.370 ;
        RECT 259.910 77.360 260.240 77.690 ;
        RECT 259.925 73.610 260.225 77.360 ;
        RECT 259.910 73.280 260.240 73.610 ;
        RECT 260.915 5.690 262.515 123.580 ;
        RECT 263.590 92.320 263.920 92.650 ;
        RECT 263.605 70.890 263.905 92.320 ;
        RECT 263.590 70.560 263.920 70.890 ;
        RECT 297.615 2.590 299.215 120.775 ;
        RECT 300.915 5.690 302.515 123.580 ;
        RECT 116.850 1.000 117.750 1.750 ;
        RECT 136.170 1.000 137.070 1.750 ;
  END
END tt_um_cw_vref
END LIBRARY

